magic
tech sky130B
magscale 1 2
timestamp 1682098054
<< viali >>
rect 40233 61353 40267 61387
rect 46857 61353 46891 61387
rect 49433 61353 49467 61387
rect 51457 61353 51491 61387
rect 9689 61285 9723 61319
rect 20729 61285 20763 61319
rect 38485 61285 38519 61319
rect 43729 61285 43763 61319
rect 52285 61285 52319 61319
rect 3065 61217 3099 61251
rect 10425 61217 10459 61251
rect 18153 61217 18187 61251
rect 48053 61217 48087 61251
rect 53389 61217 53423 61251
rect 1685 61149 1719 61183
rect 2789 61149 2823 61183
rect 4353 61149 4387 61183
rect 5089 61149 5123 61183
rect 5733 61149 5767 61183
rect 6653 61149 6687 61183
rect 7573 61149 7607 61183
rect 9505 61149 9539 61183
rect 10241 61149 10275 61183
rect 10977 61149 11011 61183
rect 11989 61149 12023 61183
rect 12725 61149 12759 61183
rect 13001 61149 13035 61183
rect 14933 61149 14967 61183
rect 16129 61149 16163 61183
rect 17233 61149 17267 61183
rect 17969 61149 18003 61183
rect 18705 61149 18739 61183
rect 19809 61149 19843 61183
rect 20545 61149 20579 61183
rect 21281 61149 21315 61183
rect 22385 61149 22419 61183
rect 23857 61149 23891 61183
rect 25329 61149 25363 61183
rect 26249 61149 26283 61183
rect 27261 61149 27295 61183
rect 28273 61149 28307 61183
rect 29837 61149 29871 61183
rect 31217 61149 31251 61183
rect 32413 61149 32447 61183
rect 33333 61149 33367 61183
rect 34069 61149 34103 61183
rect 35725 61149 35759 61183
rect 36461 61149 36495 61183
rect 37565 61149 37599 61183
rect 38301 61149 38335 61183
rect 38945 61149 38979 61183
rect 40141 61149 40175 61183
rect 41613 61149 41647 61183
rect 42625 61149 42659 61183
rect 43545 61149 43579 61183
rect 44373 61149 44407 61183
rect 45293 61149 45327 61183
rect 46029 61149 46063 61183
rect 46765 61149 46799 61183
rect 47869 61149 47903 61183
rect 48605 61149 48639 61183
rect 49341 61149 49375 61183
rect 50445 61149 50479 61183
rect 51365 61149 51399 61183
rect 52101 61149 52135 61183
rect 53205 61149 53239 61183
rect 54125 61149 54159 61183
rect 55505 61149 55539 61183
rect 56517 61149 56551 61183
rect 58173 61149 58207 61183
rect 2237 61081 2271 61115
rect 4537 61081 4571 61115
rect 6929 61081 6963 61115
rect 7849 61081 7883 61115
rect 15209 61081 15243 61115
rect 16313 61081 16347 61115
rect 18889 61081 18923 61115
rect 19993 61081 20027 61115
rect 22753 61081 22787 61115
rect 24041 61081 24075 61115
rect 26433 61081 26467 61115
rect 34253 61081 34287 61115
rect 34989 61081 35023 61115
rect 35909 61081 35943 61115
rect 37749 61081 37783 61115
rect 40877 61081 40911 61115
rect 42901 61081 42935 61115
rect 55781 61081 55815 61115
rect 5181 61013 5215 61047
rect 5917 61013 5951 61047
rect 11069 61013 11103 61047
rect 12173 61013 12207 61047
rect 17325 61013 17359 61047
rect 21373 61013 21407 61047
rect 25421 61013 25455 61047
rect 27353 61013 27387 61047
rect 28365 61013 28399 61047
rect 29929 61013 29963 61047
rect 31309 61013 31343 61047
rect 32505 61013 32539 61047
rect 33425 61013 33459 61047
rect 35081 61013 35115 61047
rect 36553 61013 36587 61047
rect 39129 61013 39163 61047
rect 40969 61013 41003 61047
rect 41705 61013 41739 61047
rect 44465 61013 44499 61047
rect 45385 61013 45419 61047
rect 46121 61013 46155 61047
rect 48697 61013 48731 61047
rect 50537 61013 50571 61047
rect 54309 61013 54343 61047
rect 56609 61013 56643 61047
rect 58265 61013 58299 61047
rect 3249 60741 3283 60775
rect 3985 60741 4019 60775
rect 8401 60741 8435 60775
rect 13553 60741 13587 60775
rect 14289 60741 14323 60775
rect 15761 60741 15795 60775
rect 19441 60741 19475 60775
rect 24593 60741 24627 60775
rect 27537 60741 27571 60775
rect 29009 60741 29043 60775
rect 30481 60741 30515 60775
rect 36369 60741 36403 60775
rect 41521 60741 41555 60775
rect 46673 60741 46707 60775
rect 50353 60741 50387 60775
rect 53021 60741 53055 60775
rect 1593 60673 1627 60707
rect 9045 60673 9079 60707
rect 22109 60673 22143 60707
rect 22293 60673 22327 60707
rect 22385 60673 22419 60707
rect 22529 60673 22563 60707
rect 23213 60673 23247 60707
rect 54677 60673 54711 60707
rect 55413 60673 55447 60707
rect 56149 60673 56183 60707
rect 56885 60673 56919 60707
rect 58081 60673 58115 60707
rect 1869 60605 1903 60639
rect 4169 60537 4203 60571
rect 8585 60537 8619 60571
rect 19625 60537 19659 60571
rect 56333 60537 56367 60571
rect 3341 60469 3375 60503
rect 9229 60469 9263 60503
rect 13645 60469 13679 60503
rect 14381 60469 14415 60503
rect 15853 60469 15887 60503
rect 22661 60469 22695 60503
rect 23397 60469 23431 60503
rect 24685 60469 24719 60503
rect 27629 60469 27663 60503
rect 29101 60469 29135 60503
rect 30573 60469 30607 60503
rect 36461 60469 36495 60503
rect 41613 60469 41647 60503
rect 46765 60469 46799 60503
rect 50445 60469 50479 60503
rect 53113 60469 53147 60503
rect 54861 60469 54895 60503
rect 55597 60469 55631 60503
rect 57069 60469 57103 60503
rect 58265 60469 58299 60503
rect 21005 60197 21039 60231
rect 41153 60197 41187 60231
rect 17877 60129 17911 60163
rect 42625 60129 42659 60163
rect 57437 60129 57471 60163
rect 2605 60061 2639 60095
rect 7389 60061 7423 60095
rect 7665 60061 7699 60095
rect 7757 60061 7791 60095
rect 18061 60061 18095 60095
rect 18429 60061 18463 60095
rect 18613 60061 18647 60095
rect 20453 60061 20487 60095
rect 20637 60061 20671 60095
rect 20729 60061 20763 60095
rect 20873 60061 20907 60095
rect 22017 60061 22051 60095
rect 22109 60061 22143 60095
rect 22385 60061 22419 60095
rect 22661 60061 22695 60095
rect 22845 60061 22879 60095
rect 23489 60061 23523 60095
rect 23765 60061 23799 60095
rect 23857 60061 23891 60095
rect 28089 60061 28123 60095
rect 28182 60061 28216 60095
rect 28457 60061 28491 60095
rect 28554 60061 28588 60095
rect 30113 60061 30147 60095
rect 30389 60061 30423 60095
rect 30482 60061 30516 60095
rect 30895 60061 30929 60095
rect 32505 60061 32539 60095
rect 32689 60061 32723 60095
rect 33057 60061 33091 60095
rect 33241 60061 33275 60095
rect 40601 60061 40635 60095
rect 40877 60061 40911 60095
rect 40974 60061 41008 60095
rect 42165 60061 42199 60095
rect 42349 60061 42383 60095
rect 42717 60061 42751 60095
rect 56517 60061 56551 60095
rect 57253 60061 57287 60095
rect 57897 60061 57931 60095
rect 1685 59993 1719 60027
rect 2053 59993 2087 60027
rect 7573 59993 7607 60027
rect 23673 59993 23707 60027
rect 28365 59993 28399 60027
rect 30665 59993 30699 60027
rect 30757 59993 30791 60027
rect 40785 59993 40819 60027
rect 58173 59993 58207 60027
rect 2697 59925 2731 59959
rect 7941 59925 7975 59959
rect 17509 59925 17543 59959
rect 21649 59925 21683 59959
rect 24041 59925 24075 59959
rect 28733 59925 28767 59959
rect 31033 59925 31067 59959
rect 32321 59925 32355 59959
rect 41981 59925 42015 59959
rect 56609 59925 56643 59959
rect 58265 59721 58299 59755
rect 2605 59653 2639 59687
rect 21005 59653 21039 59687
rect 23397 59653 23431 59687
rect 30113 59653 30147 59687
rect 57345 59653 57379 59687
rect 1685 59585 1719 59619
rect 19349 59585 19383 59619
rect 19533 59585 19567 59619
rect 19625 59585 19659 59619
rect 19769 59585 19803 59619
rect 20821 59585 20855 59619
rect 21097 59585 21131 59619
rect 21189 59585 21223 59619
rect 22109 59585 22143 59619
rect 22661 59585 22695 59619
rect 23213 59585 23247 59619
rect 23489 59585 23523 59619
rect 23633 59585 23667 59619
rect 28365 59585 28399 59619
rect 29745 59585 29779 59619
rect 29838 59585 29872 59619
rect 30021 59585 30055 59619
rect 30210 59585 30244 59619
rect 43269 59585 43303 59619
rect 43637 59585 43671 59619
rect 58081 59585 58115 59619
rect 28549 59517 28583 59551
rect 42717 59517 42751 59551
rect 43085 59517 43119 59551
rect 43545 59517 43579 59551
rect 21373 59449 21407 59483
rect 57529 59449 57563 59483
rect 1961 59381 1995 59415
rect 2697 59381 2731 59415
rect 19901 59381 19935 59415
rect 23765 59381 23799 59415
rect 29469 59381 29503 59415
rect 30389 59381 30423 59415
rect 30757 59381 30791 59415
rect 57345 59177 57379 59211
rect 19993 59109 20027 59143
rect 41337 59041 41371 59075
rect 41797 59041 41831 59075
rect 58081 59041 58115 59075
rect 1685 58973 1719 59007
rect 19441 58973 19475 59007
rect 19717 58973 19751 59007
rect 19861 58973 19895 59007
rect 41521 58973 41555 59007
rect 41889 58973 41923 59007
rect 57161 58973 57195 59007
rect 57897 58973 57931 59007
rect 19625 58905 19659 58939
rect 1777 58837 1811 58871
rect 41153 58837 41187 58871
rect 58173 58565 58207 58599
rect 1593 58497 1627 58531
rect 37933 58497 37967 58531
rect 38025 58497 38059 58531
rect 38301 58497 38335 58531
rect 38577 58497 38611 58531
rect 38853 58497 38887 58531
rect 41337 58497 41371 58531
rect 41521 58497 41555 58531
rect 41889 58497 41923 58531
rect 1869 58429 1903 58463
rect 41797 58429 41831 58463
rect 37565 58293 37599 58327
rect 41153 58293 41187 58327
rect 58265 58293 58299 58327
rect 1593 57885 1627 57919
rect 35633 57885 35667 57919
rect 35909 57885 35943 57919
rect 36001 57885 36035 57919
rect 36277 57885 36311 57919
rect 36553 57885 36587 57919
rect 1869 57817 1903 57851
rect 35173 57817 35207 57851
rect 57989 57817 58023 57851
rect 58081 57749 58115 57783
rect 1593 57409 1627 57443
rect 35725 57409 35759 57443
rect 36001 57341 36035 57375
rect 1777 57205 1811 57239
rect 32873 56865 32907 56899
rect 33333 56865 33367 56899
rect 33057 56797 33091 56831
rect 33425 56797 33459 56831
rect 57897 56797 57931 56831
rect 1685 56729 1719 56763
rect 2053 56729 2087 56763
rect 58173 56729 58207 56763
rect 32505 56661 32539 56695
rect 58173 56389 58207 56423
rect 24409 56321 24443 56355
rect 24777 56321 24811 56355
rect 24869 56321 24903 56355
rect 29469 56321 29503 56355
rect 29837 56321 29871 56355
rect 41337 56321 41371 56355
rect 41521 56321 41555 56355
rect 41889 56321 41923 56355
rect 24317 56253 24351 56287
rect 29561 56253 29595 56287
rect 29929 56253 29963 56287
rect 41797 56253 41831 56287
rect 23857 56117 23891 56151
rect 28917 56117 28951 56151
rect 41153 56117 41187 56151
rect 58265 56117 58299 56151
rect 58357 55913 58391 55947
rect 25237 55709 25271 55743
rect 25329 55709 25363 55743
rect 25605 55709 25639 55743
rect 25697 55709 25731 55743
rect 1685 55641 1719 55675
rect 24593 55641 24627 55675
rect 1777 55573 1811 55607
rect 1777 55369 1811 55403
rect 41061 55301 41095 55335
rect 41153 55301 41187 55335
rect 1593 55233 1627 55267
rect 40877 55233 40911 55267
rect 41250 55233 41284 55267
rect 41446 55233 41480 55267
rect 23397 54689 23431 54723
rect 23489 54621 23523 54655
rect 23857 54621 23891 54655
rect 24041 54621 24075 54655
rect 58357 54621 58391 54655
rect 1685 54553 1719 54587
rect 22845 54553 22879 54587
rect 1777 54485 1811 54519
rect 1593 54145 1627 54179
rect 1777 53941 1811 53975
rect 40877 53669 40911 53703
rect 41337 53601 41371 53635
rect 40325 53533 40359 53567
rect 40745 53533 40779 53567
rect 40509 53465 40543 53499
rect 40601 53465 40635 53499
rect 23765 53125 23799 53159
rect 23857 53125 23891 53159
rect 1685 53057 1719 53091
rect 23581 53057 23615 53091
rect 23949 53057 23983 53091
rect 24593 53057 24627 53091
rect 24777 52989 24811 53023
rect 1777 52853 1811 52887
rect 24133 52853 24167 52887
rect 58357 52853 58391 52887
rect 24961 52649 24995 52683
rect 1869 52513 1903 52547
rect 1593 52445 1627 52479
rect 24685 52377 24719 52411
rect 1869 52037 1903 52071
rect 8217 52037 8251 52071
rect 1685 51969 1719 52003
rect 8033 51969 8067 52003
rect 8309 51969 8343 52003
rect 7849 51765 7883 51799
rect 20821 51561 20855 51595
rect 21005 51493 21039 51527
rect 20913 51425 20947 51459
rect 21097 51357 21131 51391
rect 21281 51357 21315 51391
rect 58357 51357 58391 51391
rect 1685 51289 1719 51323
rect 1869 51289 1903 51323
rect 20545 51221 20579 51255
rect 3985 50949 4019 50983
rect 3709 50881 3743 50915
rect 3893 50881 3927 50915
rect 4082 50881 4116 50915
rect 4261 50677 4295 50711
rect 57897 50269 57931 50303
rect 1685 50201 1719 50235
rect 1869 50201 1903 50235
rect 58173 50201 58207 50235
rect 1593 49793 1627 49827
rect 1777 49657 1811 49691
rect 1593 49181 1627 49215
rect 57989 49113 58023 49147
rect 58357 49113 58391 49147
rect 1777 49045 1811 49079
rect 1685 48705 1719 48739
rect 1869 48569 1903 48603
rect 2605 48229 2639 48263
rect 2053 48093 2087 48127
rect 2237 48093 2271 48127
rect 2426 48093 2460 48127
rect 57897 48093 57931 48127
rect 2329 48025 2363 48059
rect 58173 48025 58207 48059
rect 1685 47617 1719 47651
rect 58081 47617 58115 47651
rect 1869 47481 1903 47515
rect 58265 47413 58299 47447
rect 1593 47005 1627 47039
rect 1777 46869 1811 46903
rect 1593 46529 1627 46563
rect 1777 46325 1811 46359
rect 58173 45985 58207 46019
rect 57897 45917 57931 45951
rect 1685 45849 1719 45883
rect 1777 45781 1811 45815
rect 36553 45509 36587 45543
rect 38209 45509 38243 45543
rect 38301 45509 38335 45543
rect 17049 45441 17083 45475
rect 17142 45441 17176 45475
rect 17325 45441 17359 45475
rect 17414 45441 17448 45475
rect 17555 45441 17589 45475
rect 36369 45441 36403 45475
rect 36645 45441 36679 45475
rect 36783 45441 36817 45475
rect 37749 45441 37783 45475
rect 38025 45441 38059 45475
rect 38398 45441 38432 45475
rect 58081 45441 58115 45475
rect 36921 45305 36955 45339
rect 38577 45305 38611 45339
rect 17693 45237 17727 45271
rect 58265 45237 58299 45271
rect 1593 44829 1627 44863
rect 56977 44829 57011 44863
rect 1869 44761 1903 44795
rect 57253 44761 57287 44795
rect 57989 44761 58023 44795
rect 58357 44761 58391 44795
rect 34345 44421 34379 44455
rect 1685 44353 1719 44387
rect 34069 44353 34103 44387
rect 34253 44353 34287 44387
rect 34442 44353 34476 44387
rect 1869 44217 1903 44251
rect 34621 44217 34655 44251
rect 34253 43877 34287 43911
rect 33701 43741 33735 43775
rect 34074 43741 34108 43775
rect 57897 43741 57931 43775
rect 1685 43673 1719 43707
rect 33885 43673 33919 43707
rect 33977 43673 34011 43707
rect 58173 43673 58207 43707
rect 1777 43605 1811 43639
rect 32505 43333 32539 43367
rect 32597 43333 32631 43367
rect 1593 43265 1627 43299
rect 32321 43265 32355 43299
rect 32741 43265 32775 43299
rect 1777 43061 1811 43095
rect 32873 43061 32907 43095
rect 33057 42653 33091 42687
rect 33149 42653 33183 42687
rect 33425 42653 33459 42687
rect 33701 42653 33735 42687
rect 33885 42653 33919 42687
rect 37289 42653 37323 42687
rect 37657 42653 37691 42687
rect 37473 42585 37507 42619
rect 37565 42585 37599 42619
rect 57069 42585 57103 42619
rect 57989 42585 58023 42619
rect 58357 42585 58391 42619
rect 32689 42517 32723 42551
rect 37841 42517 37875 42551
rect 57345 42517 57379 42551
rect 1593 42177 1627 42211
rect 1777 41973 1811 42007
rect 56977 41565 57011 41599
rect 1685 41497 1719 41531
rect 57253 41497 57287 41531
rect 57989 41497 58023 41531
rect 58357 41497 58391 41531
rect 1961 41429 1995 41463
rect 1685 41089 1719 41123
rect 1777 40885 1811 40919
rect 57897 40477 57931 40511
rect 1685 40409 1719 40443
rect 57069 40409 57103 40443
rect 58173 40409 58207 40443
rect 1777 40341 1811 40375
rect 57161 40341 57195 40375
rect 21189 40069 21223 40103
rect 20913 40001 20947 40035
rect 21097 40001 21131 40035
rect 21281 40001 21315 40035
rect 21465 39797 21499 39831
rect 2881 39525 2915 39559
rect 1869 39457 1903 39491
rect 2329 39389 2363 39423
rect 2605 39389 2639 39423
rect 2749 39389 2783 39423
rect 1685 39321 1719 39355
rect 2513 39321 2547 39355
rect 57069 39321 57103 39355
rect 57989 39321 58023 39355
rect 57161 39253 57195 39287
rect 58081 39253 58115 39287
rect 23302 38981 23336 39015
rect 1685 38913 1719 38947
rect 22937 38913 22971 38947
rect 23085 38913 23119 38947
rect 23213 38913 23247 38947
rect 23402 38913 23436 38947
rect 1869 38777 1903 38811
rect 23581 38709 23615 38743
rect 1777 38505 1811 38539
rect 20177 38505 20211 38539
rect 2605 38369 2639 38403
rect 21189 38369 21223 38403
rect 21557 38369 21591 38403
rect 2789 38301 2823 38335
rect 20177 38301 20211 38335
rect 20361 38301 20395 38335
rect 20453 38301 20487 38335
rect 21465 38301 21499 38335
rect 21741 38301 21775 38335
rect 23121 38301 23155 38335
rect 57897 38301 57931 38335
rect 1685 38233 1719 38267
rect 2973 38233 3007 38267
rect 23489 38233 23523 38267
rect 58173 38233 58207 38267
rect 20637 38165 20671 38199
rect 21925 38165 21959 38199
rect 23305 37961 23339 37995
rect 2237 37893 2271 37927
rect 21005 37893 21039 37927
rect 22937 37893 22971 37927
rect 23765 37893 23799 37927
rect 25237 37893 25271 37927
rect 2053 37825 2087 37859
rect 2329 37825 2363 37859
rect 2421 37825 2455 37859
rect 19349 37825 19383 37859
rect 19497 37825 19531 37859
rect 19625 37825 19659 37859
rect 19717 37825 19751 37859
rect 19855 37825 19889 37859
rect 20361 37825 20395 37859
rect 20821 37825 20855 37859
rect 21097 37825 21131 37859
rect 22753 37825 22787 37859
rect 23029 37825 23063 37859
rect 23121 37825 23155 37859
rect 24961 37825 24995 37859
rect 25099 37825 25133 37859
rect 25329 37825 25363 37859
rect 58081 37825 58115 37859
rect 22477 37757 22511 37791
rect 24133 37757 24167 37791
rect 19993 37689 20027 37723
rect 24041 37689 24075 37723
rect 25513 37689 25547 37723
rect 2605 37621 2639 37655
rect 20637 37621 20671 37655
rect 23930 37621 23964 37655
rect 24409 37621 24443 37655
rect 58265 37621 58299 37655
rect 1869 37281 1903 37315
rect 21097 37281 21131 37315
rect 1685 37213 1719 37247
rect 5917 37213 5951 37247
rect 6009 37213 6043 37247
rect 6285 37213 6319 37247
rect 6561 37213 6595 37247
rect 6745 37213 6779 37247
rect 19625 37213 19659 37247
rect 20913 37213 20947 37247
rect 53849 37213 53883 37247
rect 54125 37213 54159 37247
rect 54269 37213 54303 37247
rect 57897 37213 57931 37247
rect 19993 37145 20027 37179
rect 54033 37145 54067 37179
rect 58173 37145 58207 37179
rect 5549 37077 5583 37111
rect 54409 37077 54443 37111
rect 18705 36805 18739 36839
rect 53941 36805 53975 36839
rect 1593 36737 1627 36771
rect 18429 36737 18463 36771
rect 18613 36737 18647 36771
rect 18797 36737 18831 36771
rect 19441 36737 19475 36771
rect 23489 36737 23523 36771
rect 23765 36737 23799 36771
rect 24041 36737 24075 36771
rect 53665 36737 53699 36771
rect 53849 36737 53883 36771
rect 54038 36737 54072 36771
rect 23857 36669 23891 36703
rect 20729 36601 20763 36635
rect 54217 36601 54251 36635
rect 1777 36533 1811 36567
rect 18981 36533 19015 36567
rect 23765 36533 23799 36567
rect 24225 36533 24259 36567
rect 1777 36329 1811 36363
rect 3065 36329 3099 36363
rect 23857 36329 23891 36363
rect 20269 36261 20303 36295
rect 20729 36193 20763 36227
rect 2513 36125 2547 36159
rect 2886 36125 2920 36159
rect 20177 36125 20211 36159
rect 20453 36125 20487 36159
rect 22201 36125 22235 36159
rect 22477 36125 22511 36159
rect 22569 36125 22603 36159
rect 23305 36125 23339 36159
rect 23673 36125 23707 36159
rect 24593 36125 24627 36159
rect 24777 36125 24811 36159
rect 1685 36057 1719 36091
rect 2697 36057 2731 36091
rect 2789 36057 2823 36091
rect 22385 36057 22419 36091
rect 23489 36057 23523 36091
rect 23581 36057 23615 36091
rect 25145 36057 25179 36091
rect 57989 36057 58023 36091
rect 58357 36057 58391 36091
rect 22753 35989 22787 36023
rect 1777 35785 1811 35819
rect 20453 35785 20487 35819
rect 40785 35785 40819 35819
rect 19257 35717 19291 35751
rect 40417 35717 40451 35751
rect 1685 35649 1719 35683
rect 19073 35649 19107 35683
rect 19349 35649 19383 35683
rect 19441 35649 19475 35683
rect 20085 35649 20119 35683
rect 22661 35649 22695 35683
rect 40233 35649 40267 35683
rect 40509 35649 40543 35683
rect 40601 35649 40635 35683
rect 20177 35581 20211 35615
rect 23397 35581 23431 35615
rect 19625 35513 19659 35547
rect 20085 35445 20119 35479
rect 22753 35241 22787 35275
rect 40601 35241 40635 35275
rect 1869 35173 1903 35207
rect 22753 35105 22787 35139
rect 22569 35037 22603 35071
rect 22845 35037 22879 35071
rect 40049 35037 40083 35071
rect 40325 35037 40359 35071
rect 40417 35037 40451 35071
rect 57897 35037 57931 35071
rect 1685 34969 1719 35003
rect 40233 34969 40267 35003
rect 58173 34969 58207 35003
rect 23029 34901 23063 34935
rect 58265 34697 58299 34731
rect 58081 34561 58115 34595
rect 21373 33949 21407 33983
rect 21521 33949 21555 33983
rect 21838 33949 21872 33983
rect 22569 33949 22603 33983
rect 23029 33949 23063 33983
rect 24593 33949 24627 33983
rect 24741 33949 24775 33983
rect 25099 33949 25133 33983
rect 1685 33881 1719 33915
rect 21649 33881 21683 33915
rect 21761 33881 21795 33915
rect 23305 33881 23339 33915
rect 24869 33881 24903 33915
rect 24961 33881 24995 33915
rect 1777 33813 1811 33847
rect 22017 33813 22051 33847
rect 25237 33813 25271 33847
rect 1869 33541 1903 33575
rect 21189 33541 21223 33575
rect 36093 33541 36127 33575
rect 1685 33473 1719 33507
rect 20637 33473 20671 33507
rect 20913 33473 20947 33507
rect 21097 33473 21131 33507
rect 21281 33473 21315 33507
rect 22017 33473 22051 33507
rect 22165 33473 22199 33507
rect 22293 33473 22327 33507
rect 22385 33473 22419 33507
rect 22523 33473 22557 33507
rect 35725 33473 35759 33507
rect 35818 33473 35852 33507
rect 36001 33473 36035 33507
rect 36190 33473 36224 33507
rect 21465 33337 21499 33371
rect 22661 33269 22695 33303
rect 36369 33269 36403 33303
rect 21925 32997 21959 33031
rect 24869 32997 24903 33031
rect 58173 32929 58207 32963
rect 21833 32861 21867 32895
rect 22109 32861 22143 32895
rect 24777 32861 24811 32895
rect 25053 32861 25087 32895
rect 57897 32861 57931 32895
rect 1685 32793 1719 32827
rect 57069 32793 57103 32827
rect 1777 32725 1811 32759
rect 22293 32725 22327 32759
rect 25237 32725 25271 32759
rect 57161 32725 57195 32759
rect 1685 32385 1719 32419
rect 1777 32181 1811 32215
rect 22477 31841 22511 31875
rect 22753 31773 22787 31807
rect 23029 31773 23063 31807
rect 23121 31773 23155 31807
rect 57897 31773 57931 31807
rect 58173 31773 58207 31807
rect 22937 31705 22971 31739
rect 23305 31637 23339 31671
rect 1685 31297 1719 31331
rect 24133 31297 24167 31331
rect 24226 31297 24260 31331
rect 24409 31297 24443 31331
rect 24501 31297 24535 31331
rect 24617 31297 24651 31331
rect 58081 31297 58115 31331
rect 24777 31161 24811 31195
rect 1777 31093 1811 31127
rect 58265 31093 58299 31127
rect 23213 30889 23247 30923
rect 19533 30753 19567 30787
rect 19441 30685 19475 30719
rect 19717 30685 19751 30719
rect 23121 30685 23155 30719
rect 23305 30685 23339 30719
rect 23581 30685 23615 30719
rect 1685 30617 1719 30651
rect 20177 30617 20211 30651
rect 22845 30617 22879 30651
rect 1777 30549 1811 30583
rect 22569 30549 22603 30583
rect 23489 30549 23523 30583
rect 19349 30345 19383 30379
rect 19073 30277 19107 30311
rect 1593 30209 1627 30243
rect 18705 30209 18739 30243
rect 18853 30209 18887 30243
rect 18981 30209 19015 30243
rect 19211 30209 19245 30243
rect 22293 30209 22327 30243
rect 22569 30209 22603 30243
rect 1777 30141 1811 30175
rect 22385 30141 22419 30175
rect 22753 30141 22787 30175
rect 22109 29801 22143 29835
rect 23121 29801 23155 29835
rect 58173 29665 58207 29699
rect 1593 29597 1627 29631
rect 21557 29597 21591 29631
rect 21925 29597 21959 29631
rect 22569 29597 22603 29631
rect 22845 29597 22879 29631
rect 22937 29597 22971 29631
rect 57897 29597 57931 29631
rect 1869 29529 1903 29563
rect 21741 29529 21775 29563
rect 21833 29529 21867 29563
rect 22753 29529 22787 29563
rect 57069 29529 57103 29563
rect 57161 29461 57195 29495
rect 9689 29257 9723 29291
rect 9321 29121 9355 29155
rect 9475 29121 9509 29155
rect 2881 28577 2915 28611
rect 1593 28509 1627 28543
rect 2513 28509 2547 28543
rect 2667 28509 2701 28543
rect 57897 28509 57931 28543
rect 1869 28441 1903 28475
rect 58173 28441 58207 28475
rect 23305 28101 23339 28135
rect 1593 28033 1627 28067
rect 23121 28033 23155 28067
rect 23397 28033 23431 28067
rect 23489 28033 23523 28067
rect 1777 27965 1811 27999
rect 23673 27829 23707 27863
rect 1593 27421 1627 27455
rect 23121 27421 23155 27455
rect 23269 27421 23303 27455
rect 23586 27421 23620 27455
rect 57989 27421 58023 27455
rect 1869 27353 1903 27387
rect 23397 27353 23431 27387
rect 23489 27353 23523 27387
rect 23765 27285 23799 27319
rect 58081 27285 58115 27319
rect 2881 27081 2915 27115
rect 1593 26945 1627 26979
rect 2513 26945 2547 26979
rect 2606 26945 2640 26979
rect 22753 26945 22787 26979
rect 22845 26945 22879 26979
rect 23029 26945 23063 26979
rect 1777 26877 1811 26911
rect 23397 26877 23431 26911
rect 58173 26401 58207 26435
rect 57897 26333 57931 26367
rect 1593 25857 1627 25891
rect 10701 25857 10735 25891
rect 10855 25857 10889 25891
rect 58081 25857 58115 25891
rect 1777 25789 1811 25823
rect 10885 25653 10919 25687
rect 58265 25653 58299 25687
rect 2881 25313 2915 25347
rect 1593 25245 1627 25279
rect 2513 25245 2547 25279
rect 2606 25245 2640 25279
rect 57897 25245 57931 25279
rect 1869 25177 1903 25211
rect 58173 25177 58207 25211
rect 1593 24769 1627 24803
rect 58081 24769 58115 24803
rect 1777 24701 1811 24735
rect 58265 24565 58299 24599
rect 3065 24361 3099 24395
rect 1593 24157 1627 24191
rect 2881 24157 2915 24191
rect 3035 24157 3069 24191
rect 1869 24089 1903 24123
rect 12817 23749 12851 23783
rect 12265 23681 12299 23715
rect 12173 23273 12207 23307
rect 18245 23205 18279 23239
rect 58173 23137 58207 23171
rect 1593 23069 1627 23103
rect 10885 23069 10919 23103
rect 11039 23069 11073 23103
rect 11989 23069 12023 23103
rect 12143 23069 12177 23103
rect 18521 23069 18555 23103
rect 57897 23069 57931 23103
rect 1869 23001 1903 23035
rect 11253 23001 11287 23035
rect 18245 23001 18279 23035
rect 18429 22933 18463 22967
rect 18429 22661 18463 22695
rect 19441 22661 19475 22695
rect 19641 22661 19675 22695
rect 58173 22661 58207 22695
rect 1593 22593 1627 22627
rect 17049 22593 17083 22627
rect 18153 22593 18187 22627
rect 18245 22593 18279 22627
rect 25973 22593 26007 22627
rect 1777 22525 1811 22559
rect 16957 22525 16991 22559
rect 25789 22525 25823 22559
rect 19809 22457 19843 22491
rect 17417 22389 17451 22423
rect 19625 22389 19659 22423
rect 26157 22389 26191 22423
rect 58265 22389 58299 22423
rect 9689 22185 9723 22219
rect 26157 22049 26191 22083
rect 1593 21981 1627 22015
rect 9505 21981 9539 22015
rect 9659 21981 9693 22015
rect 16589 21981 16623 22015
rect 21005 21981 21039 22015
rect 21189 21981 21223 22015
rect 57897 21981 57931 22015
rect 1869 21913 1903 21947
rect 19625 21913 19659 21947
rect 19901 21913 19935 21947
rect 19993 21913 20027 21947
rect 58173 21913 58207 21947
rect 17785 21845 17819 21879
rect 19809 21845 19843 21879
rect 20177 21845 20211 21879
rect 21373 21845 21407 21879
rect 25605 21845 25639 21879
rect 25973 21845 26007 21879
rect 26065 21845 26099 21879
rect 12081 21641 12115 21675
rect 22017 21641 22051 21675
rect 22385 21641 22419 21675
rect 24961 21641 24995 21675
rect 29837 21641 29871 21675
rect 1685 21505 1719 21539
rect 11713 21505 11747 21539
rect 11867 21505 11901 21539
rect 13001 21505 13035 21539
rect 13093 21505 13127 21539
rect 13277 21505 13311 21539
rect 15215 21505 15249 21539
rect 15393 21505 15427 21539
rect 16129 21505 16163 21539
rect 16313 21505 16347 21539
rect 17224 21505 17258 21539
rect 18797 21505 18831 21539
rect 23581 21505 23615 21539
rect 27813 21505 27847 21539
rect 28641 21505 28675 21539
rect 36001 21505 36035 21539
rect 38669 21505 38703 21539
rect 58081 21505 58115 21539
rect 13185 21437 13219 21471
rect 16957 21437 16991 21471
rect 22477 21437 22511 21471
rect 22661 21437 22695 21471
rect 27905 21437 27939 21471
rect 27997 21437 28031 21471
rect 36093 21437 36127 21471
rect 36277 21437 36311 21471
rect 38761 21437 38795 21471
rect 38853 21437 38887 21471
rect 18337 21369 18371 21403
rect 1777 21301 1811 21335
rect 12817 21301 12851 21335
rect 15209 21301 15243 21335
rect 16129 21301 16163 21335
rect 19993 21301 20027 21335
rect 27445 21301 27479 21335
rect 28549 21301 28583 21335
rect 35265 21301 35299 21335
rect 35633 21301 35667 21335
rect 37933 21301 37967 21335
rect 38301 21301 38335 21335
rect 58265 21301 58299 21335
rect 15945 21097 15979 21131
rect 19993 21097 20027 21131
rect 19441 21029 19475 21063
rect 27353 21029 27387 21063
rect 30665 21029 30699 21063
rect 53297 21029 53331 21063
rect 11713 20961 11747 20995
rect 12173 20961 12207 20995
rect 17969 20961 18003 20995
rect 22017 20961 22051 20995
rect 27813 20961 27847 20995
rect 27997 20961 28031 20995
rect 31217 20961 31251 20995
rect 36001 20961 36035 20995
rect 38301 20961 38335 20995
rect 42073 20961 42107 20995
rect 54125 20961 54159 20995
rect 54585 20961 54619 20995
rect 55597 20961 55631 20995
rect 11805 20893 11839 20927
rect 12817 20893 12851 20927
rect 13001 20893 13035 20927
rect 15301 20893 15335 20927
rect 15485 20893 15519 20927
rect 15945 20893 15979 20927
rect 16129 20893 16163 20927
rect 16589 20893 16623 20927
rect 19809 20893 19843 20927
rect 20913 20893 20947 20927
rect 23673 20893 23707 20927
rect 23857 20893 23891 20927
rect 24593 20893 24627 20927
rect 26433 20893 26467 20927
rect 26525 20893 26559 20927
rect 27721 20893 27755 20927
rect 28641 20893 28675 20927
rect 28733 20893 28767 20927
rect 29837 20893 29871 20927
rect 30021 20893 30055 20927
rect 34897 20893 34931 20927
rect 38485 20893 38519 20927
rect 42717 20893 42751 20927
rect 42901 20893 42935 20927
rect 43913 20893 43947 20927
rect 47501 20893 47535 20927
rect 47869 20893 47903 20927
rect 52745 20893 52779 20927
rect 53113 20893 53147 20927
rect 53757 20893 53791 20927
rect 53941 20893 53975 20927
rect 54769 20893 54803 20927
rect 55781 20893 55815 20927
rect 57897 20893 57931 20927
rect 12633 20825 12667 20859
rect 24041 20825 24075 20859
rect 24838 20825 24872 20859
rect 27077 20825 27111 20859
rect 41889 20825 41923 20859
rect 43545 20825 43579 20859
rect 43729 20825 43763 20859
rect 47685 20825 47719 20859
rect 47777 20825 47811 20859
rect 52929 20825 52963 20859
rect 53021 20825 53055 20859
rect 58173 20825 58207 20859
rect 12909 20757 12943 20791
rect 13185 20757 13219 20791
rect 15393 20757 15427 20791
rect 19625 20757 19659 20791
rect 19717 20757 19751 20791
rect 25973 20757 26007 20791
rect 26709 20757 26743 20791
rect 28917 20757 28951 20791
rect 30205 20757 30239 20791
rect 31033 20757 31067 20791
rect 31125 20757 31159 20791
rect 38669 20757 38703 20791
rect 41521 20757 41555 20791
rect 41981 20757 42015 20791
rect 43085 20757 43119 20791
rect 48053 20757 48087 20791
rect 54953 20757 54987 20791
rect 55965 20757 55999 20791
rect 19717 20553 19751 20587
rect 25513 20553 25547 20587
rect 28549 20553 28583 20587
rect 44097 20553 44131 20587
rect 49525 20553 49559 20587
rect 54493 20553 54527 20587
rect 56333 20553 56367 20587
rect 22262 20485 22296 20519
rect 27414 20485 27448 20519
rect 42984 20485 43018 20519
rect 46029 20485 46063 20519
rect 1593 20417 1627 20451
rect 8033 20417 8067 20451
rect 10977 20417 11011 20451
rect 11161 20417 11195 20451
rect 12440 20417 12474 20451
rect 14013 20417 14047 20451
rect 17601 20417 17635 20451
rect 17877 20417 17911 20451
rect 18061 20417 18095 20451
rect 18521 20417 18555 20451
rect 21281 20417 21315 20451
rect 21465 20417 21499 20451
rect 24317 20417 24351 20451
rect 27169 20417 27203 20451
rect 29469 20417 29503 20451
rect 33517 20417 33551 20451
rect 37657 20417 37691 20451
rect 38393 20417 38427 20451
rect 41429 20417 41463 20451
rect 47041 20417 47075 20451
rect 48412 20417 48446 20451
rect 50261 20417 50295 20451
rect 50528 20417 50562 20451
rect 53113 20417 53147 20451
rect 53380 20417 53414 20451
rect 54953 20417 54987 20451
rect 55220 20417 55254 20451
rect 1777 20349 1811 20383
rect 12173 20349 12207 20383
rect 22017 20349 22051 20383
rect 33333 20349 33367 20383
rect 35173 20349 35207 20383
rect 35449 20349 35483 20383
rect 37473 20349 37507 20383
rect 38669 20349 38703 20383
rect 41245 20349 41279 20383
rect 42717 20349 42751 20383
rect 46857 20349 46891 20383
rect 48145 20349 48179 20383
rect 13553 20281 13587 20315
rect 30665 20281 30699 20315
rect 46305 20281 46339 20315
rect 51641 20281 51675 20315
rect 9413 20213 9447 20247
rect 11069 20213 11103 20247
rect 15209 20213 15243 20247
rect 17417 20213 17451 20247
rect 21281 20213 21315 20247
rect 23397 20213 23431 20247
rect 33701 20213 33735 20247
rect 36553 20213 36587 20247
rect 37841 20213 37875 20247
rect 39773 20213 39807 20247
rect 41613 20213 41647 20247
rect 47225 20213 47259 20247
rect 16037 20009 16071 20043
rect 20821 20009 20855 20043
rect 22753 20009 22787 20043
rect 31861 20009 31895 20043
rect 35357 20009 35391 20043
rect 54401 20009 54435 20043
rect 56057 20009 56091 20043
rect 9413 19941 9447 19975
rect 37749 19941 37783 19975
rect 42533 19941 42567 19975
rect 44465 19941 44499 19975
rect 48421 19941 48455 19975
rect 9597 19873 9631 19907
rect 10241 19873 10275 19907
rect 13185 19873 13219 19907
rect 25605 19873 25639 19907
rect 27629 19873 27663 19907
rect 34989 19873 35023 19907
rect 38301 19873 38335 19907
rect 51457 19873 51491 19907
rect 56609 19873 56643 19907
rect 1593 19805 1627 19839
rect 6285 19805 6319 19839
rect 10333 19805 10367 19839
rect 11437 19805 11471 19839
rect 14657 19805 14691 19839
rect 14924 19805 14958 19839
rect 16589 19805 16623 19839
rect 19441 19805 19475 19839
rect 21557 19805 21591 19839
rect 24869 19805 24903 19839
rect 24961 19805 24995 19839
rect 25145 19805 25179 19839
rect 26341 19805 26375 19839
rect 29745 19805 29779 19839
rect 29929 19805 29963 19839
rect 30665 19805 30699 19839
rect 35173 19805 35207 19839
rect 35817 19805 35851 19839
rect 41153 19805 41187 19839
rect 43085 19805 43119 19839
rect 46121 19805 46155 19839
rect 46388 19805 46422 19839
rect 48053 19805 48087 19839
rect 48237 19805 48271 19839
rect 50353 19805 50387 19839
rect 50721 19805 50755 19839
rect 53849 19805 53883 19839
rect 54217 19805 54251 19839
rect 55505 19805 55539 19839
rect 55689 19805 55723 19839
rect 55873 19805 55907 19839
rect 56865 19805 56899 19839
rect 1869 19737 1903 19771
rect 9137 19737 9171 19771
rect 18889 19737 18923 19771
rect 19686 19737 19720 19771
rect 36084 19737 36118 19771
rect 40325 19737 40359 19771
rect 40509 19737 40543 19771
rect 41420 19737 41454 19771
rect 43330 19737 43364 19771
rect 45293 19737 45327 19771
rect 45661 19737 45695 19771
rect 50537 19737 50571 19771
rect 50629 19737 50663 19771
rect 51724 19737 51758 19771
rect 54033 19737 54067 19771
rect 54125 19737 54159 19771
rect 55781 19737 55815 19771
rect 7481 19669 7515 19703
rect 10701 19669 10735 19703
rect 30113 19669 30147 19703
rect 37197 19669 37231 19703
rect 38117 19669 38151 19703
rect 38209 19669 38243 19703
rect 40693 19669 40727 19703
rect 47501 19669 47535 19703
rect 50905 19669 50939 19703
rect 52837 19669 52871 19703
rect 57989 19669 58023 19703
rect 8217 19465 8251 19499
rect 13461 19465 13495 19499
rect 33885 19465 33919 19499
rect 34621 19465 34655 19499
rect 35081 19465 35115 19499
rect 36001 19465 36035 19499
rect 36369 19465 36403 19499
rect 36461 19465 36495 19499
rect 7104 19397 7138 19431
rect 18521 19397 18555 19431
rect 22652 19397 22686 19431
rect 32772 19397 32806 19431
rect 34989 19397 35023 19431
rect 42901 19397 42935 19431
rect 43821 19397 43855 19431
rect 51181 19397 51215 19431
rect 1593 19329 1627 19363
rect 1869 19329 1903 19363
rect 6837 19329 6871 19363
rect 8861 19329 8895 19363
rect 11897 19329 11931 19363
rect 14013 19329 14047 19363
rect 16865 19329 16899 19363
rect 19165 19329 19199 19363
rect 22385 19329 22419 19363
rect 24317 19329 24351 19363
rect 27169 19329 27203 19363
rect 30297 19329 30331 19363
rect 30553 19329 30587 19363
rect 32505 19329 32539 19363
rect 41889 19329 41923 19363
rect 42625 19329 42659 19363
rect 42809 19329 42843 19363
rect 42993 19329 43027 19363
rect 43131 19329 43165 19363
rect 45385 19329 45419 19363
rect 45652 19329 45686 19363
rect 47777 19329 47811 19363
rect 48053 19329 48087 19363
rect 50261 19329 50295 19363
rect 50905 19329 50939 19363
rect 51089 19329 51123 19363
rect 51273 19329 51307 19363
rect 52101 19329 52135 19363
rect 52285 19329 52319 19363
rect 12173 19261 12207 19295
rect 17141 19261 17175 19295
rect 20729 19261 20763 19295
rect 25421 19261 25455 19295
rect 34345 19261 34379 19295
rect 35265 19261 35299 19295
rect 36645 19261 36679 19295
rect 41705 19261 41739 19295
rect 43269 19261 43303 19295
rect 50077 19261 50111 19295
rect 51917 19261 51951 19295
rect 23765 19193 23799 19227
rect 31677 19193 31711 19227
rect 51457 19193 51491 19227
rect 2421 19125 2455 19159
rect 10057 19125 10091 19159
rect 15209 19125 15243 19159
rect 28365 19125 28399 19159
rect 35725 19125 35759 19159
rect 42073 19125 42107 19159
rect 43913 19125 43947 19159
rect 46765 19125 46799 19159
rect 50445 19125 50479 19159
rect 12633 18921 12667 18955
rect 22661 18921 22695 18955
rect 45569 18921 45603 18955
rect 46581 18921 46615 18955
rect 58081 18921 58115 18955
rect 10517 18853 10551 18887
rect 15853 18853 15887 18887
rect 25329 18853 25363 18887
rect 35725 18853 35759 18887
rect 36093 18853 36127 18887
rect 36369 18853 36403 18887
rect 36829 18853 36863 18887
rect 42717 18853 42751 18887
rect 18061 18785 18095 18819
rect 25973 18785 26007 18819
rect 28365 18785 28399 18819
rect 30297 18785 30331 18819
rect 37473 18785 37507 18819
rect 38669 18785 38703 18819
rect 41245 18785 41279 18819
rect 43361 18785 43395 18819
rect 1593 18717 1627 18751
rect 6285 18717 6319 18751
rect 9137 18717 9171 18751
rect 11437 18717 11471 18751
rect 14473 18717 14507 18751
rect 14740 18717 14774 18751
rect 16589 18717 16623 18751
rect 19441 18717 19475 18751
rect 21281 18717 21315 18751
rect 24593 18717 24627 18751
rect 24777 18717 24811 18751
rect 25789 18717 25823 18751
rect 26525 18717 26559 18751
rect 30564 18717 30598 18751
rect 32229 18717 32263 18751
rect 32413 18717 32447 18751
rect 33793 18717 33827 18751
rect 37197 18717 37231 18751
rect 38853 18717 38887 18751
rect 42902 18711 42936 18745
rect 45293 18717 45327 18751
rect 45385 18717 45419 18751
rect 46029 18717 46063 18751
rect 46305 18717 46339 18751
rect 46397 18717 46431 18751
rect 48329 18717 48363 18751
rect 48513 18717 48547 18751
rect 55505 18717 55539 18751
rect 55689 18717 55723 18751
rect 56977 18717 57011 18751
rect 57989 18717 58023 18751
rect 1869 18649 1903 18683
rect 2421 18649 2455 18683
rect 9404 18649 9438 18683
rect 19708 18649 19742 18683
rect 34069 18649 34103 18683
rect 42994 18649 43028 18683
rect 43085 18649 43119 18683
rect 43223 18649 43257 18683
rect 46213 18649 46247 18683
rect 47133 18649 47167 18683
rect 47501 18649 47535 18683
rect 57253 18649 57287 18683
rect 7481 18581 7515 18615
rect 20821 18581 20855 18615
rect 24685 18581 24719 18615
rect 25697 18581 25731 18615
rect 31677 18581 31711 18615
rect 32597 18581 32631 18615
rect 37289 18581 37323 18615
rect 39037 18581 39071 18615
rect 40601 18581 40635 18615
rect 40969 18581 41003 18615
rect 41061 18581 41095 18615
rect 48697 18581 48731 18615
rect 55873 18581 55907 18615
rect 7941 18377 7975 18411
rect 22017 18377 22051 18411
rect 30849 18377 30883 18411
rect 31309 18377 31343 18411
rect 42073 18377 42107 18411
rect 46397 18377 46431 18411
rect 54033 18377 54067 18411
rect 54953 18377 54987 18411
rect 57161 18377 57195 18411
rect 16313 18309 16347 18343
rect 22385 18309 22419 18343
rect 27804 18309 27838 18343
rect 41797 18309 41831 18343
rect 42993 18309 43027 18343
rect 46029 18309 46063 18343
rect 46121 18309 46155 18343
rect 54677 18309 54711 18343
rect 6561 18241 6595 18275
rect 6828 18241 6862 18275
rect 8585 18241 8619 18275
rect 11989 18241 12023 18275
rect 12817 18241 12851 18275
rect 16037 18241 16071 18275
rect 16129 18241 16163 18275
rect 17141 18241 17175 18275
rect 17408 18241 17442 18275
rect 19165 18241 19199 18275
rect 22477 18241 22511 18275
rect 23581 18241 23615 18275
rect 23673 18241 23707 18275
rect 24317 18241 24351 18275
rect 27537 18241 27571 18275
rect 29745 18241 29779 18275
rect 29837 18241 29871 18275
rect 30021 18241 30055 18275
rect 30113 18241 30147 18275
rect 31217 18241 31251 18275
rect 32137 18241 32171 18275
rect 34713 18241 34747 18275
rect 35449 18241 35483 18275
rect 38761 18241 38795 18275
rect 39037 18241 39071 18275
rect 41521 18241 41555 18275
rect 41705 18241 41739 18275
rect 41889 18241 41923 18275
rect 42625 18241 42659 18275
rect 42718 18241 42752 18275
rect 42901 18241 42935 18275
rect 43090 18241 43124 18275
rect 45845 18241 45879 18275
rect 46213 18241 46247 18275
rect 48780 18241 48814 18275
rect 54401 18241 54435 18275
rect 54585 18241 54619 18275
rect 54769 18241 54803 18275
rect 55781 18241 55815 18275
rect 56037 18241 56071 18275
rect 11897 18173 11931 18207
rect 22661 18173 22695 18207
rect 31493 18173 31527 18207
rect 35541 18173 35575 18207
rect 35725 18173 35759 18207
rect 48513 18173 48547 18207
rect 12357 18105 12391 18139
rect 18521 18105 18555 18139
rect 25513 18105 25547 18139
rect 33333 18105 33367 18139
rect 35081 18105 35115 18139
rect 43269 18105 43303 18139
rect 9781 18037 9815 18071
rect 14013 18037 14047 18071
rect 20361 18037 20395 18071
rect 23857 18037 23891 18071
rect 28917 18037 28951 18071
rect 29561 18037 29595 18071
rect 40141 18037 40175 18071
rect 49893 18037 49927 18071
rect 8033 17833 8067 17867
rect 11345 17833 11379 17867
rect 13369 17833 13403 17867
rect 15485 17833 15519 17867
rect 15669 17833 15703 17867
rect 17325 17833 17359 17867
rect 19441 17833 19475 17867
rect 24593 17833 24627 17867
rect 28641 17833 28675 17867
rect 32137 17833 32171 17867
rect 38761 17833 38795 17867
rect 48421 17833 48455 17867
rect 52837 17833 52871 17867
rect 58265 17833 58299 17867
rect 7573 17765 7607 17799
rect 13185 17765 13219 17799
rect 21281 17765 21315 17799
rect 30297 17765 30331 17799
rect 7297 17697 7331 17731
rect 8217 17697 8251 17731
rect 8493 17697 8527 17731
rect 9137 17697 9171 17731
rect 23213 17697 23247 17731
rect 25145 17697 25179 17731
rect 31677 17697 31711 17731
rect 32321 17697 32355 17731
rect 32413 17697 32447 17731
rect 33885 17697 33919 17731
rect 39313 17697 39347 17731
rect 55689 17697 55723 17731
rect 56885 17697 56919 17731
rect 1593 17629 1627 17663
rect 7205 17629 7239 17663
rect 8309 17629 8343 17663
rect 8401 17629 8435 17663
rect 9321 17629 9355 17663
rect 9505 17629 9539 17663
rect 10149 17629 10183 17663
rect 12909 17629 12943 17663
rect 14657 17629 14691 17663
rect 14841 17629 14875 17663
rect 16154 17629 16188 17663
rect 19441 17629 19475 17663
rect 19625 17629 19659 17663
rect 20085 17629 20119 17663
rect 23397 17629 23431 17663
rect 24961 17629 24995 17663
rect 26157 17629 26191 17663
rect 26424 17629 26458 17663
rect 28089 17629 28123 17663
rect 28365 17629 28399 17663
rect 28462 17629 28496 17663
rect 30573 17629 30607 17663
rect 31401 17629 31435 17663
rect 32506 17629 32540 17663
rect 32597 17629 32631 17663
rect 34897 17629 34931 17663
rect 35081 17629 35115 17663
rect 35265 17629 35299 17663
rect 40325 17629 40359 17663
rect 40592 17629 40626 17663
rect 47869 17629 47903 17663
rect 48237 17629 48271 17663
rect 50445 17629 50479 17663
rect 50721 17629 50755 17663
rect 50813 17629 50847 17663
rect 51457 17629 51491 17663
rect 55505 17629 55539 17663
rect 1869 17561 1903 17595
rect 9413 17561 9447 17595
rect 15301 17561 15335 17595
rect 28273 17561 28307 17595
rect 30849 17561 30883 17595
rect 33057 17561 33091 17595
rect 48053 17561 48087 17595
rect 48145 17561 48179 17595
rect 50629 17561 50663 17595
rect 51724 17561 51758 17595
rect 57130 17561 57164 17595
rect 9689 17493 9723 17527
rect 14749 17493 14783 17527
rect 15511 17493 15545 17527
rect 23581 17493 23615 17527
rect 25053 17493 25087 17527
rect 27537 17493 27571 17527
rect 30757 17493 30791 17527
rect 33333 17493 33367 17527
rect 33701 17493 33735 17527
rect 33793 17493 33827 17527
rect 39129 17493 39163 17527
rect 39221 17493 39255 17527
rect 41705 17493 41739 17527
rect 50997 17493 51031 17527
rect 13737 17289 13771 17323
rect 23213 17289 23247 17323
rect 26341 17289 26375 17323
rect 51733 17289 51767 17323
rect 56149 17289 56183 17323
rect 9873 17221 9907 17255
rect 25283 17221 25317 17255
rect 25421 17221 25455 17255
rect 27813 17221 27847 17255
rect 28917 17221 28951 17255
rect 38577 17221 38611 17255
rect 40969 17221 41003 17255
rect 41061 17221 41095 17255
rect 54953 17221 54987 17255
rect 55045 17221 55079 17255
rect 1593 17153 1627 17187
rect 2421 17153 2455 17187
rect 6745 17153 6779 17187
rect 8217 17153 8251 17187
rect 12541 17153 12575 17187
rect 15853 17153 15887 17187
rect 17049 17153 17083 17187
rect 17693 17153 17727 17187
rect 21097 17153 21131 17187
rect 22017 17153 22051 17187
rect 25145 17153 25179 17187
rect 26157 17153 26191 17187
rect 26295 17153 26329 17187
rect 26525 17153 26559 17187
rect 27261 17153 27295 17187
rect 27537 17153 27571 17187
rect 27721 17153 27755 17187
rect 27905 17153 27939 17187
rect 28549 17153 28583 17187
rect 28697 17153 28731 17187
rect 28825 17153 28859 17187
rect 29014 17153 29048 17187
rect 29745 17153 29779 17187
rect 30021 17153 30055 17187
rect 32781 17153 32815 17187
rect 33968 17153 34002 17187
rect 51365 17153 51399 17187
rect 51549 17153 51583 17187
rect 54128 17143 54162 17177
rect 54769 17153 54803 17187
rect 55137 17153 55171 17187
rect 55965 17153 55999 17187
rect 57069 17153 57103 17187
rect 1777 17085 1811 17119
rect 6837 17085 6871 17119
rect 7113 17085 7147 17119
rect 8493 17085 8527 17119
rect 16865 17085 16899 17119
rect 21189 17085 21223 17119
rect 21373 17085 21407 17119
rect 29837 17085 29871 17119
rect 30481 17085 30515 17119
rect 32321 17085 32355 17119
rect 32505 17085 32539 17119
rect 32597 17085 32631 17119
rect 32689 17085 32723 17119
rect 33701 17085 33735 17119
rect 38669 17085 38703 17119
rect 38853 17085 38887 17119
rect 41245 17085 41279 17119
rect 53941 17085 53975 17119
rect 55781 17085 55815 17119
rect 57345 17085 57379 17119
rect 16221 17017 16255 17051
rect 17233 17017 17267 17051
rect 20729 17017 20763 17051
rect 25973 17017 26007 17051
rect 28089 17017 28123 17051
rect 29193 17017 29227 17051
rect 55321 17017 55355 17051
rect 16313 16949 16347 16983
rect 18889 16949 18923 16983
rect 20361 16949 20395 16983
rect 24869 16949 24903 16983
rect 35081 16949 35115 16983
rect 38209 16949 38243 16983
rect 40601 16949 40635 16983
rect 54309 16949 54343 16983
rect 52377 16745 52411 16779
rect 13185 16677 13219 16711
rect 16129 16677 16163 16711
rect 22753 16677 22787 16711
rect 24593 16677 24627 16711
rect 11069 16609 11103 16643
rect 13461 16609 13495 16643
rect 13645 16609 13679 16643
rect 22293 16609 22327 16643
rect 23397 16609 23431 16643
rect 25697 16609 25731 16643
rect 27997 16609 28031 16643
rect 28181 16609 28215 16643
rect 28733 16609 28767 16643
rect 32505 16609 32539 16643
rect 32965 16609 32999 16643
rect 36737 16609 36771 16643
rect 37381 16609 37415 16643
rect 40509 16609 40543 16643
rect 41521 16609 41555 16643
rect 45201 16609 45235 16643
rect 53021 16609 53055 16643
rect 53573 16609 53607 16643
rect 1593 16541 1627 16575
rect 9137 16541 9171 16575
rect 9321 16541 9355 16575
rect 13369 16541 13403 16575
rect 13553 16541 13587 16575
rect 14749 16541 14783 16575
rect 16589 16541 16623 16575
rect 19993 16541 20027 16575
rect 22878 16541 22912 16575
rect 23305 16541 23339 16575
rect 23857 16541 23891 16575
rect 24777 16541 24811 16575
rect 25145 16541 25179 16575
rect 27905 16541 27939 16575
rect 28917 16541 28951 16575
rect 33232 16541 33266 16575
rect 37648 16541 37682 16575
rect 40693 16541 40727 16575
rect 40785 16541 40819 16575
rect 40969 16541 41003 16575
rect 41061 16541 41095 16575
rect 41705 16541 41739 16575
rect 41797 16541 41831 16575
rect 41981 16541 42015 16575
rect 42073 16541 42107 16575
rect 51365 16541 51399 16575
rect 51549 16541 51583 16575
rect 52193 16541 52227 16575
rect 52929 16541 52963 16575
rect 53113 16541 53147 16575
rect 53840 16541 53874 16575
rect 57989 16541 58023 16575
rect 1869 16473 1903 16507
rect 11336 16473 11370 16507
rect 15016 16473 15050 16507
rect 23003 16473 23037 16507
rect 25964 16473 25998 16507
rect 32137 16473 32171 16507
rect 32321 16473 32355 16507
rect 36553 16473 36587 16507
rect 45468 16473 45502 16507
rect 57069 16473 57103 16507
rect 9321 16405 9355 16439
rect 12449 16405 12483 16439
rect 17969 16405 18003 16439
rect 23949 16405 23983 16439
rect 24869 16405 24903 16439
rect 24961 16405 24995 16439
rect 27077 16405 27111 16439
rect 27537 16405 27571 16439
rect 29101 16405 29135 16439
rect 34345 16405 34379 16439
rect 36185 16405 36219 16439
rect 36645 16405 36679 16439
rect 38761 16405 38795 16439
rect 46581 16405 46615 16439
rect 51733 16405 51767 16439
rect 54953 16405 54987 16439
rect 57161 16405 57195 16439
rect 58081 16405 58115 16439
rect 15117 16201 15151 16235
rect 16221 16201 16255 16235
rect 19717 16201 19751 16235
rect 27261 16201 27295 16235
rect 40417 16201 40451 16235
rect 43177 16201 43211 16235
rect 45477 16201 45511 16235
rect 46397 16201 46431 16235
rect 46857 16201 46891 16235
rect 48145 16201 48179 16235
rect 54125 16201 54159 16235
rect 54769 16201 54803 16235
rect 17877 16133 17911 16167
rect 22262 16133 22296 16167
rect 27721 16133 27755 16167
rect 30481 16133 30515 16167
rect 37473 16133 37507 16167
rect 38485 16133 38519 16167
rect 39037 16133 39071 16167
rect 40141 16133 40175 16167
rect 42901 16133 42935 16167
rect 51264 16133 51298 16167
rect 53849 16133 53883 16167
rect 1593 16065 1627 16099
rect 10149 16065 10183 16099
rect 11897 16065 11931 16099
rect 13185 16065 13219 16099
rect 13452 16065 13486 16099
rect 15393 16065 15427 16099
rect 15485 16065 15519 16099
rect 16129 16065 16163 16099
rect 16313 16065 16347 16099
rect 17693 16065 17727 16099
rect 18521 16065 18555 16099
rect 21281 16065 21315 16099
rect 21465 16065 21499 16099
rect 23857 16065 23891 16099
rect 27629 16065 27663 16099
rect 28457 16065 28491 16099
rect 28724 16065 28758 16099
rect 30297 16065 30331 16099
rect 32413 16065 32447 16099
rect 32597 16065 32631 16099
rect 32689 16065 32723 16099
rect 32873 16065 32907 16099
rect 32965 16065 32999 16099
rect 37657 16065 37691 16099
rect 38669 16065 38703 16099
rect 39865 16065 39899 16099
rect 40049 16065 40083 16099
rect 40233 16065 40267 16099
rect 41521 16065 41555 16099
rect 41889 16065 41923 16099
rect 41981 16065 42015 16099
rect 42625 16065 42659 16099
rect 42809 16065 42843 16099
rect 42993 16065 43027 16099
rect 44189 16065 44223 16099
rect 46765 16065 46799 16099
rect 53573 16065 53607 16099
rect 53757 16065 53791 16099
rect 53941 16065 53975 16099
rect 54585 16065 54619 16099
rect 1777 15997 1811 16031
rect 2421 15997 2455 16031
rect 9965 15997 9999 16031
rect 11989 15997 12023 16031
rect 15301 15997 15335 16031
rect 15577 15997 15611 16031
rect 17969 15997 18003 16031
rect 22017 15997 22051 16031
rect 27905 15997 27939 16031
rect 30665 15997 30699 16031
rect 41613 15997 41647 16031
rect 46949 15997 46983 16031
rect 48237 15997 48271 16031
rect 48329 15997 48363 16031
rect 50997 15997 51031 16031
rect 17417 15929 17451 15963
rect 10333 15861 10367 15895
rect 12265 15861 12299 15895
rect 14565 15861 14599 15895
rect 21281 15861 21315 15895
rect 23397 15861 23431 15895
rect 25053 15861 25087 15895
rect 29837 15861 29871 15895
rect 37749 15861 37783 15895
rect 40969 15861 41003 15895
rect 47777 15861 47811 15895
rect 52377 15861 52411 15895
rect 13185 15657 13219 15691
rect 25145 15657 25179 15691
rect 29745 15657 29779 15691
rect 41705 15657 41739 15691
rect 51549 15657 51583 15691
rect 19441 15589 19475 15623
rect 19993 15589 20027 15623
rect 26249 15589 26283 15623
rect 13369 15521 13403 15555
rect 13461 15521 13495 15555
rect 13553 15521 13587 15555
rect 14289 15521 14323 15555
rect 15945 15521 15979 15555
rect 27353 15521 27387 15555
rect 30297 15521 30331 15555
rect 9873 15453 9907 15487
rect 13645 15453 13679 15487
rect 14565 15453 14599 15487
rect 16589 15453 16623 15487
rect 19625 15453 19659 15487
rect 19809 15453 19843 15487
rect 21097 15453 21131 15487
rect 23397 15453 23431 15487
rect 23857 15453 23891 15487
rect 24593 15453 24627 15487
rect 24869 15453 24903 15487
rect 24966 15453 25000 15487
rect 25697 15453 25731 15487
rect 26117 15453 26151 15487
rect 32137 15453 32171 15487
rect 32321 15453 32355 15487
rect 36369 15453 36403 15487
rect 36625 15453 36659 15487
rect 41061 15453 41095 15487
rect 41154 15453 41188 15487
rect 41337 15453 41371 15487
rect 41567 15453 41601 15487
rect 46857 15453 46891 15487
rect 50997 15453 51031 15487
rect 51181 15453 51215 15487
rect 51365 15453 51399 15487
rect 57897 15453 57931 15487
rect 24777 15385 24811 15419
rect 25881 15385 25915 15419
rect 25973 15385 26007 15419
rect 27620 15385 27654 15419
rect 30205 15385 30239 15419
rect 41429 15385 41463 15419
rect 51273 15385 51307 15419
rect 58173 15385 58207 15419
rect 11069 15317 11103 15351
rect 17969 15317 18003 15351
rect 19717 15317 19751 15351
rect 23949 15317 23983 15351
rect 28733 15317 28767 15351
rect 30113 15317 30147 15351
rect 37749 15317 37783 15351
rect 48145 15317 48179 15351
rect 13461 15113 13495 15147
rect 15761 15113 15795 15147
rect 20177 15113 20211 15147
rect 33885 15113 33919 15147
rect 38669 15113 38703 15147
rect 17132 15045 17166 15079
rect 28089 15045 28123 15079
rect 28181 15045 28215 15079
rect 1593 14977 1627 15011
rect 8861 14977 8895 15011
rect 12265 14977 12299 15011
rect 16037 14977 16071 15011
rect 16129 14977 16163 15011
rect 16221 14977 16255 15011
rect 16865 14977 16899 15011
rect 18981 14977 19015 15011
rect 22017 14977 22051 15011
rect 24777 14977 24811 15011
rect 25044 14977 25078 15011
rect 27905 14977 27939 15011
rect 28278 14977 28312 15011
rect 29193 14977 29227 15011
rect 29929 14977 29963 15011
rect 32597 14977 32631 15011
rect 34437 14977 34471 15011
rect 34704 14977 34738 15011
rect 38666 14977 38700 15011
rect 42901 14977 42935 15011
rect 1777 14909 1811 14943
rect 15945 14909 15979 14943
rect 23121 14909 23155 14943
rect 30205 14909 30239 14943
rect 32321 14909 32355 14943
rect 39129 14909 39163 14943
rect 43085 14909 43119 14943
rect 18245 14841 18279 14875
rect 28457 14841 28491 14875
rect 10057 14773 10091 14807
rect 26157 14773 26191 14807
rect 29285 14773 29319 14807
rect 35817 14773 35851 14807
rect 38485 14773 38519 14807
rect 39037 14773 39071 14807
rect 22845 14569 22879 14603
rect 27629 14569 27663 14603
rect 31125 14569 31159 14603
rect 31769 14569 31803 14603
rect 39405 14569 39439 14603
rect 41429 14569 41463 14603
rect 44557 14569 44591 14603
rect 48145 14569 48179 14603
rect 25053 14501 25087 14535
rect 2421 14433 2455 14467
rect 9321 14433 9355 14467
rect 9597 14433 9631 14467
rect 14289 14433 14323 14467
rect 25697 14433 25731 14467
rect 28825 14433 28859 14467
rect 32781 14433 32815 14467
rect 35541 14433 35575 14467
rect 37473 14433 37507 14467
rect 1593 14365 1627 14399
rect 11437 14365 11471 14399
rect 14565 14365 14599 14399
rect 16589 14365 16623 14399
rect 19717 14365 19751 14399
rect 21649 14365 21683 14399
rect 25513 14365 25547 14399
rect 26249 14365 26283 14399
rect 26525 14365 26559 14399
rect 26617 14365 26651 14399
rect 27261 14365 27295 14399
rect 27445 14365 27479 14399
rect 29009 14365 29043 14399
rect 29745 14365 29779 14399
rect 31769 14365 31803 14399
rect 31953 14365 31987 14399
rect 32689 14365 32723 14399
rect 32965 14365 32999 14399
rect 33149 14365 33183 14399
rect 33609 14365 33643 14399
rect 34253 14365 34287 14399
rect 37381 14365 37415 14399
rect 37565 14365 37599 14399
rect 38025 14365 38059 14399
rect 40049 14365 40083 14399
rect 42993 14365 43027 14399
rect 43269 14365 43303 14399
rect 46765 14365 46799 14399
rect 57989 14365 58023 14399
rect 1869 14297 1903 14331
rect 10977 14297 11011 14331
rect 19984 14297 20018 14331
rect 25421 14297 25455 14331
rect 26433 14297 26467 14331
rect 29193 14297 29227 14331
rect 29990 14297 30024 14331
rect 35357 14297 35391 14331
rect 38270 14297 38304 14331
rect 40294 14297 40328 14331
rect 47032 14297 47066 14331
rect 12633 14229 12667 14263
rect 15669 14229 15703 14263
rect 17785 14229 17819 14263
rect 21097 14229 21131 14263
rect 26801 14229 26835 14263
rect 34897 14229 34931 14263
rect 35265 14229 35299 14263
rect 58081 14229 58115 14263
rect 10057 14025 10091 14059
rect 13093 14025 13127 14059
rect 18245 14025 18279 14059
rect 24225 14025 24259 14059
rect 25145 14025 25179 14059
rect 27445 14025 27479 14059
rect 29285 14025 29319 14059
rect 32413 14025 32447 14059
rect 37933 14025 37967 14059
rect 38117 14025 38151 14059
rect 39129 14025 39163 14059
rect 17132 13957 17166 13991
rect 41797 13957 41831 13991
rect 1593 13889 1627 13923
rect 8861 13889 8895 13923
rect 11713 13889 11747 13923
rect 11980 13889 12014 13923
rect 13737 13889 13771 13923
rect 16865 13889 16899 13923
rect 19165 13889 19199 13923
rect 21465 13889 21499 13923
rect 21833 13889 21867 13923
rect 22100 13889 22134 13923
rect 23581 13889 23615 13923
rect 25320 13889 25354 13923
rect 25421 13889 25455 13923
rect 25605 13889 25639 13923
rect 25697 13889 25731 13923
rect 26157 13889 26191 13923
rect 27353 13889 27387 13923
rect 27537 13889 27571 13923
rect 29653 13889 29687 13923
rect 31125 13889 31159 13923
rect 31217 13889 31251 13923
rect 31493 13889 31527 13923
rect 31677 13889 31711 13923
rect 32597 13889 32631 13923
rect 32781 13889 32815 13923
rect 34897 13889 34931 13923
rect 38114 13889 38148 13923
rect 39037 13889 39071 13923
rect 39221 13889 39255 13923
rect 41521 13889 41555 13923
rect 41705 13889 41739 13923
rect 41889 13889 41923 13923
rect 43085 13889 43119 13923
rect 1777 13821 1811 13855
rect 15209 13821 15243 13855
rect 24317 13821 24351 13855
rect 24501 13821 24535 13855
rect 26433 13821 26467 13855
rect 29745 13821 29779 13855
rect 29837 13821 29871 13855
rect 34989 13821 35023 13855
rect 35173 13821 35207 13855
rect 38577 13821 38611 13855
rect 43361 13821 43395 13855
rect 44741 13821 44775 13855
rect 23213 13753 23247 13787
rect 23857 13753 23891 13787
rect 30573 13753 30607 13787
rect 38485 13753 38519 13787
rect 34529 13685 34563 13719
rect 42073 13685 42107 13719
rect 19533 13481 19567 13515
rect 22201 13481 22235 13515
rect 27353 13481 27387 13515
rect 28273 13481 28307 13515
rect 43637 13481 43671 13515
rect 42809 13413 42843 13447
rect 9321 13345 9355 13379
rect 9597 13345 9631 13379
rect 14289 13345 14323 13379
rect 18153 13345 18187 13379
rect 19993 13345 20027 13379
rect 25053 13345 25087 13379
rect 58173 13345 58207 13379
rect 1593 13277 1627 13311
rect 11437 13277 11471 13311
rect 14565 13277 14599 13311
rect 16589 13277 16623 13311
rect 21005 13277 21039 13311
rect 23857 13277 23891 13311
rect 24041 13277 24075 13311
rect 24777 13277 24811 13311
rect 24869 13277 24903 13311
rect 25145 13277 25179 13311
rect 28273 13277 28307 13311
rect 28457 13277 28491 13311
rect 31861 13277 31895 13311
rect 32229 13277 32263 13311
rect 36277 13277 36311 13311
rect 36461 13277 36495 13311
rect 38117 13277 38151 13311
rect 38669 13277 38703 13311
rect 42257 13277 42291 13311
rect 42625 13277 42659 13311
rect 43269 13277 43303 13311
rect 43453 13277 43487 13311
rect 56977 13277 57011 13311
rect 57897 13277 57931 13311
rect 1869 13209 1903 13243
rect 10977 13209 11011 13243
rect 20085 13209 20119 13243
rect 23949 13209 23983 13243
rect 24593 13209 24627 13243
rect 26065 13209 26099 13243
rect 32045 13209 32079 13243
rect 32137 13209 32171 13243
rect 37197 13209 37231 13243
rect 42441 13209 42475 13243
rect 42533 13209 42567 13243
rect 57253 13209 57287 13243
rect 12633 13141 12667 13175
rect 15669 13141 15703 13175
rect 19993 13141 20027 13175
rect 32413 13141 32447 13175
rect 36645 13141 36679 13175
rect 37289 13141 37323 13175
rect 38209 13141 38243 13175
rect 9965 12937 9999 12971
rect 11161 12937 11195 12971
rect 13553 12937 13587 12971
rect 15393 12937 15427 12971
rect 17233 12937 17267 12971
rect 43177 12937 43211 12971
rect 11897 12869 11931 12903
rect 12173 12869 12207 12903
rect 12265 12869 12299 12903
rect 16865 12869 16899 12903
rect 28641 12869 28675 12903
rect 30297 12869 30331 12903
rect 36001 12869 36035 12903
rect 36093 12869 36127 12903
rect 9597 12801 9631 12835
rect 12081 12801 12115 12835
rect 12633 12801 12667 12835
rect 14013 12801 14047 12835
rect 17049 12801 17083 12835
rect 17325 12801 17359 12835
rect 17785 12801 17819 12835
rect 21005 12801 21039 12835
rect 22017 12801 22051 12835
rect 24777 12801 24811 12835
rect 25044 12801 25078 12835
rect 27353 12801 27387 12835
rect 27445 12801 27479 12835
rect 30941 12801 30975 12835
rect 31125 12801 31159 12835
rect 31217 12801 31251 12835
rect 32689 12801 32723 12835
rect 32965 12801 32999 12835
rect 33885 12801 33919 12835
rect 34152 12801 34186 12835
rect 35817 12801 35851 12835
rect 36185 12801 36219 12835
rect 41797 12801 41831 12835
rect 42993 12801 43027 12835
rect 9505 12733 9539 12767
rect 10701 12733 10735 12767
rect 13093 12733 13127 12767
rect 20821 12733 20855 12767
rect 21189 12733 21223 12767
rect 28089 12733 28123 12767
rect 32781 12733 32815 12767
rect 33425 12733 33459 12767
rect 42809 12733 42843 12767
rect 10977 12665 11011 12699
rect 13461 12665 13495 12699
rect 36369 12665 36403 12699
rect 41981 12665 42015 12699
rect 18981 12597 19015 12631
rect 23213 12597 23247 12631
rect 26157 12597 26191 12631
rect 27353 12597 27387 12631
rect 27721 12597 27755 12631
rect 30941 12597 30975 12631
rect 35265 12597 35299 12631
rect 2237 12393 2271 12427
rect 10885 12393 10919 12427
rect 11713 12393 11747 12427
rect 15209 12393 15243 12427
rect 17141 12393 17175 12427
rect 19809 12393 19843 12427
rect 25421 12393 25455 12427
rect 32413 12393 32447 12427
rect 32873 12393 32907 12427
rect 13737 12325 13771 12359
rect 21281 12325 21315 12359
rect 11897 12257 11931 12291
rect 11989 12257 12023 12291
rect 13461 12257 13495 12291
rect 14565 12257 14599 12291
rect 14933 12257 14967 12291
rect 22753 12257 22787 12291
rect 23673 12257 23707 12291
rect 24961 12257 24995 12291
rect 26065 12257 26099 12291
rect 27077 12257 27111 12291
rect 32505 12257 32539 12291
rect 36645 12257 36679 12291
rect 41889 12257 41923 12291
rect 2145 12189 2179 12223
rect 2605 12189 2639 12223
rect 10517 12189 10551 12223
rect 12081 12189 12115 12223
rect 12173 12189 12207 12223
rect 13369 12189 13403 12223
rect 15945 12189 15979 12223
rect 18705 12189 18739 12223
rect 18889 12189 18923 12223
rect 19441 12189 19475 12223
rect 19625 12189 19659 12223
rect 20085 12189 20119 12223
rect 23397 12189 23431 12223
rect 24593 12189 24627 12223
rect 24777 12189 24811 12223
rect 25881 12189 25915 12223
rect 30113 12189 30147 12223
rect 30389 12189 30423 12223
rect 31033 12189 31067 12223
rect 31309 12189 31343 12223
rect 31769 12189 31803 12223
rect 31953 12189 31987 12223
rect 32689 12189 32723 12223
rect 35357 12189 35391 12223
rect 35633 12189 35667 12223
rect 35725 12189 35759 12223
rect 36369 12189 36403 12223
rect 40049 12189 40083 12223
rect 40142 12189 40176 12223
rect 40555 12189 40589 12223
rect 41797 12189 41831 12223
rect 42165 12189 42199 12223
rect 42349 12189 42383 12223
rect 57897 12189 57931 12223
rect 10701 12121 10735 12155
rect 15025 12121 15059 12155
rect 27322 12121 27356 12155
rect 30297 12121 30331 12155
rect 31861 12121 31895 12155
rect 32413 12121 32447 12155
rect 35541 12121 35575 12155
rect 38025 12121 38059 12155
rect 40325 12121 40359 12155
rect 40417 12121 40451 12155
rect 41153 12121 41187 12155
rect 58173 12121 58207 12155
rect 14841 12053 14875 12087
rect 18797 12053 18831 12087
rect 23029 12053 23063 12087
rect 23489 12053 23523 12087
rect 25789 12053 25823 12087
rect 28457 12053 28491 12087
rect 29929 12053 29963 12087
rect 30849 12053 30883 12087
rect 31217 12053 31251 12087
rect 35909 12053 35943 12087
rect 40693 12053 40727 12087
rect 10609 11849 10643 11883
rect 14565 11849 14599 11883
rect 15025 11849 15059 11883
rect 19007 11849 19041 11883
rect 19993 11849 20027 11883
rect 20361 11849 20395 11883
rect 20453 11849 20487 11883
rect 22385 11849 22419 11883
rect 26617 11849 26651 11883
rect 1869 11781 1903 11815
rect 13185 11781 13219 11815
rect 13401 11781 13435 11815
rect 17132 11781 17166 11815
rect 18797 11781 18831 11815
rect 40509 11781 40543 11815
rect 1593 11713 1627 11747
rect 10517 11713 10551 11747
rect 10701 11713 10735 11747
rect 11897 11713 11931 11747
rect 11989 11713 12023 11747
rect 14197 11713 14231 11747
rect 15209 11713 15243 11747
rect 15384 11713 15418 11747
rect 16037 11713 16071 11747
rect 16221 11713 16255 11747
rect 16865 11713 16899 11747
rect 22201 11713 22235 11747
rect 23857 11713 23891 11747
rect 25053 11713 25087 11747
rect 25237 11713 25271 11747
rect 26249 11713 26283 11747
rect 26433 11713 26467 11747
rect 27537 11713 27571 11747
rect 30481 11713 30515 11747
rect 30573 11713 30607 11747
rect 31125 11713 31159 11747
rect 31309 11713 31343 11747
rect 32965 11713 32999 11747
rect 33241 11713 33275 11747
rect 34713 11713 34747 11747
rect 34980 11713 35014 11747
rect 38761 11713 38795 11747
rect 43269 11713 43303 11747
rect 43361 11713 43395 11747
rect 43637 11713 43671 11747
rect 45477 11713 45511 11747
rect 45744 11713 45778 11747
rect 57161 11713 57195 11747
rect 11713 11645 11747 11679
rect 12081 11645 12115 11679
rect 12173 11645 12207 11679
rect 14289 11645 14323 11679
rect 15301 11645 15335 11679
rect 15486 11645 15520 11679
rect 20637 11645 20671 11679
rect 22017 11645 22051 11679
rect 25421 11645 25455 11679
rect 25605 11645 25639 11679
rect 27997 11645 28031 11679
rect 33425 11645 33459 11679
rect 43729 11645 43763 11679
rect 16129 11577 16163 11611
rect 18245 11577 18279 11611
rect 33057 11577 33091 11611
rect 13369 11509 13403 11543
rect 13553 11509 13587 11543
rect 18981 11509 19015 11543
rect 19165 11509 19199 11543
rect 23949 11509 23983 11543
rect 31125 11509 31159 11543
rect 36093 11509 36127 11543
rect 42717 11509 42751 11543
rect 46857 11509 46891 11543
rect 57253 11509 57287 11543
rect 15209 11305 15243 11339
rect 18061 11305 18095 11339
rect 21005 11305 21039 11339
rect 24041 11305 24075 11339
rect 28273 11305 28307 11339
rect 35357 11305 35391 11339
rect 46121 11305 46155 11339
rect 23121 11237 23155 11271
rect 31401 11237 31435 11271
rect 43085 11237 43119 11271
rect 56149 11237 56183 11271
rect 58265 11237 58299 11271
rect 1777 11169 1811 11203
rect 10977 11169 11011 11203
rect 11161 11169 11195 11203
rect 11253 11169 11287 11203
rect 11345 11169 11379 11203
rect 13185 11169 13219 11203
rect 14841 11169 14875 11203
rect 17877 11169 17911 11203
rect 30757 11169 30791 11203
rect 35817 11169 35851 11203
rect 36001 11169 36035 11203
rect 46673 11169 46707 11203
rect 1593 11101 1627 11135
rect 11437 11101 11471 11135
rect 13001 11101 13035 11135
rect 15025 11101 15059 11135
rect 15945 11101 15979 11135
rect 16405 11101 16439 11135
rect 16589 11101 16623 11135
rect 16865 11101 16899 11135
rect 17785 11101 17819 11135
rect 19625 11101 19659 11135
rect 19881 11101 19915 11135
rect 23029 11101 23063 11135
rect 23213 11101 23247 11135
rect 23765 11101 23799 11135
rect 23857 11101 23891 11135
rect 24593 11101 24627 11135
rect 26065 11101 26099 11135
rect 29929 11101 29963 11135
rect 31401 11101 31435 11135
rect 31585 11101 31619 11135
rect 31677 11101 31711 11135
rect 32137 11101 32171 11135
rect 32229 11101 32263 11135
rect 33793 11101 33827 11135
rect 34069 11101 34103 11135
rect 34161 11101 34195 11135
rect 35725 11101 35759 11135
rect 38485 11101 38519 11135
rect 40601 11101 40635 11135
rect 42441 11101 42475 11135
rect 42589 11101 42623 11135
rect 42717 11101 42751 11135
rect 42809 11101 42843 11135
rect 42906 11101 42940 11135
rect 44189 11101 44223 11135
rect 44465 11101 44499 11135
rect 46489 11101 46523 11135
rect 56425 11101 56459 11135
rect 56885 11101 56919 11135
rect 57141 11101 57175 11135
rect 25421 11033 25455 11067
rect 33977 11033 34011 11067
rect 38301 11033 38335 11067
rect 38853 11033 38887 11067
rect 40868 11033 40902 11067
rect 46581 11033 46615 11067
rect 56149 11033 56183 11067
rect 56333 11033 56367 11067
rect 15761 10965 15795 10999
rect 34345 10965 34379 10999
rect 41981 10965 42015 10999
rect 9229 10761 9263 10795
rect 12173 10761 12207 10795
rect 13369 10761 13403 10795
rect 27169 10761 27203 10795
rect 31309 10761 31343 10795
rect 41153 10761 41187 10795
rect 57253 10761 57287 10795
rect 1869 10693 1903 10727
rect 17049 10693 17083 10727
rect 17509 10693 17543 10727
rect 19962 10693 19996 10727
rect 23857 10693 23891 10727
rect 34805 10693 34839 10727
rect 53389 10693 53423 10727
rect 1593 10625 1627 10659
rect 9413 10625 9447 10659
rect 12909 10625 12943 10659
rect 13185 10625 13219 10659
rect 15761 10625 15795 10659
rect 16129 10625 16163 10659
rect 17417 10625 17451 10659
rect 18889 10625 18923 10659
rect 24196 10625 24230 10659
rect 25513 10625 25547 10659
rect 25881 10625 25915 10659
rect 27537 10625 27571 10659
rect 28733 10625 28767 10659
rect 31250 10625 31284 10659
rect 33333 10625 33367 10659
rect 35121 10625 35155 10659
rect 37473 10625 37507 10659
rect 41521 10625 41555 10659
rect 44189 10625 44223 10659
rect 53113 10625 53147 10659
rect 53297 10625 53331 10659
rect 53481 10625 53515 10659
rect 57161 10625 57195 10659
rect 57345 10625 57379 10659
rect 8953 10557 8987 10591
rect 9505 10557 9539 10591
rect 9597 10557 9631 10591
rect 9689 10557 9723 10591
rect 11713 10557 11747 10591
rect 15853 10557 15887 10591
rect 16221 10557 16255 10591
rect 16957 10557 16991 10591
rect 17969 10557 18003 10591
rect 18981 10557 19015 10591
rect 19165 10557 19199 10591
rect 19717 10557 19751 10591
rect 25973 10557 26007 10591
rect 27629 10557 27663 10591
rect 27813 10557 27847 10591
rect 29009 10557 29043 10591
rect 31677 10557 31711 10591
rect 31769 10557 31803 10591
rect 33701 10557 33735 10591
rect 34897 10557 34931 10591
rect 37749 10557 37783 10591
rect 41613 10557 41647 10591
rect 41797 10557 41831 10591
rect 11989 10489 12023 10523
rect 13001 10489 13035 10523
rect 15209 10489 15243 10523
rect 18521 10489 18555 10523
rect 24133 10489 24167 10523
rect 25329 10489 25363 10523
rect 31125 10489 31159 10523
rect 53665 10489 53699 10523
rect 21097 10421 21131 10455
rect 24022 10421 24056 10455
rect 24501 10421 24535 10455
rect 30297 10421 30331 10455
rect 35081 10421 35115 10455
rect 35265 10421 35299 10455
rect 45477 10421 45511 10455
rect 11529 10217 11563 10251
rect 28181 10217 28215 10251
rect 31953 10217 31987 10251
rect 48145 10217 48179 10251
rect 11345 10149 11379 10183
rect 12909 10149 12943 10183
rect 18153 10149 18187 10183
rect 21649 10149 21683 10183
rect 23489 10149 23523 10183
rect 1777 10081 1811 10115
rect 14933 10081 14967 10115
rect 18613 10081 18647 10115
rect 18797 10081 18831 10115
rect 22201 10081 22235 10115
rect 27813 10081 27847 10115
rect 58173 10081 58207 10115
rect 1593 10013 1627 10047
rect 12817 10013 12851 10047
rect 13093 10013 13127 10047
rect 14381 10013 14415 10047
rect 15945 10013 15979 10047
rect 16313 10013 16347 10047
rect 16681 10013 16715 10047
rect 17325 10013 17359 10047
rect 18521 10013 18555 10047
rect 19809 10013 19843 10047
rect 22017 10013 22051 10047
rect 24041 10013 24075 10047
rect 24593 10013 24627 10047
rect 24780 10013 24814 10047
rect 25145 10013 25179 10047
rect 27261 10013 27295 10047
rect 27997 10013 28031 10047
rect 28825 10013 28859 10047
rect 29193 10013 29227 10047
rect 29929 10013 29963 10047
rect 30021 10013 30055 10047
rect 30205 10013 30239 10047
rect 30297 10013 30331 10047
rect 30757 10013 30791 10047
rect 32137 10013 32171 10047
rect 32413 10013 32447 10047
rect 33333 10013 33367 10047
rect 33426 10013 33460 10047
rect 33609 10013 33643 10047
rect 33839 10013 33873 10047
rect 34989 10013 35023 10047
rect 37105 10013 37139 10047
rect 37381 10013 37415 10047
rect 37473 10013 37507 10047
rect 38117 10013 38151 10047
rect 38393 10013 38427 10047
rect 38531 10013 38565 10047
rect 44097 10013 44131 10047
rect 44189 10013 44223 10047
rect 44281 10013 44315 10047
rect 44459 10013 44493 10047
rect 45937 10013 45971 10047
rect 46213 10013 46247 10047
rect 46857 10013 46891 10047
rect 57897 10013 57931 10047
rect 11069 9945 11103 9979
rect 16865 9945 16899 9979
rect 20076 9945 20110 9979
rect 23673 9945 23707 9979
rect 24979 9945 25013 9979
rect 25605 9945 25639 9979
rect 28641 9945 28675 9979
rect 31033 9945 31067 9979
rect 32321 9945 32355 9979
rect 33701 9945 33735 9979
rect 35173 9945 35207 9979
rect 35357 9945 35391 9979
rect 37289 9945 37323 9979
rect 38301 9945 38335 9979
rect 57069 9945 57103 9979
rect 13277 9877 13311 9911
rect 21189 9877 21223 9911
rect 22109 9877 22143 9911
rect 23765 9877 23799 9911
rect 23857 9877 23891 9911
rect 24869 9877 24903 9911
rect 28917 9877 28951 9911
rect 29009 9877 29043 9911
rect 29745 9877 29779 9911
rect 33977 9877 34011 9911
rect 37657 9877 37691 9911
rect 38669 9877 38703 9911
rect 43821 9877 43855 9911
rect 45753 9877 45787 9911
rect 46121 9877 46155 9911
rect 57161 9877 57195 9911
rect 22017 9673 22051 9707
rect 22385 9673 22419 9707
rect 27537 9673 27571 9707
rect 29285 9673 29319 9707
rect 29469 9673 29503 9707
rect 29561 9673 29595 9707
rect 32505 9673 32539 9707
rect 33339 9673 33373 9707
rect 46581 9673 46615 9707
rect 20076 9605 20110 9639
rect 23673 9605 23707 9639
rect 27353 9605 27387 9639
rect 28365 9605 28399 9639
rect 29745 9605 29779 9639
rect 37749 9605 37783 9639
rect 38945 9605 38979 9639
rect 44005 9605 44039 9639
rect 45468 9605 45502 9639
rect 1593 9537 1627 9571
rect 13369 9537 13403 9571
rect 13461 9537 13495 9571
rect 13645 9537 13679 9571
rect 13737 9537 13771 9571
rect 14197 9537 14231 9571
rect 15301 9537 15335 9571
rect 15577 9537 15611 9571
rect 15669 9537 15703 9571
rect 15945 9537 15979 9571
rect 16221 9537 16255 9571
rect 17049 9537 17083 9571
rect 18889 9537 18923 9571
rect 24041 9537 24075 9571
rect 24133 9537 24167 9571
rect 24225 9537 24259 9571
rect 25237 9537 25271 9571
rect 25421 9537 25455 9571
rect 25605 9537 25639 9571
rect 25881 9537 25915 9571
rect 26157 9537 26191 9571
rect 27491 9537 27525 9571
rect 27721 9537 27755 9571
rect 28181 9537 28215 9571
rect 28457 9537 28491 9571
rect 28595 9537 28629 9571
rect 29377 9537 29411 9571
rect 30205 9537 30239 9571
rect 31033 9537 31067 9571
rect 32597 9537 32631 9571
rect 32781 9537 32815 9571
rect 33241 9537 33275 9571
rect 33425 9537 33459 9571
rect 33517 9537 33551 9571
rect 36001 9537 36035 9571
rect 36185 9537 36219 9571
rect 37473 9537 37507 9571
rect 37621 9537 37655 9571
rect 37841 9537 37875 9571
rect 37979 9537 38013 9571
rect 38577 9537 38611 9571
rect 38670 9537 38704 9571
rect 38853 9537 38887 9571
rect 39083 9537 39117 9571
rect 44097 9537 44131 9571
rect 44189 9537 44223 9571
rect 45201 9537 45235 9571
rect 56977 9537 57011 9571
rect 57161 9537 57195 9571
rect 1777 9469 1811 9503
rect 8769 9469 8803 9503
rect 9229 9469 9263 9503
rect 14289 9469 14323 9503
rect 18061 9469 18095 9503
rect 19165 9469 19199 9503
rect 19809 9469 19843 9503
rect 22477 9469 22511 9503
rect 22569 9469 22603 9503
rect 23489 9469 23523 9503
rect 24777 9469 24811 9503
rect 9045 9401 9079 9435
rect 14933 9401 14967 9435
rect 27169 9401 27203 9435
rect 28733 9401 28767 9435
rect 39221 9401 39255 9435
rect 43821 9401 43855 9435
rect 13185 9333 13219 9367
rect 21189 9333 21223 9367
rect 30389 9333 30423 9367
rect 31309 9333 31343 9367
rect 32321 9333 32355 9367
rect 36001 9333 36035 9367
rect 38117 9333 38151 9367
rect 44373 9333 44407 9367
rect 57069 9333 57103 9367
rect 13369 9129 13403 9163
rect 21281 9129 21315 9163
rect 28457 9129 28491 9163
rect 39037 9129 39071 9163
rect 46213 9129 46247 9163
rect 13277 9061 13311 9095
rect 14749 9061 14783 9095
rect 31401 9061 31435 9095
rect 32873 9061 32907 9095
rect 40049 9061 40083 9095
rect 56149 9061 56183 9095
rect 18337 8993 18371 9027
rect 24685 8993 24719 9027
rect 27905 8993 27939 9027
rect 29101 8993 29135 9027
rect 30757 8993 30791 9027
rect 36277 8993 36311 9027
rect 44465 8993 44499 9027
rect 56885 8993 56919 9027
rect 1593 8925 1627 8959
rect 15301 8925 15335 8959
rect 18061 8925 18095 8959
rect 19901 8925 19935 8959
rect 23489 8925 23523 8959
rect 23673 8925 23707 8959
rect 24777 8925 24811 8959
rect 25237 8925 25271 8959
rect 25697 8925 25731 8959
rect 25881 8925 25915 8959
rect 26249 8925 26283 8959
rect 26433 8925 26467 8959
rect 26617 8925 26651 8959
rect 27629 8925 27663 8959
rect 27813 8925 27847 8959
rect 30021 8925 30055 8959
rect 31585 8925 31619 8959
rect 33149 8925 33183 8959
rect 33333 8925 33367 8959
rect 33793 8925 33827 8959
rect 35817 8925 35851 8959
rect 36369 8925 36403 8959
rect 37749 8925 37783 8959
rect 37842 8925 37876 8959
rect 38117 8925 38151 8959
rect 38233 8925 38267 8959
rect 39037 8925 39071 8959
rect 40049 8925 40083 8959
rect 40325 8925 40359 8959
rect 40785 8925 40819 8959
rect 45201 8925 45235 8959
rect 46121 8925 46155 8959
rect 46305 8925 46339 8959
rect 56149 8925 56183 8959
rect 56333 8925 56367 8959
rect 56425 8925 56459 8959
rect 57141 8925 57175 8959
rect 1869 8857 1903 8891
rect 12909 8857 12943 8891
rect 14933 8857 14967 8891
rect 15761 8857 15795 8891
rect 17509 8857 17543 8891
rect 24041 8857 24075 8891
rect 28917 8857 28951 8891
rect 31953 8857 31987 8891
rect 34069 8857 34103 8891
rect 38025 8857 38059 8891
rect 43729 8857 43763 8891
rect 45477 8857 45511 8891
rect 15025 8789 15059 8823
rect 15117 8789 15151 8823
rect 23765 8789 23799 8823
rect 23857 8789 23891 8823
rect 27077 8789 27111 8823
rect 28825 8789 28859 8823
rect 31677 8789 31711 8823
rect 31769 8789 31803 8823
rect 33057 8789 33091 8823
rect 36001 8789 36035 8823
rect 38393 8789 38427 8823
rect 40233 8789 40267 8823
rect 40877 8789 40911 8823
rect 58265 8789 58299 8823
rect 14105 8585 14139 8619
rect 16221 8585 16255 8619
rect 19441 8585 19475 8619
rect 23397 8585 23431 8619
rect 23489 8585 23523 8619
rect 25329 8585 25363 8619
rect 33425 8585 33459 8619
rect 44281 8585 44315 8619
rect 56333 8585 56367 8619
rect 17049 8517 17083 8551
rect 23673 8517 23707 8551
rect 30941 8517 30975 8551
rect 33057 8517 33091 8551
rect 34161 8517 34195 8551
rect 57345 8517 57379 8551
rect 1593 8449 1627 8483
rect 14013 8449 14047 8483
rect 15209 8449 15243 8483
rect 15393 8449 15427 8483
rect 16129 8449 16163 8483
rect 16957 8449 16991 8483
rect 17417 8449 17451 8483
rect 17509 8449 17543 8483
rect 17601 8449 17635 8483
rect 18337 8449 18371 8483
rect 18705 8449 18739 8483
rect 19073 8449 19107 8483
rect 19901 8449 19935 8483
rect 22385 8449 22419 8483
rect 23305 8449 23339 8483
rect 24133 8449 24167 8483
rect 27169 8449 27203 8483
rect 29469 8449 29503 8483
rect 31677 8449 31711 8483
rect 32781 8449 32815 8483
rect 32874 8449 32908 8483
rect 33149 8449 33183 8483
rect 33287 8449 33321 8483
rect 33885 8449 33919 8483
rect 33978 8449 34012 8483
rect 34261 8449 34295 8483
rect 34391 8449 34425 8483
rect 35909 8449 35943 8483
rect 36737 8449 36771 8483
rect 37473 8449 37507 8483
rect 37565 8449 37599 8483
rect 37749 8449 37783 8483
rect 39385 8449 39419 8483
rect 42901 8449 42935 8483
rect 44465 8449 44499 8483
rect 44557 8449 44591 8483
rect 44741 8449 44775 8483
rect 44833 8449 44867 8483
rect 45293 8449 45327 8483
rect 46397 8449 46431 8483
rect 56241 8449 56275 8483
rect 57069 8449 57103 8483
rect 1777 8381 1811 8415
rect 27629 8381 27663 8415
rect 30113 8381 30147 8415
rect 31309 8381 31343 8415
rect 35357 8381 35391 8415
rect 35633 8381 35667 8415
rect 35817 8381 35851 8415
rect 36553 8381 36587 8415
rect 37933 8381 37967 8415
rect 39129 8381 39163 8415
rect 43177 8381 43211 8415
rect 45477 8381 45511 8415
rect 46581 8381 46615 8415
rect 15577 8313 15611 8347
rect 23121 8313 23155 8347
rect 31217 8313 31251 8347
rect 34529 8313 34563 8347
rect 40509 8313 40543 8347
rect 15393 8245 15427 8279
rect 22569 8245 22603 8279
rect 31106 8245 31140 8279
rect 36921 8245 36955 8279
rect 34161 8041 34195 8075
rect 38669 8041 38703 8075
rect 42901 8041 42935 8075
rect 45385 8041 45419 8075
rect 58265 8041 58299 8075
rect 12817 7973 12851 8007
rect 20821 7973 20855 8007
rect 26157 7973 26191 8007
rect 30941 7973 30975 8007
rect 31493 7973 31527 8007
rect 32597 7973 32631 8007
rect 35265 7973 35299 8007
rect 38945 7973 38979 8007
rect 56149 7973 56183 8007
rect 11161 7905 11195 7939
rect 19441 7905 19475 7939
rect 23305 7905 23339 7939
rect 28733 7905 28767 7939
rect 29837 7905 29871 7939
rect 39037 7905 39071 7939
rect 46673 7905 46707 7939
rect 56885 7905 56919 7939
rect 1593 7837 1627 7871
rect 7849 7837 7883 7871
rect 7941 7837 7975 7871
rect 8125 7837 8159 7871
rect 9965 7837 9999 7871
rect 10241 7837 10275 7871
rect 10885 7837 10919 7871
rect 15209 7837 15243 7871
rect 15485 7837 15519 7871
rect 16497 7837 16531 7871
rect 17049 7837 17083 7871
rect 17233 7837 17267 7871
rect 17969 7837 18003 7871
rect 24961 7837 24995 7871
rect 28365 7837 28399 7871
rect 30021 7837 30055 7871
rect 30113 7837 30147 7871
rect 31401 7837 31435 7871
rect 31677 7837 31711 7871
rect 32781 7837 32815 7871
rect 34161 7837 34195 7871
rect 34345 7837 34379 7871
rect 36277 7837 36311 7871
rect 36544 7837 36578 7871
rect 38862 7837 38896 7871
rect 39129 7837 39163 7871
rect 39313 7837 39347 7871
rect 42809 7837 42843 7871
rect 43729 7837 43763 7871
rect 44005 7837 44039 7871
rect 45293 7837 45327 7871
rect 45569 7837 45603 7871
rect 46305 7837 46339 7871
rect 55505 7837 55539 7871
rect 55689 7837 55723 7871
rect 56425 7837 56459 7871
rect 57141 7837 57175 7871
rect 1869 7769 1903 7803
rect 8585 7769 8619 7803
rect 9781 7769 9815 7803
rect 12541 7769 12575 7803
rect 15669 7769 15703 7803
rect 15945 7769 15979 7803
rect 19708 7769 19742 7803
rect 30481 7769 30515 7803
rect 33149 7769 33183 7803
rect 34989 7769 35023 7803
rect 43913 7769 43947 7803
rect 44465 7769 44499 7803
rect 45477 7769 45511 7803
rect 56149 7769 56183 7803
rect 10149 7701 10183 7735
rect 13001 7701 13035 7735
rect 15577 7701 15611 7735
rect 16497 7701 16531 7735
rect 22661 7701 22695 7735
rect 23029 7701 23063 7735
rect 23121 7701 23155 7735
rect 31861 7701 31895 7735
rect 32873 7701 32907 7735
rect 32965 7701 32999 7735
rect 37657 7701 37691 7735
rect 55689 7701 55723 7735
rect 56333 7701 56367 7735
rect 10609 7497 10643 7531
rect 19257 7497 19291 7531
rect 23489 7497 23523 7531
rect 27905 7497 27939 7531
rect 29929 7497 29963 7531
rect 35449 7497 35483 7531
rect 36185 7497 36219 7531
rect 11989 7429 12023 7463
rect 15301 7429 15335 7463
rect 15853 7429 15887 7463
rect 16957 7429 16991 7463
rect 17509 7429 17543 7463
rect 18521 7429 18555 7463
rect 19073 7429 19107 7463
rect 55873 7429 55907 7463
rect 58173 7429 58207 7463
rect 9505 7361 9539 7395
rect 10977 7361 11011 7395
rect 11805 7361 11839 7395
rect 15761 7361 15795 7395
rect 17371 7361 17405 7395
rect 18981 7361 19015 7395
rect 20085 7361 20119 7395
rect 20352 7361 20386 7395
rect 23305 7361 23339 7395
rect 23673 7361 23707 7395
rect 24317 7361 24351 7395
rect 27445 7361 27479 7395
rect 27537 7361 27571 7395
rect 27721 7361 27755 7395
rect 28641 7361 28675 7395
rect 30849 7361 30883 7395
rect 32597 7361 32631 7395
rect 32781 7361 32815 7395
rect 32873 7361 32907 7395
rect 34069 7361 34103 7395
rect 34336 7361 34370 7395
rect 36553 7361 36587 7395
rect 36645 7361 36679 7395
rect 44373 7361 44407 7395
rect 44465 7361 44499 7395
rect 45017 7361 45051 7395
rect 45284 7361 45318 7395
rect 55689 7361 55723 7395
rect 55965 7361 55999 7395
rect 56517 7361 56551 7395
rect 58081 7361 58115 7395
rect 58265 7361 58299 7395
rect 10793 7293 10827 7327
rect 10885 7293 10919 7327
rect 11069 7293 11103 7327
rect 12449 7293 12483 7327
rect 15393 7293 15427 7327
rect 16313 7293 16347 7327
rect 17049 7293 17083 7327
rect 17969 7293 18003 7327
rect 31033 7293 31067 7327
rect 36737 7293 36771 7327
rect 56793 7293 56827 7327
rect 12725 7225 12759 7259
rect 12909 7225 12943 7259
rect 18503 7225 18537 7259
rect 25513 7225 25547 7259
rect 9689 7157 9723 7191
rect 21465 7157 21499 7191
rect 23857 7157 23891 7191
rect 32413 7157 32447 7191
rect 35909 7157 35943 7191
rect 46397 7157 46431 7191
rect 55689 7157 55723 7191
rect 21189 6953 21223 6987
rect 34345 6953 34379 6987
rect 45201 6953 45235 6987
rect 45845 6953 45879 6987
rect 23857 6885 23891 6919
rect 30849 6885 30883 6919
rect 34897 6885 34931 6919
rect 10793 6817 10827 6851
rect 18705 6817 18739 6851
rect 19809 6817 19843 6851
rect 21741 6817 21775 6851
rect 26525 6817 26559 6851
rect 27261 6817 27295 6851
rect 28549 6817 28583 6851
rect 30205 6817 30239 6851
rect 31861 6817 31895 6851
rect 31953 6817 31987 6851
rect 32597 6817 32631 6851
rect 33977 6817 34011 6851
rect 35449 6817 35483 6851
rect 36553 6817 36587 6851
rect 46305 6817 46339 6851
rect 46489 6817 46523 6851
rect 1593 6749 1627 6783
rect 9597 6749 9631 6783
rect 10977 6749 11011 6783
rect 11069 6749 11103 6783
rect 11161 6749 11195 6783
rect 11253 6749 11287 6783
rect 16589 6749 16623 6783
rect 19533 6749 19567 6783
rect 22477 6749 22511 6783
rect 24685 6749 24719 6783
rect 27169 6749 27203 6783
rect 27503 6749 27537 6783
rect 27629 6749 27663 6783
rect 28181 6749 28215 6783
rect 30021 6749 30055 6783
rect 30113 6749 30147 6783
rect 31769 6749 31803 6783
rect 32781 6749 32815 6783
rect 32965 6749 32999 6783
rect 34161 6749 34195 6783
rect 36461 6749 36495 6783
rect 36645 6749 36679 6783
rect 45201 6749 45235 6783
rect 45385 6749 45419 6783
rect 56885 6749 56919 6783
rect 57141 6749 57175 6783
rect 1869 6681 1903 6715
rect 17325 6681 17359 6715
rect 17877 6681 17911 6715
rect 21557 6681 21591 6715
rect 22744 6681 22778 6715
rect 24952 6681 24986 6715
rect 30481 6681 30515 6715
rect 35357 6681 35391 6715
rect 46213 6681 46247 6715
rect 9781 6613 9815 6647
rect 18153 6613 18187 6647
rect 18521 6613 18555 6647
rect 18613 6613 18647 6647
rect 21649 6613 21683 6647
rect 26065 6613 26099 6647
rect 31401 6613 31435 6647
rect 35265 6613 35299 6647
rect 58265 6613 58299 6647
rect 9137 6409 9171 6443
rect 14381 6409 14415 6443
rect 24685 6409 24719 6443
rect 25605 6409 25639 6443
rect 30481 6409 30515 6443
rect 37657 6409 37691 6443
rect 46765 6409 46799 6443
rect 13553 6341 13587 6375
rect 15393 6341 15427 6375
rect 18245 6341 18279 6375
rect 23397 6341 23431 6375
rect 57161 6341 57195 6375
rect 1593 6273 1627 6307
rect 9321 6273 9355 6307
rect 9413 6273 9447 6307
rect 14289 6273 14323 6307
rect 15301 6273 15335 6307
rect 15761 6273 15795 6307
rect 15853 6273 15887 6307
rect 16313 6273 16347 6307
rect 17509 6273 17543 6307
rect 19697 6273 19731 6307
rect 22385 6273 22419 6307
rect 25973 6273 26007 6307
rect 27169 6273 27203 6307
rect 29101 6273 29135 6307
rect 33885 6273 33919 6307
rect 34529 6273 34563 6307
rect 35541 6273 35575 6307
rect 35909 6273 35943 6307
rect 36461 6273 36495 6307
rect 37565 6273 37599 6307
rect 46489 6273 46523 6307
rect 46581 6273 46615 6307
rect 1777 6205 1811 6239
rect 9505 6205 9539 6239
rect 9597 6205 9631 6239
rect 19441 6205 19475 6239
rect 26065 6205 26099 6239
rect 26157 6205 26191 6239
rect 27445 6205 27479 6239
rect 34713 6205 34747 6239
rect 13737 6137 13771 6171
rect 22569 6137 22603 6171
rect 27721 6137 27755 6171
rect 34069 6137 34103 6171
rect 20821 6069 20855 6103
rect 27537 6069 27571 6103
rect 36553 6069 36587 6103
rect 57253 6069 57287 6103
rect 9137 5865 9171 5899
rect 10885 5865 10919 5899
rect 13737 5865 13771 5899
rect 23029 5865 23063 5899
rect 26157 5865 26191 5899
rect 29910 5865 29944 5899
rect 30021 5865 30055 5899
rect 10701 5797 10735 5831
rect 13553 5797 13587 5831
rect 14565 5797 14599 5831
rect 36001 5797 36035 5831
rect 38393 5797 38427 5831
rect 40325 5797 40359 5831
rect 41613 5797 41647 5831
rect 9413 5729 9447 5763
rect 9505 5729 9539 5763
rect 15669 5729 15703 5763
rect 15761 5729 15795 5763
rect 21649 5729 21683 5763
rect 23581 5729 23615 5763
rect 30113 5729 30147 5763
rect 31217 5729 31251 5763
rect 36553 5729 36587 5763
rect 39313 5729 39347 5763
rect 58173 5729 58207 5763
rect 1593 5661 1627 5695
rect 9321 5661 9355 5695
rect 9597 5661 9631 5695
rect 16129 5661 16163 5695
rect 16217 5661 16251 5695
rect 16359 5661 16393 5695
rect 17049 5661 17083 5695
rect 17601 5661 17635 5695
rect 17877 5661 17911 5695
rect 18613 5661 18647 5695
rect 19625 5661 19659 5695
rect 19881 5661 19915 5695
rect 21465 5661 21499 5695
rect 22569 5661 22603 5695
rect 23489 5661 23523 5695
rect 24961 5661 24995 5695
rect 27905 5661 27939 5695
rect 28549 5661 28583 5695
rect 28917 5661 28951 5695
rect 30481 5661 30515 5695
rect 31484 5661 31518 5695
rect 33425 5661 33459 5695
rect 34161 5661 34195 5695
rect 34989 5661 35023 5695
rect 35725 5661 35759 5695
rect 36461 5661 36495 5695
rect 37473 5661 37507 5695
rect 37657 5661 37691 5695
rect 56977 5661 57011 5695
rect 57897 5661 57931 5695
rect 1869 5593 1903 5627
rect 10425 5593 10459 5627
rect 13277 5593 13311 5627
rect 14289 5593 14323 5627
rect 29745 5593 29779 5627
rect 33609 5593 33643 5627
rect 35173 5593 35207 5627
rect 39129 5593 39163 5627
rect 39221 5593 39255 5627
rect 40141 5593 40175 5627
rect 41429 5593 41463 5627
rect 57253 5593 57287 5627
rect 14749 5525 14783 5559
rect 18337 5525 18371 5559
rect 21005 5525 21039 5559
rect 23397 5525 23431 5559
rect 32597 5525 32631 5559
rect 34253 5525 34287 5559
rect 36369 5525 36403 5559
rect 37841 5525 37875 5559
rect 38761 5525 38795 5559
rect 9413 5321 9447 5355
rect 10149 5321 10183 5355
rect 14197 5321 14231 5355
rect 19257 5321 19291 5355
rect 19717 5321 19751 5355
rect 20637 5321 20671 5355
rect 25881 5321 25915 5355
rect 31125 5321 31159 5355
rect 31217 5321 31251 5355
rect 41981 5321 42015 5355
rect 42809 5321 42843 5355
rect 43545 5321 43579 5355
rect 58265 5321 58299 5355
rect 8953 5253 8987 5287
rect 12909 5253 12943 5287
rect 21097 5253 21131 5287
rect 28457 5253 28491 5287
rect 30849 5253 30883 5287
rect 32873 5253 32907 5287
rect 33609 5253 33643 5287
rect 34345 5253 34379 5287
rect 1593 5185 1627 5219
rect 8309 5185 8343 5219
rect 10333 5185 10367 5219
rect 10517 5185 10551 5219
rect 12173 5185 12207 5219
rect 14013 5185 14047 5219
rect 17049 5185 17083 5219
rect 17325 5185 17359 5219
rect 18061 5185 18095 5219
rect 19625 5185 19659 5219
rect 21005 5185 21039 5219
rect 22569 5185 22603 5219
rect 25145 5185 25179 5219
rect 26249 5185 26283 5219
rect 27169 5185 27203 5219
rect 27261 5185 27295 5219
rect 28549 5185 28583 5219
rect 29745 5185 29779 5219
rect 29929 5185 29963 5219
rect 30021 5185 30055 5219
rect 30165 5185 30199 5219
rect 31033 5185 31067 5219
rect 31401 5185 31435 5219
rect 34989 5185 35023 5219
rect 35909 5185 35943 5219
rect 37473 5185 37507 5219
rect 37657 5185 37691 5219
rect 38945 5185 38979 5219
rect 39681 5185 39715 5219
rect 40325 5185 40359 5219
rect 41153 5185 41187 5219
rect 41797 5185 41831 5219
rect 42717 5185 42751 5219
rect 43453 5185 43487 5219
rect 44189 5185 44223 5219
rect 44925 5185 44959 5219
rect 45845 5185 45879 5219
rect 48789 5185 48823 5219
rect 49045 5185 49079 5219
rect 58081 5185 58115 5219
rect 1777 5117 1811 5151
rect 10425 5117 10459 5151
rect 10609 5117 10643 5151
rect 13369 5117 13403 5151
rect 18337 5117 18371 5151
rect 19901 5117 19935 5151
rect 21281 5117 21315 5151
rect 22753 5117 22787 5151
rect 26341 5117 26375 5151
rect 26525 5117 26559 5151
rect 28733 5117 28767 5151
rect 35173 5117 35207 5151
rect 36093 5117 36127 5151
rect 38761 5117 38795 5151
rect 46029 5117 46063 5151
rect 8493 5049 8527 5083
rect 9229 5049 9263 5083
rect 12357 5049 12391 5083
rect 13185 5049 13219 5083
rect 24041 5049 24075 5083
rect 33057 5049 33091 5083
rect 33793 5049 33827 5083
rect 44373 5049 44407 5083
rect 16313 4981 16347 5015
rect 20269 4981 20303 5015
rect 24685 4981 24719 5015
rect 25329 4981 25363 5015
rect 27169 4981 27203 5015
rect 27537 4981 27571 5015
rect 28089 4981 28123 5015
rect 30297 4981 30331 5015
rect 34437 4981 34471 5015
rect 37841 4981 37875 5015
rect 39129 4981 39163 5015
rect 39773 4981 39807 5015
rect 40509 4981 40543 5015
rect 41245 4981 41279 5015
rect 45017 4981 45051 5015
rect 50169 4981 50203 5015
rect 11069 4777 11103 4811
rect 15393 4777 15427 4811
rect 21833 4777 21867 4811
rect 27537 4777 27571 4811
rect 27721 4777 27755 4811
rect 30481 4777 30515 4811
rect 37657 4777 37691 4811
rect 44189 4777 44223 4811
rect 45385 4777 45419 4811
rect 58265 4777 58299 4811
rect 8585 4709 8619 4743
rect 10885 4709 10919 4743
rect 13553 4709 13587 4743
rect 14565 4709 14599 4743
rect 14749 4709 14783 4743
rect 32137 4709 32171 4743
rect 9597 4641 9631 4675
rect 9781 4641 9815 4675
rect 9965 4641 9999 4675
rect 10609 4641 10643 4675
rect 12817 4641 12851 4675
rect 17785 4641 17819 4675
rect 21005 4641 21039 4675
rect 21189 4641 21223 4675
rect 23857 4641 23891 4675
rect 26709 4641 26743 4675
rect 32689 4641 32723 4675
rect 38853 4641 38887 4675
rect 41705 4641 41739 4675
rect 42441 4641 42475 4675
rect 42625 4641 42659 4675
rect 9873 4573 9907 4607
rect 10057 4573 10091 4607
rect 12081 4573 12115 4607
rect 13277 4573 13311 4607
rect 14289 4573 14323 4607
rect 15301 4573 15335 4607
rect 16129 4573 16163 4607
rect 16589 4573 16623 4607
rect 17509 4573 17543 4607
rect 18429 4573 18463 4607
rect 19625 4573 19659 4607
rect 21741 4573 21775 4607
rect 22385 4573 22419 4607
rect 24685 4573 24719 4607
rect 26433 4573 26467 4607
rect 26525 4573 26559 4607
rect 27169 4573 27203 4607
rect 28549 4573 28583 4607
rect 29837 4573 29871 4607
rect 30481 4573 30515 4607
rect 30665 4573 30699 4607
rect 32597 4573 32631 4607
rect 33333 4573 33367 4607
rect 33517 4573 33551 4607
rect 35541 4573 35575 4607
rect 35808 4573 35842 4607
rect 38301 4573 38335 4607
rect 40877 4573 40911 4607
rect 42349 4573 42383 4607
rect 42717 4573 42751 4607
rect 43637 4573 43671 4607
rect 43821 4573 43855 4607
rect 44010 4573 44044 4607
rect 46213 4573 46247 4607
rect 51273 4573 51307 4607
rect 51457 4573 51491 4607
rect 58081 4573 58115 4607
rect 6929 4505 6963 4539
rect 7665 4505 7699 4539
rect 8401 4505 8435 4539
rect 11897 4505 11931 4539
rect 12633 4505 12667 4539
rect 16865 4505 16899 4539
rect 18705 4505 18739 4539
rect 19901 4505 19935 4539
rect 20913 4505 20947 4539
rect 22661 4505 22695 4539
rect 23673 4505 23707 4539
rect 25053 4505 25087 4539
rect 27583 4505 27617 4539
rect 28917 4505 28951 4539
rect 32505 4505 32539 4539
rect 37565 4505 37599 4539
rect 40141 4505 40175 4539
rect 43913 4505 43947 4539
rect 45293 4505 45327 4539
rect 46029 4505 46063 4539
rect 7021 4437 7055 4471
rect 7757 4437 7791 4471
rect 13737 4437 13771 4471
rect 20545 4437 20579 4471
rect 23305 4437 23339 4471
rect 23765 4437 23799 4471
rect 29929 4437 29963 4471
rect 33701 4437 33735 4471
rect 36921 4437 36955 4471
rect 40233 4437 40267 4471
rect 40969 4437 41003 4471
rect 51641 4437 51675 4471
rect 24685 4233 24719 4267
rect 26433 4233 26467 4267
rect 32689 4233 32723 4267
rect 53113 4233 53147 4267
rect 5825 4165 5859 4199
rect 6653 4165 6687 4199
rect 7389 4165 7423 4199
rect 10977 4165 11011 4199
rect 11805 4165 11839 4199
rect 13369 4165 13403 4199
rect 14289 4165 14323 4199
rect 20260 4165 20294 4199
rect 27620 4165 27654 4199
rect 30757 4165 30791 4199
rect 41337 4165 41371 4199
rect 44465 4165 44499 4199
rect 46857 4165 46891 4199
rect 52193 4165 52227 4199
rect 53021 4165 53055 4199
rect 53757 4165 53791 4199
rect 58173 4165 58207 4199
rect 1593 4097 1627 4131
rect 6837 4097 6871 4131
rect 8033 4097 8067 4131
rect 9321 4097 9355 4131
rect 11161 4097 11195 4131
rect 11989 4097 12023 4131
rect 15853 4097 15887 4131
rect 16957 4097 16991 4131
rect 17877 4097 17911 4131
rect 19165 4097 19199 4131
rect 22385 4097 22419 4131
rect 23572 4097 23606 4131
rect 25145 4097 25179 4131
rect 29745 4097 29779 4131
rect 31585 4097 31619 4131
rect 33517 4097 33551 4131
rect 34437 4097 34471 4131
rect 35357 4097 35391 4131
rect 36277 4097 36311 4131
rect 37473 4097 37507 4131
rect 38844 4097 38878 4131
rect 40601 4097 40635 4131
rect 41521 4097 41555 4131
rect 43361 4097 43395 4131
rect 43729 4097 43763 4131
rect 45201 4097 45235 4131
rect 45937 4097 45971 4131
rect 46673 4097 46707 4131
rect 48237 4097 48271 4131
rect 53941 4097 53975 4131
rect 54585 4097 54619 4131
rect 58357 4097 58391 4131
rect 1777 4029 1811 4063
rect 8493 4029 8527 4063
rect 9137 4029 9171 4063
rect 9229 4029 9263 4063
rect 9413 4029 9447 4063
rect 9965 4029 9999 4063
rect 10425 4029 10459 4063
rect 12449 4029 12483 4063
rect 12909 4029 12943 4063
rect 14749 4029 14783 4063
rect 16129 4029 16163 4063
rect 17233 4029 17267 4063
rect 18153 4029 18187 4063
rect 19257 4029 19291 4063
rect 19349 4029 19383 4063
rect 19993 4029 20027 4063
rect 22661 4029 22695 4063
rect 23305 4029 23339 4063
rect 25329 4029 25363 4063
rect 27353 4029 27387 4063
rect 29929 4029 29963 4063
rect 32781 4029 32815 4063
rect 32873 4029 32907 4063
rect 33701 4029 33735 4063
rect 34621 4029 34655 4063
rect 35541 4029 35575 4063
rect 36461 4029 36495 4063
rect 37657 4029 37691 4063
rect 38577 4029 38611 4063
rect 40785 4029 40819 4063
rect 43453 4029 43487 4063
rect 43637 4029 43671 4063
rect 44649 4029 44683 4063
rect 45385 4029 45419 4063
rect 46121 4029 46155 4063
rect 6009 3961 6043 3995
rect 8401 3961 8435 3995
rect 10241 3961 10275 3995
rect 12817 3961 12851 3995
rect 13645 3961 13679 3995
rect 14565 3961 14599 3995
rect 31769 3961 31803 3995
rect 39957 3961 39991 3995
rect 42993 3961 43027 3995
rect 48421 3961 48455 3995
rect 54769 3961 54803 3995
rect 7481 3893 7515 3927
rect 8953 3893 8987 3927
rect 13829 3893 13863 3927
rect 18797 3893 18831 3927
rect 21373 3893 21407 3927
rect 28733 3893 28767 3927
rect 30849 3893 30883 3927
rect 32321 3893 32355 3927
rect 52285 3893 52319 3927
rect 5181 3689 5215 3723
rect 10885 3689 10919 3723
rect 12817 3689 12851 3723
rect 13737 3689 13771 3723
rect 16129 3689 16163 3723
rect 24593 3689 24627 3723
rect 27721 3689 27755 3723
rect 33701 3689 33735 3723
rect 42901 3689 42935 3723
rect 46121 3689 46155 3723
rect 47041 3689 47075 3723
rect 47961 3689 47995 3723
rect 48697 3689 48731 3723
rect 49433 3689 49467 3723
rect 53481 3689 53515 3723
rect 54217 3689 54251 3723
rect 55689 3689 55723 3723
rect 6009 3621 6043 3655
rect 7573 3621 7607 3655
rect 7665 3621 7699 3655
rect 8401 3621 8435 3655
rect 8585 3621 8619 3655
rect 10701 3621 10735 3655
rect 11897 3621 11931 3655
rect 12633 3621 12667 3655
rect 13645 3621 13679 3655
rect 15945 3621 15979 3655
rect 21005 3621 21039 3655
rect 38669 3621 38703 3655
rect 41981 3621 42015 3655
rect 50629 3621 50663 3655
rect 6745 3553 6779 3587
rect 9413 3553 9447 3587
rect 9689 3553 9723 3587
rect 17785 3553 17819 3587
rect 22109 3553 22143 3587
rect 25053 3553 25087 3587
rect 25237 3553 25271 3587
rect 28365 3553 28399 3587
rect 32321 3553 32355 3587
rect 32597 3553 32631 3587
rect 35081 3553 35115 3587
rect 37289 3553 37323 3587
rect 40141 3553 40175 3587
rect 40877 3553 40911 3587
rect 41061 3553 41095 3587
rect 51365 3553 51399 3587
rect 52837 3553 52871 3587
rect 56885 3553 56919 3587
rect 1593 3485 1627 3519
rect 5089 3485 5123 3519
rect 9597 3485 9631 3519
rect 9781 3485 9815 3519
rect 9873 3485 9907 3519
rect 10425 3485 10459 3519
rect 11713 3485 11747 3519
rect 14749 3485 14783 3519
rect 15669 3485 15703 3519
rect 17049 3485 17083 3519
rect 17509 3485 17543 3519
rect 18429 3485 18463 3519
rect 19625 3485 19659 3519
rect 22661 3485 22695 3519
rect 24961 3485 24995 3519
rect 25789 3485 25823 3519
rect 26893 3485 26927 3519
rect 27005 3485 27039 3519
rect 29193 3485 29227 3519
rect 30297 3485 30331 3519
rect 31585 3485 31619 3519
rect 31677 3485 31711 3519
rect 34897 3485 34931 3519
rect 36185 3485 36219 3519
rect 37565 3485 37599 3519
rect 40785 3485 40819 3519
rect 41153 3485 41187 3519
rect 41797 3485 41831 3519
rect 43257 3485 43291 3519
rect 43545 3485 43579 3519
rect 43658 3485 43692 3519
rect 43913 3485 43947 3519
rect 44189 3485 44223 3519
rect 45293 3485 45327 3519
rect 48513 3485 48547 3519
rect 49249 3485 49283 3519
rect 52653 3485 52687 3519
rect 54125 3485 54159 3519
rect 55505 3485 55539 3519
rect 1869 3417 1903 3451
rect 5825 3417 5859 3451
rect 6561 3417 6595 3451
rect 7205 3417 7239 3451
rect 8125 3417 8159 3451
rect 12357 3417 12391 3451
rect 13277 3417 13311 3451
rect 15025 3417 15059 3451
rect 18705 3417 18739 3451
rect 19881 3417 19915 3451
rect 21833 3417 21867 3451
rect 22928 3417 22962 3451
rect 26065 3417 26099 3451
rect 26709 3417 26743 3451
rect 27095 3417 27129 3451
rect 27261 3417 27295 3451
rect 28181 3417 28215 3451
rect 29009 3417 29043 3451
rect 30573 3417 30607 3451
rect 31861 3417 31895 3451
rect 36737 3417 36771 3451
rect 46029 3417 46063 3451
rect 46949 3417 46983 3451
rect 47869 3417 47903 3451
rect 50445 3417 50479 3451
rect 51181 3417 51215 3451
rect 51917 3417 51951 3451
rect 53389 3417 53423 3451
rect 57130 3417 57164 3451
rect 21465 3349 21499 3383
rect 21925 3349 21959 3383
rect 24041 3349 24075 3383
rect 28089 3349 28123 3383
rect 45385 3349 45419 3383
rect 52009 3349 52043 3383
rect 58265 3349 58299 3383
rect 8953 3145 8987 3179
rect 10885 3145 10919 3179
rect 13001 3145 13035 3179
rect 23213 3145 23247 3179
rect 24593 3145 24627 3179
rect 36921 3145 36955 3179
rect 37841 3145 37875 3179
rect 38209 3145 38243 3179
rect 44465 3145 44499 3179
rect 45201 3145 45235 3179
rect 46489 3145 46523 3179
rect 47961 3145 47995 3179
rect 48881 3145 48915 3179
rect 49801 3145 49835 3179
rect 50721 3145 50755 3179
rect 52193 3145 52227 3179
rect 55321 3145 55355 3179
rect 4353 3077 4387 3111
rect 10425 3077 10459 3111
rect 18981 3077 19015 3111
rect 19892 3077 19926 3111
rect 23673 3077 23707 3111
rect 36553 3077 36587 3111
rect 36645 3077 36679 3111
rect 40417 3077 40451 3111
rect 45109 3077 45143 3111
rect 50629 3077 50663 3111
rect 52101 3077 52135 3111
rect 54493 3077 54527 3111
rect 58173 3077 58207 3111
rect 1593 3009 1627 3043
rect 4537 3009 4571 3043
rect 5089 3009 5123 3043
rect 5825 3009 5859 3043
rect 7113 3009 7147 3043
rect 7849 3009 7883 3043
rect 9597 3009 9631 3043
rect 9689 3009 9723 3043
rect 9873 3009 9907 3043
rect 12173 3009 12207 3043
rect 12909 3009 12943 3043
rect 13553 3009 13587 3043
rect 14473 3009 14507 3043
rect 15393 3009 15427 3043
rect 16865 3009 16899 3043
rect 17785 3009 17819 3043
rect 18705 3009 18739 3043
rect 19625 3009 19659 3043
rect 22293 3009 22327 3043
rect 23581 3009 23615 3043
rect 25237 3009 25271 3043
rect 26157 3009 26191 3043
rect 27537 3009 27571 3043
rect 28457 3009 28491 3043
rect 30849 3009 30883 3043
rect 32321 3009 32355 3043
rect 33241 3009 33275 3043
rect 34897 3009 34931 3043
rect 35357 3009 35391 3043
rect 36277 3009 36311 3043
rect 36425 3009 36459 3043
rect 36742 3009 36776 3043
rect 39037 3009 39071 3043
rect 40049 3009 40083 3043
rect 40969 3009 41003 3043
rect 41153 3009 41187 3043
rect 41705 3009 41739 3043
rect 42073 3009 42107 3043
rect 42625 3009 42659 3043
rect 43269 3009 43303 3043
rect 43637 3009 43671 3043
rect 44281 3009 44315 3043
rect 46397 3009 46431 3043
rect 47869 3009 47903 3043
rect 48789 3009 48823 3043
rect 49709 3009 49743 3043
rect 51365 3009 51399 3043
rect 53021 3009 53055 3043
rect 54125 3009 54159 3043
rect 55045 3009 55079 3043
rect 55873 3009 55907 3043
rect 57253 3009 57287 3043
rect 1777 2941 1811 2975
rect 8493 2941 8527 2975
rect 9772 2941 9806 2975
rect 13829 2941 13863 2975
rect 14749 2941 14783 2975
rect 17141 2941 17175 2975
rect 18061 2941 18095 2975
rect 22569 2941 22603 2975
rect 23765 2941 23799 2975
rect 25421 2941 25455 2975
rect 26433 2941 26467 2975
rect 27813 2941 27847 2975
rect 28733 2941 28767 2975
rect 29837 2941 29871 2975
rect 31033 2941 31067 2975
rect 32505 2941 32539 2975
rect 33517 2941 33551 2975
rect 35541 2941 35575 2975
rect 38301 2941 38335 2975
rect 38485 2941 38519 2975
rect 39221 2941 39255 2975
rect 43361 2941 43395 2975
rect 43545 2941 43579 2975
rect 51549 2941 51583 2975
rect 56057 2941 56091 2975
rect 57069 2941 57103 2975
rect 58357 2941 58391 2975
rect 5273 2873 5307 2907
rect 8769 2873 8803 2907
rect 10701 2873 10735 2907
rect 12357 2873 12391 2907
rect 15669 2873 15703 2907
rect 53205 2873 53239 2907
rect 57437 2873 57471 2907
rect 5917 2805 5951 2839
rect 7205 2805 7239 2839
rect 7941 2805 7975 2839
rect 9413 2805 9447 2839
rect 15853 2805 15887 2839
rect 21005 2805 21039 2839
rect 3341 2601 3375 2635
rect 11897 2601 11931 2635
rect 14473 2601 14507 2635
rect 45385 2601 45419 2635
rect 46213 2601 46247 2635
rect 47133 2601 47167 2635
rect 47961 2601 47995 2635
rect 48881 2601 48915 2635
rect 58265 2601 58299 2635
rect 6009 2533 6043 2567
rect 9689 2533 9723 2567
rect 10425 2533 10459 2567
rect 11161 2533 11195 2567
rect 50629 2533 50663 2567
rect 52101 2533 52135 2567
rect 15209 2465 15243 2499
rect 17049 2465 17083 2499
rect 18705 2465 18739 2499
rect 20177 2465 20211 2499
rect 22937 2465 22971 2499
rect 28089 2465 28123 2499
rect 32505 2465 32539 2499
rect 36001 2465 36035 2499
rect 37657 2465 37691 2499
rect 38577 2465 38611 2499
rect 41337 2465 41371 2499
rect 54033 2465 54067 2499
rect 55689 2465 55723 2499
rect 1593 2397 1627 2431
rect 3249 2397 3283 2431
rect 5273 2397 5307 2431
rect 6929 2397 6963 2431
rect 10241 2397 10275 2431
rect 10977 2397 11011 2431
rect 12357 2397 12391 2431
rect 13277 2397 13311 2431
rect 14933 2397 14967 2431
rect 15853 2397 15887 2431
rect 17509 2397 17543 2431
rect 18429 2397 18463 2431
rect 19901 2397 19935 2431
rect 20729 2397 20763 2431
rect 21005 2397 21039 2431
rect 22661 2397 22695 2431
rect 23581 2397 23615 2431
rect 25237 2397 25271 2431
rect 26157 2397 26191 2431
rect 27813 2397 27847 2431
rect 28733 2397 28767 2431
rect 30205 2397 30239 2431
rect 31125 2397 31159 2431
rect 32321 2397 32355 2431
rect 33241 2397 33275 2431
rect 34897 2397 34931 2431
rect 35817 2397 35851 2431
rect 37473 2397 37507 2431
rect 38393 2397 38427 2431
rect 41061 2397 41095 2431
rect 42625 2397 42659 2431
rect 42773 2397 42807 2431
rect 42901 2397 42935 2431
rect 43131 2397 43165 2431
rect 45201 2397 45235 2431
rect 47869 2397 47903 2431
rect 50445 2397 50479 2431
rect 51181 2397 51215 2431
rect 53849 2397 53883 2431
rect 55505 2397 55539 2431
rect 57069 2397 57103 2431
rect 58173 2397 58207 2431
rect 1869 2329 1903 2363
rect 4353 2329 4387 2363
rect 5089 2329 5123 2363
rect 5825 2329 5859 2363
rect 7665 2329 7699 2363
rect 8401 2329 8435 2363
rect 9505 2329 9539 2363
rect 12633 2329 12667 2363
rect 13553 2329 13587 2363
rect 16129 2329 16163 2363
rect 17785 2329 17819 2363
rect 21281 2329 21315 2363
rect 23857 2329 23891 2363
rect 25513 2329 25547 2363
rect 26433 2329 26467 2363
rect 29009 2329 29043 2363
rect 30481 2329 30515 2363
rect 31401 2329 31435 2363
rect 33517 2329 33551 2363
rect 35173 2329 35207 2363
rect 40141 2329 40175 2363
rect 42993 2329 43027 2363
rect 43913 2329 43947 2363
rect 46121 2329 46155 2363
rect 47041 2329 47075 2363
rect 48789 2329 48823 2363
rect 51917 2329 51951 2363
rect 53021 2329 53055 2363
rect 57345 2329 57379 2363
rect 4445 2261 4479 2295
rect 7021 2261 7055 2295
rect 7757 2261 7791 2295
rect 8493 2261 8527 2295
rect 19441 2261 19475 2295
rect 22017 2261 22051 2295
rect 24593 2261 24627 2295
rect 27169 2261 27203 2295
rect 40233 2261 40267 2295
rect 43269 2261 43303 2295
rect 44005 2261 44039 2295
rect 51273 2261 51307 2295
rect 53113 2261 53147 2295
<< metal1 >>
rect 30098 61752 30104 61804
rect 30156 61792 30162 61804
rect 49418 61792 49424 61804
rect 30156 61764 49424 61792
rect 30156 61752 30162 61764
rect 49418 61752 49424 61764
rect 49476 61752 49482 61804
rect 33410 61684 33416 61736
rect 33468 61724 33474 61736
rect 42702 61724 42708 61736
rect 33468 61696 42708 61724
rect 33468 61684 33474 61696
rect 42702 61684 42708 61696
rect 42760 61684 42766 61736
rect 11054 61616 11060 61668
rect 11112 61656 11118 61668
rect 19426 61656 19432 61668
rect 11112 61628 19432 61656
rect 11112 61616 11118 61628
rect 19426 61616 19432 61628
rect 19484 61616 19490 61668
rect 28442 61616 28448 61668
rect 28500 61656 28506 61668
rect 46842 61656 46848 61668
rect 28500 61628 46848 61656
rect 28500 61616 28506 61628
rect 46842 61616 46848 61628
rect 46900 61616 46906 61668
rect 21174 61548 21180 61600
rect 21232 61588 21238 61600
rect 40218 61588 40224 61600
rect 21232 61560 40224 61588
rect 21232 61548 21238 61560
rect 40218 61548 40224 61560
rect 40276 61548 40282 61600
rect 41874 61548 41880 61600
rect 41932 61588 41938 61600
rect 51442 61588 51448 61600
rect 41932 61560 51448 61588
rect 41932 61548 41938 61560
rect 51442 61548 51448 61560
rect 51500 61548 51506 61600
rect 1104 61498 58880 61520
rect 1104 61446 4214 61498
rect 4266 61446 4278 61498
rect 4330 61446 4342 61498
rect 4394 61446 4406 61498
rect 4458 61446 4470 61498
rect 4522 61446 34934 61498
rect 34986 61446 34998 61498
rect 35050 61446 35062 61498
rect 35114 61446 35126 61498
rect 35178 61446 35190 61498
rect 35242 61446 58880 61498
rect 1104 61424 58880 61446
rect 7650 61344 7656 61396
rect 7708 61384 7714 61396
rect 40218 61384 40224 61396
rect 7708 61356 39804 61384
rect 40179 61356 40224 61384
rect 7708 61344 7714 61356
rect 9677 61319 9735 61325
rect 9677 61285 9689 61319
rect 9723 61316 9735 61319
rect 15838 61316 15844 61328
rect 9723 61288 15844 61316
rect 9723 61285 9735 61288
rect 9677 61279 9735 61285
rect 15838 61276 15844 61288
rect 15896 61276 15902 61328
rect 18230 61316 18236 61328
rect 16546 61288 18236 61316
rect 3053 61251 3111 61257
rect 3053 61217 3065 61251
rect 3099 61248 3111 61251
rect 10413 61251 10471 61257
rect 3099 61220 10364 61248
rect 3099 61217 3111 61220
rect 3053 61211 3111 61217
rect 1670 61180 1676 61192
rect 1631 61152 1676 61180
rect 1670 61140 1676 61152
rect 1728 61140 1734 61192
rect 2774 61180 2780 61192
rect 2735 61152 2780 61180
rect 2774 61140 2780 61152
rect 2832 61140 2838 61192
rect 4341 61183 4399 61189
rect 4341 61149 4353 61183
rect 4387 61180 4399 61183
rect 4614 61180 4620 61192
rect 4387 61152 4620 61180
rect 4387 61149 4399 61152
rect 4341 61143 4399 61149
rect 4614 61140 4620 61152
rect 4672 61140 4678 61192
rect 5074 61180 5080 61192
rect 5035 61152 5080 61180
rect 5074 61140 5080 61152
rect 5132 61140 5138 61192
rect 5718 61180 5724 61192
rect 5679 61152 5724 61180
rect 5718 61140 5724 61152
rect 5776 61140 5782 61192
rect 6638 61180 6644 61192
rect 6599 61152 6644 61180
rect 6638 61140 6644 61152
rect 6696 61140 6702 61192
rect 7558 61180 7564 61192
rect 7519 61152 7564 61180
rect 7558 61140 7564 61152
rect 7616 61140 7622 61192
rect 9493 61183 9551 61189
rect 9493 61149 9505 61183
rect 9539 61180 9551 61183
rect 9674 61180 9680 61192
rect 9539 61152 9680 61180
rect 9539 61149 9551 61152
rect 9493 61143 9551 61149
rect 9674 61140 9680 61152
rect 9732 61140 9738 61192
rect 10226 61180 10232 61192
rect 10187 61152 10232 61180
rect 10226 61140 10232 61152
rect 10284 61140 10290 61192
rect 2225 61115 2283 61121
rect 2225 61081 2237 61115
rect 2271 61081 2283 61115
rect 2225 61075 2283 61081
rect 4525 61115 4583 61121
rect 4525 61081 4537 61115
rect 4571 61112 4583 61115
rect 5626 61112 5632 61124
rect 4571 61084 5632 61112
rect 4571 61081 4583 61084
rect 4525 61075 4583 61081
rect 2240 61044 2268 61075
rect 5626 61072 5632 61084
rect 5684 61072 5690 61124
rect 6914 61072 6920 61124
rect 6972 61112 6978 61124
rect 7837 61115 7895 61121
rect 6972 61084 7017 61112
rect 6972 61072 6978 61084
rect 7837 61081 7849 61115
rect 7883 61112 7895 61115
rect 8938 61112 8944 61124
rect 7883 61084 8944 61112
rect 7883 61081 7895 61084
rect 7837 61075 7895 61081
rect 8938 61072 8944 61084
rect 8996 61072 9002 61124
rect 10336 61112 10364 61220
rect 10413 61217 10425 61251
rect 10459 61248 10471 61251
rect 16546 61248 16574 61288
rect 18230 61276 18236 61288
rect 18288 61276 18294 61328
rect 20717 61319 20775 61325
rect 20717 61285 20729 61319
rect 20763 61316 20775 61319
rect 22094 61316 22100 61328
rect 20763 61288 22100 61316
rect 20763 61285 20775 61288
rect 20717 61279 20775 61285
rect 22094 61276 22100 61288
rect 22152 61276 22158 61328
rect 38473 61319 38531 61325
rect 38473 61316 38485 61319
rect 26206 61288 38485 61316
rect 10459 61220 16574 61248
rect 18141 61251 18199 61257
rect 10459 61217 10471 61220
rect 10413 61211 10471 61217
rect 18141 61217 18153 61251
rect 18187 61248 18199 61251
rect 22830 61248 22836 61260
rect 18187 61220 22836 61248
rect 18187 61217 18199 61220
rect 18141 61211 18199 61217
rect 22830 61208 22836 61220
rect 22888 61208 22894 61260
rect 26206 61248 26234 61288
rect 38473 61285 38485 61288
rect 38519 61285 38531 61319
rect 39776 61316 39804 61356
rect 40218 61344 40224 61356
rect 40276 61344 40282 61396
rect 42610 61344 42616 61396
rect 42668 61384 42674 61396
rect 46842 61384 46848 61396
rect 42668 61356 45554 61384
rect 46803 61356 46848 61384
rect 42668 61344 42674 61356
rect 43717 61319 43775 61325
rect 43717 61316 43729 61319
rect 39776 61288 43729 61316
rect 38473 61279 38531 61285
rect 43717 61285 43729 61288
rect 43763 61285 43775 61319
rect 45526 61316 45554 61356
rect 46842 61344 46848 61356
rect 46900 61344 46906 61396
rect 49418 61384 49424 61396
rect 49379 61356 49424 61384
rect 49418 61344 49424 61356
rect 49476 61344 49482 61396
rect 51442 61384 51448 61396
rect 51403 61356 51448 61384
rect 51442 61344 51448 61356
rect 51500 61344 51506 61396
rect 52273 61319 52331 61325
rect 52273 61316 52285 61319
rect 45526 61288 52285 61316
rect 43717 61279 43775 61285
rect 52273 61285 52285 61288
rect 52319 61285 52331 61319
rect 52273 61279 52331 61285
rect 23676 61220 26234 61248
rect 10965 61183 11023 61189
rect 10965 61149 10977 61183
rect 11011 61180 11023 61183
rect 11146 61180 11152 61192
rect 11011 61152 11152 61180
rect 11011 61149 11023 61152
rect 10965 61143 11023 61149
rect 11146 61140 11152 61152
rect 11204 61140 11210 61192
rect 11974 61180 11980 61192
rect 11935 61152 11980 61180
rect 11974 61140 11980 61152
rect 12032 61140 12038 61192
rect 12710 61180 12716 61192
rect 12671 61152 12716 61180
rect 12710 61140 12716 61152
rect 12768 61140 12774 61192
rect 12986 61180 12992 61192
rect 12947 61152 12992 61180
rect 12986 61140 12992 61152
rect 13044 61140 13050 61192
rect 14918 61180 14924 61192
rect 14879 61152 14924 61180
rect 14918 61140 14924 61152
rect 14976 61140 14982 61192
rect 16114 61180 16120 61192
rect 16075 61152 16120 61180
rect 16114 61140 16120 61152
rect 16172 61140 16178 61192
rect 17218 61180 17224 61192
rect 17179 61152 17224 61180
rect 17218 61140 17224 61152
rect 17276 61140 17282 61192
rect 17954 61180 17960 61192
rect 17915 61152 17960 61180
rect 17954 61140 17960 61152
rect 18012 61140 18018 61192
rect 18690 61180 18696 61192
rect 18651 61152 18696 61180
rect 18690 61140 18696 61152
rect 18748 61140 18754 61192
rect 19794 61180 19800 61192
rect 19755 61152 19800 61180
rect 19794 61140 19800 61152
rect 19852 61140 19858 61192
rect 20533 61183 20591 61189
rect 20533 61149 20545 61183
rect 20579 61180 20591 61183
rect 20714 61180 20720 61192
rect 20579 61152 20720 61180
rect 20579 61149 20591 61152
rect 20533 61143 20591 61149
rect 20714 61140 20720 61152
rect 20772 61140 20778 61192
rect 21266 61180 21272 61192
rect 21227 61152 21272 61180
rect 21266 61140 21272 61152
rect 21324 61140 21330 61192
rect 22370 61180 22376 61192
rect 22331 61152 22376 61180
rect 22370 61140 22376 61152
rect 22428 61140 22434 61192
rect 23676 61180 23704 61220
rect 35894 61208 35900 61260
rect 35952 61248 35958 61260
rect 35952 61220 36492 61248
rect 35952 61208 35958 61220
rect 23842 61180 23848 61192
rect 22572 61152 23704 61180
rect 23803 61152 23848 61180
rect 14642 61112 14648 61124
rect 10336 61084 14648 61112
rect 14642 61072 14648 61084
rect 14700 61072 14706 61124
rect 15194 61112 15200 61124
rect 15155 61084 15200 61112
rect 15194 61072 15200 61084
rect 15252 61072 15258 61124
rect 16301 61115 16359 61121
rect 16301 61081 16313 61115
rect 16347 61112 16359 61115
rect 17402 61112 17408 61124
rect 16347 61084 17408 61112
rect 16347 61081 16359 61084
rect 16301 61075 16359 61081
rect 17402 61072 17408 61084
rect 17460 61072 17466 61124
rect 18874 61112 18880 61124
rect 18835 61084 18880 61112
rect 18874 61072 18880 61084
rect 18932 61072 18938 61124
rect 19981 61115 20039 61121
rect 19981 61081 19993 61115
rect 20027 61112 20039 61115
rect 20438 61112 20444 61124
rect 20027 61084 20444 61112
rect 20027 61081 20039 61084
rect 19981 61075 20039 61081
rect 20438 61072 20444 61084
rect 20496 61072 20502 61124
rect 21082 61072 21088 61124
rect 21140 61112 21146 61124
rect 22572 61112 22600 61152
rect 23842 61140 23848 61152
rect 23900 61140 23906 61192
rect 25130 61140 25136 61192
rect 25188 61180 25194 61192
rect 25317 61183 25375 61189
rect 25317 61180 25329 61183
rect 25188 61152 25329 61180
rect 25188 61140 25194 61152
rect 25317 61149 25329 61152
rect 25363 61149 25375 61183
rect 25317 61143 25375 61149
rect 26234 61140 26240 61192
rect 26292 61180 26298 61192
rect 26292 61152 26337 61180
rect 26292 61140 26298 61152
rect 26602 61140 26608 61192
rect 26660 61180 26666 61192
rect 27249 61183 27307 61189
rect 27249 61180 27261 61183
rect 26660 61152 27261 61180
rect 26660 61140 26666 61152
rect 27249 61149 27261 61152
rect 27295 61149 27307 61183
rect 27249 61143 27307 61149
rect 28074 61140 28080 61192
rect 28132 61180 28138 61192
rect 28261 61183 28319 61189
rect 28261 61180 28273 61183
rect 28132 61152 28273 61180
rect 28132 61140 28138 61152
rect 28261 61149 28273 61152
rect 28307 61149 28319 61183
rect 29822 61180 29828 61192
rect 29783 61152 29828 61180
rect 28261 61143 28319 61149
rect 29822 61140 29828 61152
rect 29880 61140 29886 61192
rect 31202 61180 31208 61192
rect 31163 61152 31208 61180
rect 31202 61140 31208 61152
rect 31260 61140 31266 61192
rect 31754 61140 31760 61192
rect 31812 61180 31818 61192
rect 32401 61183 32459 61189
rect 32401 61180 32413 61183
rect 31812 61152 32413 61180
rect 31812 61140 31818 61152
rect 32401 61149 32413 61152
rect 32447 61149 32459 61183
rect 32401 61143 32459 61149
rect 32858 61140 32864 61192
rect 32916 61180 32922 61192
rect 33321 61183 33379 61189
rect 33321 61180 33333 61183
rect 32916 61152 33333 61180
rect 32916 61140 32922 61152
rect 33321 61149 33333 61152
rect 33367 61149 33379 61183
rect 33321 61143 33379 61149
rect 33502 61140 33508 61192
rect 33560 61180 33566 61192
rect 34057 61183 34115 61189
rect 34057 61180 34069 61183
rect 33560 61152 34069 61180
rect 33560 61140 33566 61152
rect 34057 61149 34069 61152
rect 34103 61149 34115 61183
rect 34057 61143 34115 61149
rect 34698 61140 34704 61192
rect 34756 61180 34762 61192
rect 36464 61189 36492 61220
rect 41506 61208 41512 61260
rect 41564 61248 41570 61260
rect 48041 61251 48099 61257
rect 48041 61248 48053 61251
rect 41564 61220 48053 61248
rect 41564 61208 41570 61220
rect 48041 61217 48053 61220
rect 48087 61217 48099 61251
rect 53374 61248 53380 61260
rect 53335 61220 53380 61248
rect 48041 61211 48099 61217
rect 53374 61208 53380 61220
rect 53432 61208 53438 61260
rect 35713 61183 35771 61189
rect 35713 61180 35725 61183
rect 34756 61152 35725 61180
rect 34756 61140 34762 61152
rect 35713 61149 35725 61152
rect 35759 61149 35771 61183
rect 35713 61143 35771 61149
rect 36449 61183 36507 61189
rect 36449 61149 36461 61183
rect 36495 61149 36507 61183
rect 36449 61143 36507 61149
rect 37274 61140 37280 61192
rect 37332 61180 37338 61192
rect 37553 61183 37611 61189
rect 37553 61180 37565 61183
rect 37332 61152 37565 61180
rect 37332 61140 37338 61152
rect 37553 61149 37565 61152
rect 37599 61149 37611 61183
rect 37553 61143 37611 61149
rect 37642 61140 37648 61192
rect 37700 61180 37706 61192
rect 38289 61183 38347 61189
rect 38289 61180 38301 61183
rect 37700 61152 38301 61180
rect 37700 61140 37706 61152
rect 38289 61149 38301 61152
rect 38335 61149 38347 61183
rect 38289 61143 38347 61149
rect 38654 61140 38660 61192
rect 38712 61180 38718 61192
rect 38933 61183 38991 61189
rect 38933 61180 38945 61183
rect 38712 61152 38945 61180
rect 38712 61140 38718 61152
rect 38933 61149 38945 61152
rect 38979 61149 38991 61183
rect 38933 61143 38991 61149
rect 39482 61140 39488 61192
rect 39540 61180 39546 61192
rect 40129 61183 40187 61189
rect 40129 61180 40141 61183
rect 39540 61152 40141 61180
rect 39540 61140 39546 61152
rect 40129 61149 40141 61152
rect 40175 61149 40187 61183
rect 40129 61143 40187 61149
rect 40586 61140 40592 61192
rect 40644 61180 40650 61192
rect 41601 61183 41659 61189
rect 41601 61180 41613 61183
rect 40644 61152 41613 61180
rect 40644 61140 40650 61152
rect 41601 61149 41613 61152
rect 41647 61149 41659 61183
rect 41601 61143 41659 61149
rect 42058 61140 42064 61192
rect 42116 61180 42122 61192
rect 42613 61183 42671 61189
rect 42613 61180 42625 61183
rect 42116 61152 42625 61180
rect 42116 61140 42122 61152
rect 42613 61149 42625 61152
rect 42659 61149 42671 61183
rect 42613 61143 42671 61149
rect 42794 61140 42800 61192
rect 42852 61180 42858 61192
rect 43533 61183 43591 61189
rect 43533 61180 43545 61183
rect 42852 61152 43545 61180
rect 42852 61140 42858 61152
rect 43533 61149 43545 61152
rect 43579 61149 43591 61183
rect 43533 61143 43591 61149
rect 43622 61140 43628 61192
rect 43680 61180 43686 61192
rect 44361 61183 44419 61189
rect 44361 61180 44373 61183
rect 43680 61152 44373 61180
rect 43680 61140 43686 61152
rect 44361 61149 44373 61152
rect 44407 61149 44419 61183
rect 44361 61143 44419 61149
rect 44542 61140 44548 61192
rect 44600 61180 44606 61192
rect 45281 61183 45339 61189
rect 45281 61180 45293 61183
rect 44600 61152 45293 61180
rect 44600 61140 44606 61152
rect 45281 61149 45293 61152
rect 45327 61149 45339 61183
rect 45281 61143 45339 61149
rect 45554 61140 45560 61192
rect 45612 61180 45618 61192
rect 46017 61183 46075 61189
rect 46017 61180 46029 61183
rect 45612 61152 46029 61180
rect 45612 61140 45618 61152
rect 46017 61149 46029 61152
rect 46063 61149 46075 61183
rect 46017 61143 46075 61149
rect 46106 61140 46112 61192
rect 46164 61180 46170 61192
rect 46753 61183 46811 61189
rect 46753 61180 46765 61183
rect 46164 61152 46765 61180
rect 46164 61140 46170 61152
rect 46753 61149 46765 61152
rect 46799 61149 46811 61183
rect 46753 61143 46811 61149
rect 47210 61140 47216 61192
rect 47268 61180 47274 61192
rect 47857 61183 47915 61189
rect 47857 61180 47869 61183
rect 47268 61152 47869 61180
rect 47268 61140 47274 61152
rect 47857 61149 47869 61152
rect 47903 61149 47915 61183
rect 47857 61143 47915 61149
rect 48314 61140 48320 61192
rect 48372 61180 48378 61192
rect 48593 61183 48651 61189
rect 48593 61180 48605 61183
rect 48372 61152 48605 61180
rect 48372 61140 48378 61152
rect 48593 61149 48605 61152
rect 48639 61149 48651 61183
rect 48593 61143 48651 61149
rect 48682 61140 48688 61192
rect 48740 61180 48746 61192
rect 49329 61183 49387 61189
rect 49329 61180 49341 61183
rect 48740 61152 49341 61180
rect 48740 61140 48746 61152
rect 49329 61149 49341 61152
rect 49375 61149 49387 61183
rect 49329 61143 49387 61149
rect 49694 61140 49700 61192
rect 49752 61180 49758 61192
rect 50433 61183 50491 61189
rect 50433 61180 50445 61183
rect 49752 61152 50445 61180
rect 49752 61140 49758 61152
rect 50433 61149 50445 61152
rect 50479 61149 50491 61183
rect 50433 61143 50491 61149
rect 51074 61140 51080 61192
rect 51132 61180 51138 61192
rect 51353 61183 51411 61189
rect 51353 61180 51365 61183
rect 51132 61152 51365 61180
rect 51132 61140 51138 61152
rect 51353 61149 51365 61152
rect 51399 61149 51411 61183
rect 51353 61143 51411 61149
rect 51626 61140 51632 61192
rect 51684 61180 51690 61192
rect 52089 61183 52147 61189
rect 52089 61180 52101 61183
rect 51684 61152 52101 61180
rect 51684 61140 51690 61152
rect 52089 61149 52101 61152
rect 52135 61149 52147 61183
rect 53190 61180 53196 61192
rect 53151 61152 53196 61180
rect 52089 61143 52147 61149
rect 53190 61140 53196 61152
rect 53248 61140 53254 61192
rect 54110 61180 54116 61192
rect 54071 61152 54116 61180
rect 54110 61140 54116 61152
rect 54168 61140 54174 61192
rect 55490 61180 55496 61192
rect 55451 61152 55496 61180
rect 55490 61140 55496 61152
rect 55548 61140 55554 61192
rect 56042 61140 56048 61192
rect 56100 61180 56106 61192
rect 56505 61183 56563 61189
rect 56505 61180 56517 61183
rect 56100 61152 56517 61180
rect 56100 61140 56106 61152
rect 56505 61149 56517 61152
rect 56551 61149 56563 61183
rect 56505 61143 56563 61149
rect 57514 61140 57520 61192
rect 57572 61180 57578 61192
rect 58161 61183 58219 61189
rect 58161 61180 58173 61183
rect 57572 61152 58173 61180
rect 57572 61140 57578 61152
rect 58161 61149 58173 61152
rect 58207 61149 58219 61183
rect 58161 61143 58219 61149
rect 22738 61112 22744 61124
rect 21140 61084 22600 61112
rect 22699 61084 22744 61112
rect 21140 61072 21146 61084
rect 22738 61072 22744 61084
rect 22796 61072 22802 61124
rect 24029 61115 24087 61121
rect 24029 61081 24041 61115
rect 24075 61112 24087 61115
rect 24762 61112 24768 61124
rect 24075 61084 24768 61112
rect 24075 61081 24087 61084
rect 24029 61075 24087 61081
rect 24762 61072 24768 61084
rect 24820 61072 24826 61124
rect 26421 61115 26479 61121
rect 26421 61081 26433 61115
rect 26467 61112 26479 61115
rect 28166 61112 28172 61124
rect 26467 61084 28172 61112
rect 26467 61081 26479 61084
rect 26421 61075 26479 61081
rect 28166 61072 28172 61084
rect 28224 61072 28230 61124
rect 33134 61072 33140 61124
rect 33192 61112 33198 61124
rect 34241 61115 34299 61121
rect 34241 61112 34253 61115
rect 33192 61084 34253 61112
rect 33192 61072 33198 61084
rect 34241 61081 34253 61084
rect 34287 61081 34299 61115
rect 34241 61075 34299 61081
rect 34514 61072 34520 61124
rect 34572 61112 34578 61124
rect 34977 61115 35035 61121
rect 34977 61112 34989 61115
rect 34572 61084 34989 61112
rect 34572 61072 34578 61084
rect 34977 61081 34989 61084
rect 35023 61081 35035 61115
rect 34977 61075 35035 61081
rect 35894 61072 35900 61124
rect 35952 61112 35958 61124
rect 37737 61115 37795 61121
rect 35952 61084 35997 61112
rect 35952 61072 35958 61084
rect 37737 61081 37749 61115
rect 37783 61112 37795 61115
rect 38010 61112 38016 61124
rect 37783 61084 38016 61112
rect 37783 61081 37795 61084
rect 37737 61075 37795 61081
rect 38010 61072 38016 61084
rect 38068 61072 38074 61124
rect 39942 61072 39948 61124
rect 40000 61112 40006 61124
rect 40865 61115 40923 61121
rect 40865 61112 40877 61115
rect 40000 61084 40877 61112
rect 40000 61072 40006 61084
rect 40865 61081 40877 61084
rect 40911 61081 40923 61115
rect 42886 61112 42892 61124
rect 42847 61084 42892 61112
rect 40865 61075 40923 61081
rect 42886 61072 42892 61084
rect 42944 61072 42950 61124
rect 55766 61112 55772 61124
rect 53208 61084 55214 61112
rect 55727 61084 55772 61112
rect 53208 61056 53236 61084
rect 4706 61044 4712 61056
rect 2240 61016 4712 61044
rect 4706 61004 4712 61016
rect 4764 61004 4770 61056
rect 5166 61044 5172 61056
rect 5127 61016 5172 61044
rect 5166 61004 5172 61016
rect 5224 61004 5230 61056
rect 5902 61044 5908 61056
rect 5863 61016 5908 61044
rect 5902 61004 5908 61016
rect 5960 61004 5966 61056
rect 11054 61044 11060 61056
rect 11015 61016 11060 61044
rect 11054 61004 11060 61016
rect 11112 61004 11118 61056
rect 12158 61044 12164 61056
rect 12119 61016 12164 61044
rect 12158 61004 12164 61016
rect 12216 61004 12222 61056
rect 17310 61044 17316 61056
rect 17271 61016 17316 61044
rect 17310 61004 17316 61016
rect 17368 61004 17374 61056
rect 20898 61004 20904 61056
rect 20956 61044 20962 61056
rect 21361 61047 21419 61053
rect 21361 61044 21373 61047
rect 20956 61016 21373 61044
rect 20956 61004 20962 61016
rect 21361 61013 21373 61016
rect 21407 61013 21419 61047
rect 25406 61044 25412 61056
rect 25367 61016 25412 61044
rect 21361 61007 21419 61013
rect 25406 61004 25412 61016
rect 25464 61004 25470 61056
rect 27338 61044 27344 61056
rect 27299 61016 27344 61044
rect 27338 61004 27344 61016
rect 27396 61004 27402 61056
rect 28350 61044 28356 61056
rect 28311 61016 28356 61044
rect 28350 61004 28356 61016
rect 28408 61004 28414 61056
rect 29914 61044 29920 61056
rect 29875 61016 29920 61044
rect 29914 61004 29920 61016
rect 29972 61004 29978 61056
rect 31294 61044 31300 61056
rect 31255 61016 31300 61044
rect 31294 61004 31300 61016
rect 31352 61004 31358 61056
rect 32493 61047 32551 61053
rect 32493 61013 32505 61047
rect 32539 61044 32551 61047
rect 32582 61044 32588 61056
rect 32539 61016 32588 61044
rect 32539 61013 32551 61016
rect 32493 61007 32551 61013
rect 32582 61004 32588 61016
rect 32640 61004 32646 61056
rect 33410 61044 33416 61056
rect 33371 61016 33416 61044
rect 33410 61004 33416 61016
rect 33468 61004 33474 61056
rect 35066 61044 35072 61056
rect 35027 61016 35072 61044
rect 35066 61004 35072 61016
rect 35124 61004 35130 61056
rect 36078 61004 36084 61056
rect 36136 61044 36142 61056
rect 36541 61047 36599 61053
rect 36541 61044 36553 61047
rect 36136 61016 36553 61044
rect 36136 61004 36142 61016
rect 36541 61013 36553 61016
rect 36587 61013 36599 61047
rect 39114 61044 39120 61056
rect 39075 61016 39120 61044
rect 36541 61007 36599 61013
rect 39114 61004 39120 61016
rect 39172 61004 39178 61056
rect 40310 61004 40316 61056
rect 40368 61044 40374 61056
rect 40957 61047 41015 61053
rect 40957 61044 40969 61047
rect 40368 61016 40969 61044
rect 40368 61004 40374 61016
rect 40957 61013 40969 61016
rect 41003 61013 41015 61047
rect 41690 61044 41696 61056
rect 41651 61016 41696 61044
rect 40957 61007 41015 61013
rect 41690 61004 41696 61016
rect 41748 61004 41754 61056
rect 44450 61044 44456 61056
rect 44411 61016 44456 61044
rect 44450 61004 44456 61016
rect 44508 61004 44514 61056
rect 45370 61044 45376 61056
rect 45331 61016 45376 61044
rect 45370 61004 45376 61016
rect 45428 61004 45434 61056
rect 46106 61044 46112 61056
rect 46067 61016 46112 61044
rect 46106 61004 46112 61016
rect 46164 61004 46170 61056
rect 46842 61004 46848 61056
rect 46900 61044 46906 61056
rect 48685 61047 48743 61053
rect 48685 61044 48697 61047
rect 46900 61016 48697 61044
rect 46900 61004 46906 61016
rect 48685 61013 48697 61016
rect 48731 61013 48743 61047
rect 48685 61007 48743 61013
rect 50062 61004 50068 61056
rect 50120 61044 50126 61056
rect 50525 61047 50583 61053
rect 50525 61044 50537 61047
rect 50120 61016 50537 61044
rect 50120 61004 50126 61016
rect 50525 61013 50537 61016
rect 50571 61013 50583 61047
rect 50525 61007 50583 61013
rect 53190 61004 53196 61056
rect 53248 61004 53254 61056
rect 54294 61044 54300 61056
rect 54255 61016 54300 61044
rect 54294 61004 54300 61016
rect 54352 61004 54358 61056
rect 55186 61044 55214 61084
rect 55766 61072 55772 61084
rect 55824 61072 55830 61124
rect 56597 61047 56655 61053
rect 56597 61044 56609 61047
rect 55186 61016 56609 61044
rect 56597 61013 56609 61016
rect 56643 61013 56655 61047
rect 56597 61007 56655 61013
rect 56686 61004 56692 61056
rect 56744 61044 56750 61056
rect 58253 61047 58311 61053
rect 58253 61044 58265 61047
rect 56744 61016 58265 61044
rect 56744 61004 56750 61016
rect 58253 61013 58265 61016
rect 58299 61013 58311 61047
rect 58253 61007 58311 61013
rect 1104 60954 58880 60976
rect 1104 60902 19574 60954
rect 19626 60902 19638 60954
rect 19690 60902 19702 60954
rect 19754 60902 19766 60954
rect 19818 60902 19830 60954
rect 19882 60902 50294 60954
rect 50346 60902 50358 60954
rect 50410 60902 50422 60954
rect 50474 60902 50486 60954
rect 50538 60902 50550 60954
rect 50602 60902 58880 60954
rect 1104 60880 58880 60902
rect 5166 60800 5172 60852
rect 5224 60840 5230 60852
rect 23474 60840 23480 60852
rect 5224 60812 23480 60840
rect 5224 60800 5230 60812
rect 23474 60800 23480 60812
rect 23532 60800 23538 60852
rect 23750 60800 23756 60852
rect 23808 60840 23814 60852
rect 44450 60840 44456 60852
rect 23808 60812 44456 60840
rect 23808 60800 23814 60812
rect 44450 60800 44456 60812
rect 44508 60800 44514 60852
rect 3234 60772 3240 60784
rect 3195 60744 3240 60772
rect 3234 60732 3240 60744
rect 3292 60732 3298 60784
rect 3970 60772 3976 60784
rect 3931 60744 3976 60772
rect 3970 60732 3976 60744
rect 4028 60732 4034 60784
rect 8294 60732 8300 60784
rect 8352 60772 8358 60784
rect 8389 60775 8447 60781
rect 8389 60772 8401 60775
rect 8352 60744 8401 60772
rect 8352 60732 8358 60744
rect 8389 60741 8401 60744
rect 8435 60741 8447 60775
rect 13538 60772 13544 60784
rect 13499 60744 13544 60772
rect 8389 60735 8447 60741
rect 13538 60732 13544 60744
rect 13596 60732 13602 60784
rect 14274 60772 14280 60784
rect 14235 60744 14280 60772
rect 14274 60732 14280 60744
rect 14332 60732 14338 60784
rect 15746 60772 15752 60784
rect 15707 60744 15752 60772
rect 15746 60732 15752 60744
rect 15804 60732 15810 60784
rect 15838 60732 15844 60784
rect 15896 60772 15902 60784
rect 15896 60744 19288 60772
rect 15896 60732 15902 60744
rect 1578 60704 1584 60716
rect 1539 60676 1584 60704
rect 1578 60664 1584 60676
rect 1636 60664 1642 60716
rect 9030 60704 9036 60716
rect 8991 60676 9036 60704
rect 9030 60664 9036 60676
rect 9088 60664 9094 60716
rect 19260 60704 19288 60744
rect 19334 60732 19340 60784
rect 19392 60772 19398 60784
rect 19429 60775 19487 60781
rect 19429 60772 19441 60775
rect 19392 60744 19441 60772
rect 19392 60732 19398 60744
rect 19429 60741 19441 60744
rect 19475 60741 19487 60775
rect 23290 60772 23296 60784
rect 19429 60735 19487 60741
rect 21376 60744 23296 60772
rect 21376 60704 21404 60744
rect 23290 60732 23296 60744
rect 23348 60732 23354 60784
rect 24394 60732 24400 60784
rect 24452 60772 24458 60784
rect 24581 60775 24639 60781
rect 24581 60772 24593 60775
rect 24452 60744 24593 60772
rect 24452 60732 24458 60744
rect 24581 60741 24593 60744
rect 24627 60741 24639 60775
rect 27522 60772 27528 60784
rect 27483 60744 27528 60772
rect 24581 60735 24639 60741
rect 27522 60732 27528 60744
rect 27580 60732 27586 60784
rect 28810 60732 28816 60784
rect 28868 60772 28874 60784
rect 28997 60775 29055 60781
rect 28997 60772 29009 60775
rect 28868 60744 29009 60772
rect 28868 60732 28874 60744
rect 28997 60741 29009 60744
rect 29043 60741 29055 60775
rect 28997 60735 29055 60741
rect 30374 60732 30380 60784
rect 30432 60772 30438 60784
rect 30469 60775 30527 60781
rect 30469 60772 30481 60775
rect 30432 60744 30481 60772
rect 30432 60732 30438 60744
rect 30469 60741 30481 60744
rect 30515 60741 30527 60775
rect 36354 60772 36360 60784
rect 36315 60744 36360 60772
rect 30469 60735 30527 60741
rect 36354 60732 36360 60744
rect 36412 60732 36418 60784
rect 41414 60732 41420 60784
rect 41472 60772 41478 60784
rect 41509 60775 41567 60781
rect 41509 60772 41521 60775
rect 41472 60744 41521 60772
rect 41472 60732 41478 60744
rect 41509 60741 41521 60744
rect 41555 60741 41567 60775
rect 46658 60772 46664 60784
rect 46619 60744 46664 60772
rect 41509 60735 41567 60741
rect 46658 60732 46664 60744
rect 46716 60732 46722 60784
rect 50154 60732 50160 60784
rect 50212 60772 50218 60784
rect 50341 60775 50399 60781
rect 50341 60772 50353 60775
rect 50212 60744 50353 60772
rect 50212 60732 50218 60744
rect 50341 60741 50353 60744
rect 50387 60741 50399 60775
rect 50341 60735 50399 60741
rect 52454 60732 52460 60784
rect 52512 60772 52518 60784
rect 53009 60775 53067 60781
rect 53009 60772 53021 60775
rect 52512 60744 53021 60772
rect 52512 60732 52518 60744
rect 53009 60741 53021 60744
rect 53055 60741 53067 60775
rect 53009 60735 53067 60741
rect 19260 60676 21404 60704
rect 22094 60664 22100 60716
rect 22152 60704 22158 60716
rect 22554 60713 22560 60716
rect 22281 60707 22339 60713
rect 22152 60676 22197 60704
rect 22152 60664 22158 60676
rect 22281 60673 22293 60707
rect 22327 60673 22339 60707
rect 22281 60667 22339 60673
rect 22373 60707 22431 60713
rect 22373 60673 22385 60707
rect 22419 60673 22431 60707
rect 22373 60667 22431 60673
rect 22517 60707 22560 60713
rect 22517 60673 22529 60707
rect 22517 60667 22560 60673
rect 1857 60639 1915 60645
rect 1857 60605 1869 60639
rect 1903 60636 1915 60639
rect 5534 60636 5540 60648
rect 1903 60608 5540 60636
rect 1903 60605 1915 60608
rect 1857 60599 1915 60605
rect 5534 60596 5540 60608
rect 5592 60596 5598 60648
rect 4157 60571 4215 60577
rect 4157 60537 4169 60571
rect 4203 60568 4215 60571
rect 4614 60568 4620 60580
rect 4203 60540 4620 60568
rect 4203 60537 4215 60540
rect 4157 60531 4215 60537
rect 4614 60528 4620 60540
rect 4672 60528 4678 60580
rect 8573 60571 8631 60577
rect 8573 60537 8585 60571
rect 8619 60568 8631 60571
rect 18414 60568 18420 60580
rect 8619 60540 18420 60568
rect 8619 60537 8631 60540
rect 8573 60531 8631 60537
rect 18414 60528 18420 60540
rect 18472 60528 18478 60580
rect 19613 60571 19671 60577
rect 19613 60537 19625 60571
rect 19659 60568 19671 60571
rect 20622 60568 20628 60580
rect 19659 60540 20628 60568
rect 19659 60537 19671 60540
rect 19613 60531 19671 60537
rect 20622 60528 20628 60540
rect 20680 60528 20686 60580
rect 3326 60500 3332 60512
rect 3287 60472 3332 60500
rect 3326 60460 3332 60472
rect 3384 60460 3390 60512
rect 9214 60500 9220 60512
rect 9175 60472 9220 60500
rect 9214 60460 9220 60472
rect 9272 60460 9278 60512
rect 13630 60500 13636 60512
rect 13591 60472 13636 60500
rect 13630 60460 13636 60472
rect 13688 60460 13694 60512
rect 14366 60500 14372 60512
rect 14327 60472 14372 60500
rect 14366 60460 14372 60472
rect 14424 60460 14430 60512
rect 15841 60503 15899 60509
rect 15841 60469 15853 60503
rect 15887 60500 15899 60503
rect 17862 60500 17868 60512
rect 15887 60472 17868 60500
rect 15887 60469 15899 60472
rect 15841 60463 15899 60469
rect 17862 60460 17868 60472
rect 17920 60460 17926 60512
rect 20530 60460 20536 60512
rect 20588 60500 20594 60512
rect 22296 60500 22324 60667
rect 22388 60568 22416 60667
rect 22554 60664 22560 60667
rect 22612 60664 22618 60716
rect 23198 60704 23204 60716
rect 23159 60676 23204 60704
rect 23198 60664 23204 60676
rect 23256 60664 23262 60716
rect 54662 60704 54668 60716
rect 54623 60676 54668 60704
rect 54662 60664 54668 60676
rect 54720 60664 54726 60716
rect 55398 60704 55404 60716
rect 55359 60676 55404 60704
rect 55398 60664 55404 60676
rect 55456 60664 55462 60716
rect 56134 60704 56140 60716
rect 56095 60676 56140 60704
rect 56134 60664 56140 60676
rect 56192 60664 56198 60716
rect 56870 60704 56876 60716
rect 56831 60676 56876 60704
rect 56870 60664 56876 60676
rect 56928 60664 56934 60716
rect 58066 60704 58072 60716
rect 58027 60676 58072 60704
rect 58066 60664 58072 60676
rect 58124 60664 58130 60716
rect 22572 60636 22600 60664
rect 40770 60636 40776 60648
rect 22572 60608 40776 60636
rect 40770 60596 40776 60608
rect 40828 60596 40834 60648
rect 56321 60571 56379 60577
rect 56321 60568 56333 60571
rect 22388 60540 56333 60568
rect 56321 60537 56333 60540
rect 56367 60537 56379 60571
rect 56321 60531 56379 60537
rect 22462 60500 22468 60512
rect 20588 60472 22468 60500
rect 20588 60460 20594 60472
rect 22462 60460 22468 60472
rect 22520 60460 22526 60512
rect 22649 60503 22707 60509
rect 22649 60469 22661 60503
rect 22695 60500 22707 60503
rect 22922 60500 22928 60512
rect 22695 60472 22928 60500
rect 22695 60469 22707 60472
rect 22649 60463 22707 60469
rect 22922 60460 22928 60472
rect 22980 60460 22986 60512
rect 23382 60500 23388 60512
rect 23343 60472 23388 60500
rect 23382 60460 23388 60472
rect 23440 60460 23446 60512
rect 24673 60503 24731 60509
rect 24673 60469 24685 60503
rect 24719 60500 24731 60503
rect 25222 60500 25228 60512
rect 24719 60472 25228 60500
rect 24719 60469 24731 60472
rect 24673 60463 24731 60469
rect 25222 60460 25228 60472
rect 25280 60460 25286 60512
rect 27617 60503 27675 60509
rect 27617 60469 27629 60503
rect 27663 60500 27675 60503
rect 28994 60500 29000 60512
rect 27663 60472 29000 60500
rect 27663 60469 27675 60472
rect 27617 60463 27675 60469
rect 28994 60460 29000 60472
rect 29052 60460 29058 60512
rect 29089 60503 29147 60509
rect 29089 60469 29101 60503
rect 29135 60500 29147 60503
rect 29822 60500 29828 60512
rect 29135 60472 29828 60500
rect 29135 60469 29147 60472
rect 29089 60463 29147 60469
rect 29822 60460 29828 60472
rect 29880 60460 29886 60512
rect 30558 60500 30564 60512
rect 30519 60472 30564 60500
rect 30558 60460 30564 60472
rect 30616 60460 30622 60512
rect 33042 60460 33048 60512
rect 33100 60500 33106 60512
rect 35066 60500 35072 60512
rect 33100 60472 35072 60500
rect 33100 60460 33106 60472
rect 35066 60460 35072 60472
rect 35124 60460 35130 60512
rect 35710 60460 35716 60512
rect 35768 60500 35774 60512
rect 36449 60503 36507 60509
rect 36449 60500 36461 60503
rect 35768 60472 36461 60500
rect 35768 60460 35774 60472
rect 36449 60469 36461 60472
rect 36495 60469 36507 60503
rect 36449 60463 36507 60469
rect 40862 60460 40868 60512
rect 40920 60500 40926 60512
rect 41601 60503 41659 60509
rect 41601 60500 41613 60503
rect 40920 60472 41613 60500
rect 40920 60460 40926 60472
rect 41601 60469 41613 60472
rect 41647 60469 41659 60503
rect 41601 60463 41659 60469
rect 44174 60460 44180 60512
rect 44232 60500 44238 60512
rect 46753 60503 46811 60509
rect 46753 60500 46765 60503
rect 44232 60472 46765 60500
rect 44232 60460 44238 60472
rect 46753 60469 46765 60472
rect 46799 60469 46811 60503
rect 50430 60500 50436 60512
rect 50391 60472 50436 60500
rect 46753 60463 46811 60469
rect 50430 60460 50436 60472
rect 50488 60460 50494 60512
rect 53098 60500 53104 60512
rect 53059 60472 53104 60500
rect 53098 60460 53104 60472
rect 53156 60460 53162 60512
rect 54846 60500 54852 60512
rect 54807 60472 54852 60500
rect 54846 60460 54852 60472
rect 54904 60460 54910 60512
rect 55582 60500 55588 60512
rect 55543 60472 55588 60500
rect 55582 60460 55588 60472
rect 55640 60460 55646 60512
rect 57054 60500 57060 60512
rect 57015 60472 57060 60500
rect 57054 60460 57060 60472
rect 57112 60460 57118 60512
rect 58250 60500 58256 60512
rect 58211 60472 58256 60500
rect 58250 60460 58256 60472
rect 58308 60460 58314 60512
rect 1104 60410 58880 60432
rect 1104 60358 4214 60410
rect 4266 60358 4278 60410
rect 4330 60358 4342 60410
rect 4394 60358 4406 60410
rect 4458 60358 4470 60410
rect 4522 60358 34934 60410
rect 34986 60358 34998 60410
rect 35050 60358 35062 60410
rect 35114 60358 35126 60410
rect 35178 60358 35190 60410
rect 35242 60358 58880 60410
rect 1104 60336 58880 60358
rect 3326 60256 3332 60308
rect 3384 60296 3390 60308
rect 20254 60296 20260 60308
rect 3384 60268 20260 60296
rect 3384 60256 3390 60268
rect 20254 60256 20260 60268
rect 20312 60256 20318 60308
rect 20714 60256 20720 60308
rect 20772 60296 20778 60308
rect 55582 60296 55588 60308
rect 20772 60268 55588 60296
rect 20772 60256 20778 60268
rect 55582 60256 55588 60268
rect 55640 60256 55646 60308
rect 13630 60188 13636 60240
rect 13688 60228 13694 60240
rect 20993 60231 21051 60237
rect 13688 60200 20668 60228
rect 13688 60188 13694 60200
rect 17862 60160 17868 60172
rect 7760 60132 17724 60160
rect 17823 60132 17868 60160
rect 2590 60092 2596 60104
rect 2551 60064 2596 60092
rect 2590 60052 2596 60064
rect 2648 60052 2654 60104
rect 5626 60052 5632 60104
rect 5684 60092 5690 60104
rect 7377 60095 7435 60101
rect 7377 60092 7389 60095
rect 5684 60064 7389 60092
rect 5684 60052 5690 60064
rect 7377 60061 7389 60064
rect 7423 60061 7435 60095
rect 7650 60092 7656 60104
rect 7611 60064 7656 60092
rect 7377 60055 7435 60061
rect 7650 60052 7656 60064
rect 7708 60052 7714 60104
rect 7760 60101 7788 60132
rect 7745 60095 7803 60101
rect 7745 60061 7757 60095
rect 7791 60061 7803 60095
rect 7745 60055 7803 60061
rect 1670 60024 1676 60036
rect 1631 59996 1676 60024
rect 1670 59984 1676 59996
rect 1728 59984 1734 60036
rect 2038 60024 2044 60036
rect 1999 59996 2044 60024
rect 2038 59984 2044 59996
rect 2096 59984 2102 60036
rect 7561 60027 7619 60033
rect 7561 59993 7573 60027
rect 7607 59993 7619 60027
rect 17586 60024 17592 60036
rect 7561 59987 7619 59993
rect 7852 59996 17592 60024
rect 2498 59916 2504 59968
rect 2556 59956 2562 59968
rect 2685 59959 2743 59965
rect 2685 59956 2697 59959
rect 2556 59928 2697 59956
rect 2556 59916 2562 59928
rect 2685 59925 2697 59928
rect 2731 59925 2743 59959
rect 7576 59956 7604 59987
rect 7852 59956 7880 59996
rect 17586 59984 17592 59996
rect 17644 59984 17650 60036
rect 7576 59928 7880 59956
rect 7929 59959 7987 59965
rect 2685 59919 2743 59925
rect 7929 59925 7941 59959
rect 7975 59956 7987 59959
rect 8018 59956 8024 59968
rect 7975 59928 8024 59956
rect 7975 59925 7987 59928
rect 7929 59919 7987 59925
rect 8018 59916 8024 59928
rect 8076 59916 8082 59968
rect 17494 59956 17500 59968
rect 17455 59928 17500 59956
rect 17494 59916 17500 59928
rect 17552 59916 17558 59968
rect 17696 59956 17724 60132
rect 17862 60120 17868 60132
rect 17920 60120 17926 60172
rect 20640 60160 20668 60200
rect 20993 60197 21005 60231
rect 21039 60228 21051 60231
rect 21358 60228 21364 60240
rect 21039 60200 21364 60228
rect 21039 60197 21051 60200
rect 20993 60191 21051 60197
rect 21358 60188 21364 60200
rect 21416 60188 21422 60240
rect 22646 60188 22652 60240
rect 22704 60228 22710 60240
rect 23382 60228 23388 60240
rect 22704 60200 23388 60228
rect 22704 60188 22710 60200
rect 23382 60188 23388 60200
rect 23440 60188 23446 60240
rect 30190 60228 30196 60240
rect 28552 60200 30196 60228
rect 26878 60160 26884 60172
rect 18064 60132 20576 60160
rect 20640 60132 26884 60160
rect 18064 60101 18092 60132
rect 20548 60104 20576 60132
rect 26878 60120 26884 60132
rect 26936 60120 26942 60172
rect 28552 60160 28580 60200
rect 30190 60188 30196 60200
rect 30248 60228 30254 60240
rect 41138 60228 41144 60240
rect 30248 60200 30788 60228
rect 41099 60200 41144 60228
rect 30248 60188 30254 60200
rect 27724 60132 28580 60160
rect 18049 60095 18107 60101
rect 18049 60061 18061 60095
rect 18095 60061 18107 60095
rect 18414 60092 18420 60104
rect 18375 60064 18420 60092
rect 18049 60055 18107 60061
rect 18414 60052 18420 60064
rect 18472 60052 18478 60104
rect 18598 60092 18604 60104
rect 18559 60064 18604 60092
rect 18598 60052 18604 60064
rect 18656 60052 18662 60104
rect 19978 60092 19984 60104
rect 18708 60064 19984 60092
rect 18708 59956 18736 60064
rect 19978 60052 19984 60064
rect 20036 60052 20042 60104
rect 20438 60092 20444 60104
rect 20399 60064 20444 60092
rect 20438 60052 20444 60064
rect 20496 60052 20502 60104
rect 20530 60052 20536 60104
rect 20588 60092 20594 60104
rect 20625 60095 20683 60101
rect 20625 60092 20637 60095
rect 20588 60064 20637 60092
rect 20588 60052 20594 60064
rect 20625 60061 20637 60064
rect 20671 60061 20683 60095
rect 20625 60055 20683 60061
rect 20714 60052 20720 60104
rect 20772 60092 20778 60104
rect 20861 60095 20919 60101
rect 20772 60064 20817 60092
rect 20772 60052 20778 60064
rect 20861 60061 20873 60095
rect 20907 60092 20919 60095
rect 21818 60092 21824 60104
rect 20907 60064 21824 60092
rect 20907 60061 20919 60064
rect 20861 60055 20919 60061
rect 21818 60052 21824 60064
rect 21876 60052 21882 60104
rect 22002 60092 22008 60104
rect 21963 60064 22008 60092
rect 22002 60052 22008 60064
rect 22060 60052 22066 60104
rect 22094 60052 22100 60104
rect 22152 60092 22158 60104
rect 22370 60092 22376 60104
rect 22152 60064 22197 60092
rect 22331 60064 22376 60092
rect 22152 60052 22158 60064
rect 22370 60052 22376 60064
rect 22428 60052 22434 60104
rect 22462 60052 22468 60104
rect 22520 60092 22526 60104
rect 22649 60095 22707 60101
rect 22649 60092 22661 60095
rect 22520 60064 22661 60092
rect 22520 60052 22526 60064
rect 22649 60061 22661 60064
rect 22695 60061 22707 60095
rect 22830 60092 22836 60104
rect 22791 60064 22836 60092
rect 22649 60055 22707 60061
rect 19242 59984 19248 60036
rect 19300 60024 19306 60036
rect 21266 60024 21272 60036
rect 19300 59996 21272 60024
rect 19300 59984 19306 59996
rect 21266 59984 21272 59996
rect 21324 60024 21330 60036
rect 22664 60024 22692 60055
rect 22830 60052 22836 60064
rect 22888 60052 22894 60104
rect 23474 60092 23480 60104
rect 23435 60064 23480 60092
rect 23474 60052 23480 60064
rect 23532 60052 23538 60104
rect 23750 60092 23756 60104
rect 23711 60064 23756 60092
rect 23750 60052 23756 60064
rect 23808 60052 23814 60104
rect 23845 60095 23903 60101
rect 23845 60061 23857 60095
rect 23891 60092 23903 60095
rect 23934 60092 23940 60104
rect 23891 60064 23940 60092
rect 23891 60061 23903 60064
rect 23845 60055 23903 60061
rect 23934 60052 23940 60064
rect 23992 60092 23998 60104
rect 27724 60092 27752 60132
rect 28074 60092 28080 60104
rect 23992 60064 27752 60092
rect 28035 60064 28080 60092
rect 23992 60052 23998 60064
rect 28074 60052 28080 60064
rect 28132 60052 28138 60104
rect 28166 60052 28172 60104
rect 28224 60092 28230 60104
rect 28442 60092 28448 60104
rect 28224 60064 28269 60092
rect 28403 60064 28448 60092
rect 28224 60052 28230 60064
rect 28442 60052 28448 60064
rect 28500 60052 28506 60104
rect 28552 60101 28580 60132
rect 28994 60120 29000 60172
rect 29052 60160 29058 60172
rect 29052 60132 30512 60160
rect 29052 60120 29058 60132
rect 28542 60095 28600 60101
rect 28542 60061 28554 60095
rect 28588 60061 28600 60095
rect 28542 60055 28600 60061
rect 30101 60095 30159 60101
rect 30101 60061 30113 60095
rect 30147 60092 30159 60095
rect 30374 60092 30380 60104
rect 30147 60064 30380 60092
rect 30147 60061 30159 60064
rect 30101 60055 30159 60061
rect 30374 60052 30380 60064
rect 30432 60052 30438 60104
rect 30484 60101 30512 60132
rect 30470 60095 30528 60101
rect 30470 60061 30482 60095
rect 30516 60061 30528 60095
rect 30760 60092 30788 60200
rect 41138 60188 41144 60200
rect 41196 60188 41202 60240
rect 50430 60228 50436 60240
rect 42720 60200 50436 60228
rect 41506 60160 41512 60172
rect 31588 60132 33272 60160
rect 30883 60095 30941 60101
rect 30883 60092 30895 60095
rect 30760 60064 30895 60092
rect 30470 60055 30528 60061
rect 30883 60061 30895 60064
rect 30929 60092 30941 60095
rect 31588 60092 31616 60132
rect 32490 60092 32496 60104
rect 30929 60064 31616 60092
rect 32451 60064 32496 60092
rect 30929 60061 30941 60064
rect 30883 60055 30941 60061
rect 32490 60052 32496 60064
rect 32548 60052 32554 60104
rect 32674 60092 32680 60104
rect 32635 60064 32680 60092
rect 32674 60052 32680 60064
rect 32732 60052 32738 60104
rect 33042 60052 33048 60104
rect 33100 60092 33106 60104
rect 33244 60101 33272 60132
rect 35866 60132 41512 60160
rect 33229 60095 33287 60101
rect 33100 60064 33145 60092
rect 33100 60052 33106 60064
rect 33229 60061 33241 60095
rect 33275 60092 33287 60095
rect 34514 60092 34520 60104
rect 33275 60064 34520 60092
rect 33275 60061 33287 60064
rect 33229 60055 33287 60061
rect 34514 60052 34520 60064
rect 34572 60052 34578 60104
rect 23566 60024 23572 60036
rect 21324 59996 21864 60024
rect 22664 59996 23572 60024
rect 21324 59984 21330 59996
rect 21634 59956 21640 59968
rect 17696 59928 18736 59956
rect 21595 59928 21640 59956
rect 21634 59916 21640 59928
rect 21692 59916 21698 59968
rect 21836 59956 21864 59996
rect 23566 59984 23572 59996
rect 23624 59984 23630 60036
rect 23661 60027 23719 60033
rect 23661 59993 23673 60027
rect 23707 59993 23719 60027
rect 23661 59987 23719 59993
rect 28353 60027 28411 60033
rect 28353 59993 28365 60027
rect 28399 60024 28411 60027
rect 30006 60024 30012 60036
rect 28399 59996 30012 60024
rect 28399 59993 28411 59996
rect 28353 59987 28411 59993
rect 23676 59956 23704 59987
rect 28552 59968 28580 59996
rect 30006 59984 30012 59996
rect 30064 60024 30070 60036
rect 30650 60024 30656 60036
rect 30064 59996 30656 60024
rect 30064 59984 30070 59996
rect 30650 59984 30656 59996
rect 30708 59984 30714 60036
rect 30745 60027 30803 60033
rect 30745 59993 30757 60027
rect 30791 60024 30803 60027
rect 35866 60024 35894 60132
rect 41506 60120 41512 60132
rect 41564 60120 41570 60172
rect 42613 60163 42671 60169
rect 42613 60160 42625 60163
rect 41616 60132 42625 60160
rect 40586 60092 40592 60104
rect 40547 60064 40592 60092
rect 40586 60052 40592 60064
rect 40644 60052 40650 60104
rect 40862 60092 40868 60104
rect 40823 60064 40868 60092
rect 40862 60052 40868 60064
rect 40920 60052 40926 60104
rect 40954 60052 40960 60104
rect 41012 60101 41018 60104
rect 41012 60092 41020 60101
rect 41616 60092 41644 60132
rect 42613 60129 42625 60132
rect 42659 60129 42671 60163
rect 42613 60123 42671 60129
rect 42150 60092 42156 60104
rect 41012 60064 41644 60092
rect 42111 60064 42156 60092
rect 41012 60055 41020 60064
rect 41012 60052 41018 60055
rect 42150 60052 42156 60064
rect 42208 60052 42214 60104
rect 42334 60092 42340 60104
rect 42295 60064 42340 60092
rect 42334 60052 42340 60064
rect 42392 60052 42398 60104
rect 40770 60024 40776 60036
rect 30791 59996 35894 60024
rect 40731 59996 40776 60024
rect 30791 59993 30803 59996
rect 30745 59987 30803 59993
rect 40770 59984 40776 59996
rect 40828 59984 40834 60036
rect 42628 60024 42656 60123
rect 42720 60101 42748 60200
rect 50430 60188 50436 60200
rect 50488 60188 50494 60240
rect 53926 60120 53932 60172
rect 53984 60160 53990 60172
rect 57425 60163 57483 60169
rect 57425 60160 57437 60163
rect 53984 60132 57437 60160
rect 53984 60120 53990 60132
rect 57425 60129 57437 60132
rect 57471 60129 57483 60163
rect 57425 60123 57483 60129
rect 42705 60095 42763 60101
rect 42705 60061 42717 60095
rect 42751 60061 42763 60095
rect 56502 60092 56508 60104
rect 56463 60064 56508 60092
rect 42705 60055 42763 60061
rect 56502 60052 56508 60064
rect 56560 60052 56566 60104
rect 57238 60092 57244 60104
rect 57199 60064 57244 60092
rect 57238 60052 57244 60064
rect 57296 60052 57302 60104
rect 57885 60095 57943 60101
rect 57885 60061 57897 60095
rect 57931 60092 57943 60095
rect 57974 60092 57980 60104
rect 57931 60064 57980 60092
rect 57931 60061 57943 60064
rect 57885 60055 57943 60061
rect 57974 60052 57980 60064
rect 58032 60052 58038 60104
rect 43530 60024 43536 60036
rect 42628 59996 43536 60024
rect 43530 59984 43536 59996
rect 43588 59984 43594 60036
rect 58161 60027 58219 60033
rect 58161 59993 58173 60027
rect 58207 60024 58219 60027
rect 58250 60024 58256 60036
rect 58207 59996 58256 60024
rect 58207 59993 58219 59996
rect 58161 59987 58219 59993
rect 58250 59984 58256 59996
rect 58308 59984 58314 60036
rect 21836 59928 23704 59956
rect 24029 59959 24087 59965
rect 24029 59925 24041 59959
rect 24075 59956 24087 59959
rect 24394 59956 24400 59968
rect 24075 59928 24400 59956
rect 24075 59925 24087 59928
rect 24029 59919 24087 59925
rect 24394 59916 24400 59928
rect 24452 59916 24458 59968
rect 28534 59916 28540 59968
rect 28592 59916 28598 59968
rect 28718 59956 28724 59968
rect 28679 59928 28724 59956
rect 28718 59916 28724 59928
rect 28776 59916 28782 59968
rect 31018 59956 31024 59968
rect 30979 59928 31024 59956
rect 31018 59916 31024 59928
rect 31076 59916 31082 59968
rect 32306 59956 32312 59968
rect 32267 59928 32312 59956
rect 32306 59916 32312 59928
rect 32364 59916 32370 59968
rect 41966 59956 41972 59968
rect 41927 59928 41972 59956
rect 41966 59916 41972 59928
rect 42024 59916 42030 59968
rect 54110 59916 54116 59968
rect 54168 59956 54174 59968
rect 56597 59959 56655 59965
rect 56597 59956 56609 59959
rect 54168 59928 56609 59956
rect 54168 59916 54174 59928
rect 56597 59925 56609 59928
rect 56643 59925 56655 59959
rect 56597 59919 56655 59925
rect 1104 59866 58880 59888
rect 1104 59814 19574 59866
rect 19626 59814 19638 59866
rect 19690 59814 19702 59866
rect 19754 59814 19766 59866
rect 19818 59814 19830 59866
rect 19882 59814 50294 59866
rect 50346 59814 50358 59866
rect 50410 59814 50422 59866
rect 50474 59814 50486 59866
rect 50538 59814 50550 59866
rect 50602 59814 58880 59866
rect 1104 59792 58880 59814
rect 14366 59712 14372 59764
rect 14424 59752 14430 59764
rect 32490 59752 32496 59764
rect 14424 59724 32496 59752
rect 14424 59712 14430 59724
rect 32490 59712 32496 59724
rect 32548 59712 32554 59764
rect 32674 59712 32680 59764
rect 32732 59752 32738 59764
rect 33042 59752 33048 59764
rect 32732 59724 33048 59752
rect 32732 59712 32738 59724
rect 33042 59712 33048 59724
rect 33100 59752 33106 59764
rect 42334 59752 42340 59764
rect 33100 59724 42340 59752
rect 33100 59712 33106 59724
rect 42334 59712 42340 59724
rect 42392 59712 42398 59764
rect 58253 59755 58311 59761
rect 58253 59752 58265 59755
rect 45526 59724 58265 59752
rect 1762 59644 1768 59696
rect 1820 59684 1826 59696
rect 2593 59687 2651 59693
rect 2593 59684 2605 59687
rect 1820 59656 2605 59684
rect 1820 59644 1826 59656
rect 2593 59653 2605 59656
rect 2639 59653 2651 59687
rect 2593 59647 2651 59653
rect 18230 59644 18236 59696
rect 18288 59684 18294 59696
rect 20993 59687 21051 59693
rect 18288 59656 20852 59684
rect 18288 59644 18294 59656
rect 1670 59616 1676 59628
rect 1631 59588 1676 59616
rect 1670 59576 1676 59588
rect 1728 59576 1734 59628
rect 17954 59576 17960 59628
rect 18012 59616 18018 59628
rect 19337 59619 19395 59625
rect 19337 59616 19349 59619
rect 18012 59588 19349 59616
rect 18012 59576 18018 59588
rect 19337 59585 19349 59588
rect 19383 59585 19395 59619
rect 19337 59579 19395 59585
rect 19521 59619 19579 59625
rect 19521 59585 19533 59619
rect 19567 59585 19579 59619
rect 19521 59579 19579 59585
rect 19613 59619 19671 59625
rect 19613 59585 19625 59619
rect 19659 59585 19671 59619
rect 19613 59579 19671 59585
rect 19757 59619 19815 59625
rect 19757 59585 19769 59619
rect 19803 59616 19815 59619
rect 19978 59616 19984 59628
rect 19803 59588 19984 59616
rect 19803 59585 19815 59588
rect 19757 59579 19815 59585
rect 17586 59508 17592 59560
rect 17644 59548 17650 59560
rect 19242 59548 19248 59560
rect 17644 59520 19248 59548
rect 17644 59508 17650 59520
rect 19242 59508 19248 59520
rect 19300 59548 19306 59560
rect 19536 59548 19564 59579
rect 19300 59520 19564 59548
rect 19300 59508 19306 59520
rect 1946 59412 1952 59424
rect 1907 59384 1952 59412
rect 1946 59372 1952 59384
rect 2004 59372 2010 59424
rect 2314 59372 2320 59424
rect 2372 59412 2378 59424
rect 2685 59415 2743 59421
rect 2685 59412 2697 59415
rect 2372 59384 2697 59412
rect 2372 59372 2378 59384
rect 2685 59381 2697 59384
rect 2731 59381 2743 59415
rect 19628 59412 19656 59579
rect 19978 59576 19984 59588
rect 20036 59616 20042 59628
rect 20824 59625 20852 59656
rect 20993 59653 21005 59687
rect 21039 59684 21051 59687
rect 21450 59684 21456 59696
rect 21039 59656 21456 59684
rect 21039 59653 21051 59656
rect 20993 59647 21051 59653
rect 21450 59644 21456 59656
rect 21508 59644 21514 59696
rect 23382 59684 23388 59696
rect 21560 59656 23152 59684
rect 23343 59656 23388 59684
rect 20809 59619 20867 59625
rect 20036 59588 20668 59616
rect 20036 59576 20042 59588
rect 20640 59548 20668 59588
rect 20809 59585 20821 59619
rect 20855 59585 20867 59619
rect 21082 59616 21088 59628
rect 21043 59588 21088 59616
rect 20809 59579 20867 59585
rect 21082 59576 21088 59588
rect 21140 59576 21146 59628
rect 21177 59619 21235 59625
rect 21177 59585 21189 59619
rect 21223 59616 21235 59619
rect 21560 59616 21588 59656
rect 21223 59588 21588 59616
rect 21223 59585 21235 59588
rect 21177 59579 21235 59585
rect 21284 59548 21312 59588
rect 22094 59576 22100 59628
rect 22152 59616 22158 59628
rect 22649 59619 22707 59625
rect 22152 59588 22197 59616
rect 22152 59576 22158 59588
rect 22649 59585 22661 59619
rect 22695 59616 22707 59619
rect 22738 59616 22744 59628
rect 22695 59588 22744 59616
rect 22695 59585 22707 59588
rect 22649 59579 22707 59585
rect 22738 59576 22744 59588
rect 22796 59576 22802 59628
rect 20640 59520 21312 59548
rect 21361 59483 21419 59489
rect 19812 59452 20392 59480
rect 19812 59412 19840 59452
rect 19628 59384 19840 59412
rect 19889 59415 19947 59421
rect 2685 59375 2743 59381
rect 19889 59381 19901 59415
rect 19935 59412 19947 59415
rect 20162 59412 20168 59424
rect 19935 59384 20168 59412
rect 19935 59381 19947 59384
rect 19889 59375 19947 59381
rect 20162 59372 20168 59384
rect 20220 59372 20226 59424
rect 20364 59412 20392 59452
rect 21361 59449 21373 59483
rect 21407 59480 21419 59483
rect 22370 59480 22376 59492
rect 21407 59452 22376 59480
rect 21407 59449 21419 59452
rect 21361 59443 21419 59449
rect 22370 59440 22376 59452
rect 22428 59440 22434 59492
rect 23124 59480 23152 59656
rect 23382 59644 23388 59656
rect 23440 59644 23446 59696
rect 30098 59684 30104 59696
rect 30059 59656 30104 59684
rect 30098 59644 30104 59656
rect 30156 59644 30162 59696
rect 45526 59684 45554 59724
rect 58253 59721 58265 59724
rect 58299 59721 58311 59755
rect 58253 59715 58311 59721
rect 30392 59656 45554 59684
rect 23201 59619 23259 59625
rect 23201 59585 23213 59619
rect 23247 59585 23259 59619
rect 23201 59579 23259 59585
rect 23216 59548 23244 59579
rect 23290 59576 23296 59628
rect 23348 59616 23354 59628
rect 23658 59625 23664 59628
rect 23477 59619 23535 59625
rect 23477 59616 23489 59619
rect 23348 59588 23489 59616
rect 23348 59576 23354 59588
rect 23477 59585 23489 59588
rect 23523 59585 23535 59619
rect 23477 59579 23535 59585
rect 23621 59619 23664 59625
rect 23621 59585 23633 59619
rect 23621 59579 23664 59585
rect 23658 59576 23664 59579
rect 23716 59576 23722 59628
rect 28353 59619 28411 59625
rect 28353 59585 28365 59619
rect 28399 59616 28411 59619
rect 28442 59616 28448 59628
rect 28399 59588 28448 59616
rect 28399 59585 28411 59588
rect 28353 59579 28411 59585
rect 28442 59576 28448 59588
rect 28500 59576 28506 59628
rect 29730 59616 29736 59628
rect 29691 59588 29736 59616
rect 29730 59576 29736 59588
rect 29788 59576 29794 59628
rect 29822 59576 29828 59628
rect 29880 59616 29886 59628
rect 29880 59588 29925 59616
rect 29880 59576 29886 59588
rect 30006 59576 30012 59628
rect 30064 59616 30070 59628
rect 30064 59588 30109 59616
rect 30064 59576 30070 59588
rect 30190 59576 30196 59628
rect 30248 59625 30254 59628
rect 30248 59616 30256 59625
rect 30248 59588 30293 59616
rect 30248 59579 30256 59588
rect 30248 59576 30254 59579
rect 28534 59548 28540 59560
rect 23216 59520 23612 59548
rect 28495 59520 28540 59548
rect 23474 59480 23480 59492
rect 23124 59452 23480 59480
rect 23474 59440 23480 59452
rect 23532 59440 23538 59492
rect 23584 59480 23612 59520
rect 28534 59508 28540 59520
rect 28592 59508 28598 59560
rect 28626 59508 28632 59560
rect 28684 59548 28690 59560
rect 30098 59548 30104 59560
rect 28684 59520 30104 59548
rect 28684 59508 28690 59520
rect 30098 59508 30104 59520
rect 30156 59508 30162 59560
rect 30392 59548 30420 59656
rect 56410 59644 56416 59696
rect 56468 59684 56474 59696
rect 57333 59687 57391 59693
rect 57333 59684 57345 59687
rect 56468 59656 57345 59684
rect 56468 59644 56474 59656
rect 57333 59653 57345 59656
rect 57379 59653 57391 59687
rect 57333 59647 57391 59653
rect 30558 59576 30564 59628
rect 30616 59616 30622 59628
rect 42150 59616 42156 59628
rect 30616 59588 42156 59616
rect 30616 59576 30622 59588
rect 42150 59576 42156 59588
rect 42208 59576 42214 59628
rect 42334 59576 42340 59628
rect 42392 59616 42398 59628
rect 43257 59619 43315 59625
rect 43257 59616 43269 59619
rect 42392 59588 43269 59616
rect 42392 59576 42398 59588
rect 43257 59585 43269 59588
rect 43303 59585 43315 59619
rect 43257 59579 43315 59585
rect 43625 59619 43683 59625
rect 43625 59585 43637 59619
rect 43671 59616 43683 59619
rect 53098 59616 53104 59628
rect 43671 59588 53104 59616
rect 43671 59585 43683 59588
rect 43625 59579 43683 59585
rect 53098 59576 53104 59588
rect 53156 59576 53162 59628
rect 58066 59616 58072 59628
rect 58027 59588 58072 59616
rect 58066 59576 58072 59588
rect 58124 59576 58130 59628
rect 30650 59548 30656 59560
rect 30300 59520 30420 59548
rect 30484 59520 30656 59548
rect 30300 59480 30328 59520
rect 30484 59480 30512 59520
rect 30650 59508 30656 59520
rect 30708 59508 30714 59560
rect 42702 59548 42708 59560
rect 42663 59520 42708 59548
rect 42702 59508 42708 59520
rect 42760 59508 42766 59560
rect 42794 59508 42800 59560
rect 42852 59548 42858 59560
rect 43073 59551 43131 59557
rect 43073 59548 43085 59551
rect 42852 59520 43085 59548
rect 42852 59508 42858 59520
rect 43073 59517 43085 59520
rect 43119 59517 43131 59551
rect 43530 59548 43536 59560
rect 43491 59520 43536 59548
rect 43073 59511 43131 59517
rect 43530 59508 43536 59520
rect 43588 59508 43594 59560
rect 23584 59452 30328 59480
rect 30392 59452 30512 59480
rect 21174 59412 21180 59424
rect 20364 59384 21180 59412
rect 21174 59372 21180 59384
rect 21232 59372 21238 59424
rect 21450 59372 21456 59424
rect 21508 59412 21514 59424
rect 23658 59412 23664 59424
rect 21508 59384 23664 59412
rect 21508 59372 21514 59384
rect 23658 59372 23664 59384
rect 23716 59372 23722 59424
rect 23753 59415 23811 59421
rect 23753 59381 23765 59415
rect 23799 59412 23811 59415
rect 24486 59412 24492 59424
rect 23799 59384 24492 59412
rect 23799 59381 23811 59384
rect 23753 59375 23811 59381
rect 24486 59372 24492 59384
rect 24544 59372 24550 59424
rect 29457 59415 29515 59421
rect 29457 59381 29469 59415
rect 29503 59412 29515 59415
rect 29730 59412 29736 59424
rect 29503 59384 29736 59412
rect 29503 59381 29515 59384
rect 29457 59375 29515 59381
rect 29730 59372 29736 59384
rect 29788 59412 29794 59424
rect 30282 59412 30288 59424
rect 29788 59384 30288 59412
rect 29788 59372 29794 59384
rect 30282 59372 30288 59384
rect 30340 59372 30346 59424
rect 30392 59421 30420 59452
rect 30558 59440 30564 59492
rect 30616 59480 30622 59492
rect 32950 59480 32956 59492
rect 30616 59452 32956 59480
rect 30616 59440 30622 59452
rect 32950 59440 32956 59452
rect 33008 59440 33014 59492
rect 40586 59440 40592 59492
rect 40644 59480 40650 59492
rect 57517 59483 57575 59489
rect 57517 59480 57529 59483
rect 40644 59452 57529 59480
rect 40644 59440 40650 59452
rect 57517 59449 57529 59452
rect 57563 59449 57575 59483
rect 57517 59443 57575 59449
rect 30377 59415 30435 59421
rect 30377 59381 30389 59415
rect 30423 59381 30435 59415
rect 30377 59375 30435 59381
rect 30466 59372 30472 59424
rect 30524 59412 30530 59424
rect 30745 59415 30803 59421
rect 30745 59412 30757 59415
rect 30524 59384 30757 59412
rect 30524 59372 30530 59384
rect 30745 59381 30757 59384
rect 30791 59412 30803 59415
rect 31570 59412 31576 59424
rect 30791 59384 31576 59412
rect 30791 59381 30803 59384
rect 30745 59375 30803 59381
rect 31570 59372 31576 59384
rect 31628 59372 31634 59424
rect 57146 59372 57152 59424
rect 57204 59412 57210 59424
rect 58986 59412 58992 59424
rect 57204 59384 58992 59412
rect 57204 59372 57210 59384
rect 58986 59372 58992 59384
rect 59044 59372 59050 59424
rect 1104 59322 58880 59344
rect 1104 59270 4214 59322
rect 4266 59270 4278 59322
rect 4330 59270 4342 59322
rect 4394 59270 4406 59322
rect 4458 59270 4470 59322
rect 4522 59270 34934 59322
rect 34986 59270 34998 59322
rect 35050 59270 35062 59322
rect 35114 59270 35126 59322
rect 35178 59270 35190 59322
rect 35242 59270 58880 59322
rect 1104 59248 58880 59270
rect 57333 59211 57391 59217
rect 57333 59208 57345 59211
rect 19444 59180 57345 59208
rect 1946 59032 1952 59084
rect 2004 59072 2010 59084
rect 2004 59044 6914 59072
rect 2004 59032 2010 59044
rect 842 58964 848 59016
rect 900 59004 906 59016
rect 1673 59007 1731 59013
rect 1673 59004 1685 59007
rect 900 58976 1685 59004
rect 900 58964 906 58976
rect 1673 58973 1685 58976
rect 1719 58973 1731 59007
rect 1673 58967 1731 58973
rect 6886 58936 6914 59044
rect 19444 59013 19472 59180
rect 57333 59177 57345 59180
rect 57379 59177 57391 59211
rect 57333 59171 57391 59177
rect 19518 59100 19524 59152
rect 19576 59140 19582 59152
rect 19981 59143 20039 59149
rect 19981 59140 19993 59143
rect 19576 59112 19993 59140
rect 19576 59100 19582 59112
rect 19981 59109 19993 59112
rect 20027 59109 20039 59143
rect 19981 59103 20039 59109
rect 41325 59075 41383 59081
rect 41325 59072 41337 59075
rect 19536 59044 41337 59072
rect 19429 59007 19487 59013
rect 19429 58973 19441 59007
rect 19475 58973 19487 59007
rect 19429 58967 19487 58973
rect 19536 58936 19564 59044
rect 41325 59041 41337 59044
rect 41371 59041 41383 59075
rect 41782 59072 41788 59084
rect 41743 59044 41788 59072
rect 41325 59035 41383 59041
rect 41782 59032 41788 59044
rect 41840 59032 41846 59084
rect 58066 59072 58072 59084
rect 58027 59044 58072 59072
rect 58066 59032 58072 59044
rect 58124 59032 58130 59084
rect 19702 59004 19708 59016
rect 19663 58976 19708 59004
rect 19702 58964 19708 58976
rect 19760 58964 19766 59016
rect 19849 59007 19907 59013
rect 19849 58973 19861 59007
rect 19895 59004 19907 59007
rect 21450 59004 21456 59016
rect 19895 58976 21456 59004
rect 19895 58973 19907 58976
rect 19849 58967 19907 58973
rect 21450 58964 21456 58976
rect 21508 58964 21514 59016
rect 41230 58964 41236 59016
rect 41288 59004 41294 59016
rect 41509 59007 41567 59013
rect 41509 59004 41521 59007
rect 41288 58976 41521 59004
rect 41288 58964 41294 58976
rect 41509 58973 41521 58976
rect 41555 58973 41567 59007
rect 41874 59004 41880 59016
rect 41835 58976 41880 59004
rect 41509 58967 41567 58973
rect 41874 58964 41880 58976
rect 41932 58964 41938 59016
rect 57146 59004 57152 59016
rect 57107 58976 57152 59004
rect 57146 58964 57152 58976
rect 57204 58964 57210 59016
rect 57882 59004 57888 59016
rect 57843 58976 57888 59004
rect 57882 58964 57888 58976
rect 57940 58964 57946 59016
rect 6886 58908 19564 58936
rect 19613 58939 19671 58945
rect 19613 58905 19625 58939
rect 19659 58905 19671 58939
rect 19613 58899 19671 58905
rect 1765 58871 1823 58877
rect 1765 58837 1777 58871
rect 1811 58868 1823 58871
rect 17954 58868 17960 58880
rect 1811 58840 17960 58868
rect 1811 58837 1823 58840
rect 1765 58831 1823 58837
rect 17954 58828 17960 58840
rect 18012 58828 18018 58880
rect 19628 58868 19656 58899
rect 19978 58868 19984 58880
rect 19628 58840 19984 58868
rect 19978 58828 19984 58840
rect 20036 58828 20042 58880
rect 41141 58871 41199 58877
rect 41141 58837 41153 58871
rect 41187 58868 41199 58871
rect 42334 58868 42340 58880
rect 41187 58840 42340 58868
rect 41187 58837 41199 58840
rect 41141 58831 41199 58837
rect 42334 58828 42340 58840
rect 42392 58828 42398 58880
rect 1104 58778 58880 58800
rect 1104 58726 19574 58778
rect 19626 58726 19638 58778
rect 19690 58726 19702 58778
rect 19754 58726 19766 58778
rect 19818 58726 19830 58778
rect 19882 58726 50294 58778
rect 50346 58726 50358 58778
rect 50410 58726 50422 58778
rect 50474 58726 50486 58778
rect 50538 58726 50550 58778
rect 50602 58726 58880 58778
rect 1104 58704 58880 58726
rect 2038 58624 2044 58676
rect 2096 58664 2102 58676
rect 2096 58636 38700 58664
rect 2096 58624 2102 58636
rect 1578 58528 1584 58540
rect 1539 58500 1584 58528
rect 1578 58488 1584 58500
rect 1636 58488 1642 58540
rect 37918 58528 37924 58540
rect 37879 58500 37924 58528
rect 37918 58488 37924 58500
rect 37976 58488 37982 58540
rect 38010 58488 38016 58540
rect 38068 58528 38074 58540
rect 38289 58531 38347 58537
rect 38068 58500 38113 58528
rect 38068 58488 38074 58500
rect 38289 58497 38301 58531
rect 38335 58497 38347 58531
rect 38289 58491 38347 58497
rect 38565 58531 38623 58537
rect 38565 58497 38577 58531
rect 38611 58497 38623 58531
rect 38565 58491 38623 58497
rect 1857 58463 1915 58469
rect 1857 58429 1869 58463
rect 1903 58460 1915 58463
rect 4798 58460 4804 58472
rect 1903 58432 4804 58460
rect 1903 58429 1915 58432
rect 1857 58423 1915 58429
rect 4798 58420 4804 58432
rect 4856 58420 4862 58472
rect 36906 58420 36912 58472
rect 36964 58460 36970 58472
rect 38304 58460 38332 58491
rect 36964 58432 38332 58460
rect 36964 58420 36970 58432
rect 37182 58352 37188 58404
rect 37240 58392 37246 58404
rect 38580 58392 38608 58491
rect 38672 58460 38700 58636
rect 58158 58596 58164 58608
rect 38856 58568 45554 58596
rect 58119 58568 58164 58596
rect 38856 58537 38884 58568
rect 38841 58531 38899 58537
rect 38841 58497 38853 58531
rect 38887 58497 38899 58531
rect 41325 58531 41383 58537
rect 41325 58528 41337 58531
rect 38841 58491 38899 58497
rect 38948 58500 41337 58528
rect 38948 58460 38976 58500
rect 41325 58497 41337 58500
rect 41371 58497 41383 58531
rect 41506 58528 41512 58540
rect 41467 58500 41512 58528
rect 41325 58491 41383 58497
rect 41506 58488 41512 58500
rect 41564 58488 41570 58540
rect 41877 58531 41935 58537
rect 41877 58497 41889 58531
rect 41923 58528 41935 58531
rect 42610 58528 42616 58540
rect 41923 58500 42616 58528
rect 41923 58497 41935 58500
rect 41877 58491 41935 58497
rect 42610 58488 42616 58500
rect 42668 58488 42674 58540
rect 45526 58528 45554 58568
rect 58158 58556 58164 58568
rect 58216 58556 58222 58608
rect 56686 58528 56692 58540
rect 45526 58500 56692 58528
rect 56686 58488 56692 58500
rect 56744 58488 56750 58540
rect 40954 58460 40960 58472
rect 38672 58432 38976 58460
rect 40512 58432 40960 58460
rect 37240 58364 38608 58392
rect 37240 58352 37246 58364
rect 37550 58324 37556 58336
rect 37511 58296 37556 58324
rect 37550 58284 37556 58296
rect 37608 58284 37614 58336
rect 37918 58284 37924 58336
rect 37976 58324 37982 58336
rect 40512 58324 40540 58432
rect 40954 58420 40960 58432
rect 41012 58460 41018 58472
rect 41782 58460 41788 58472
rect 41012 58432 41788 58460
rect 41012 58420 41018 58432
rect 41782 58420 41788 58432
rect 41840 58420 41846 58472
rect 37976 58296 40540 58324
rect 41141 58327 41199 58333
rect 37976 58284 37982 58296
rect 41141 58293 41153 58327
rect 41187 58324 41199 58327
rect 41322 58324 41328 58336
rect 41187 58296 41328 58324
rect 41187 58293 41199 58296
rect 41141 58287 41199 58293
rect 41322 58284 41328 58296
rect 41380 58284 41386 58336
rect 52454 58284 52460 58336
rect 52512 58324 52518 58336
rect 58253 58327 58311 58333
rect 58253 58324 58265 58327
rect 52512 58296 58265 58324
rect 52512 58284 52518 58296
rect 58253 58293 58265 58296
rect 58299 58293 58311 58327
rect 58253 58287 58311 58293
rect 1104 58234 58880 58256
rect 1104 58182 4214 58234
rect 4266 58182 4278 58234
rect 4330 58182 4342 58234
rect 4394 58182 4406 58234
rect 4458 58182 4470 58234
rect 4522 58182 34934 58234
rect 34986 58182 34998 58234
rect 35050 58182 35062 58234
rect 35114 58182 35126 58234
rect 35178 58182 35190 58234
rect 35242 58182 58880 58234
rect 1104 58160 58880 58182
rect 35342 58080 35348 58132
rect 35400 58120 35406 58132
rect 41506 58120 41512 58132
rect 35400 58092 41512 58120
rect 35400 58080 35406 58092
rect 41506 58080 41512 58092
rect 41564 58080 41570 58132
rect 1578 57916 1584 57928
rect 1539 57888 1584 57916
rect 1578 57876 1584 57888
rect 1636 57876 1642 57928
rect 35618 57916 35624 57928
rect 35579 57888 35624 57916
rect 35618 57876 35624 57888
rect 35676 57876 35682 57928
rect 35897 57919 35955 57925
rect 35897 57885 35909 57919
rect 35943 57885 35955 57919
rect 35897 57879 35955 57885
rect 1857 57851 1915 57857
rect 1857 57817 1869 57851
rect 1903 57848 1915 57851
rect 10134 57848 10140 57860
rect 1903 57820 10140 57848
rect 1903 57817 1915 57820
rect 1857 57811 1915 57817
rect 10134 57808 10140 57820
rect 10192 57808 10198 57860
rect 34698 57808 34704 57860
rect 34756 57848 34762 57860
rect 35161 57851 35219 57857
rect 35161 57848 35173 57851
rect 34756 57820 35173 57848
rect 34756 57808 34762 57820
rect 35161 57817 35173 57820
rect 35207 57817 35219 57851
rect 35161 57811 35219 57817
rect 35710 57740 35716 57792
rect 35768 57780 35774 57792
rect 35912 57780 35940 57879
rect 35986 57876 35992 57928
rect 36044 57916 36050 57928
rect 36262 57916 36268 57928
rect 36044 57888 36089 57916
rect 36223 57888 36268 57916
rect 36044 57876 36050 57888
rect 36262 57876 36268 57888
rect 36320 57876 36326 57928
rect 36541 57919 36599 57925
rect 36541 57885 36553 57919
rect 36587 57916 36599 57919
rect 52454 57916 52460 57928
rect 36587 57888 52460 57916
rect 36587 57885 36599 57888
rect 36541 57879 36599 57885
rect 52454 57876 52460 57888
rect 52512 57876 52518 57928
rect 57974 57848 57980 57860
rect 57935 57820 57980 57848
rect 57974 57808 57980 57820
rect 58032 57808 58038 57860
rect 58066 57780 58072 57792
rect 35768 57752 35940 57780
rect 58027 57752 58072 57780
rect 35768 57740 35774 57752
rect 58066 57740 58072 57752
rect 58124 57740 58130 57792
rect 1104 57690 58880 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 58880 57690
rect 1104 57616 58880 57638
rect 34606 57468 34612 57520
rect 34664 57508 34670 57520
rect 35986 57508 35992 57520
rect 34664 57480 35992 57508
rect 34664 57468 34670 57480
rect 35986 57468 35992 57480
rect 36044 57468 36050 57520
rect 1578 57440 1584 57452
rect 1539 57412 1584 57440
rect 1578 57400 1584 57412
rect 1636 57400 1642 57452
rect 34514 57400 34520 57452
rect 34572 57440 34578 57452
rect 35713 57443 35771 57449
rect 35713 57440 35725 57443
rect 34572 57412 35725 57440
rect 34572 57400 34578 57412
rect 35713 57409 35725 57412
rect 35759 57409 35771 57443
rect 35713 57403 35771 57409
rect 35618 57332 35624 57384
rect 35676 57372 35682 57384
rect 35989 57375 36047 57381
rect 35989 57372 36001 57375
rect 35676 57344 36001 57372
rect 35676 57332 35682 57344
rect 35989 57341 36001 57344
rect 36035 57372 36047 57375
rect 37918 57372 37924 57384
rect 36035 57344 37924 57372
rect 36035 57341 36047 57344
rect 35989 57335 36047 57341
rect 37918 57332 37924 57344
rect 37976 57332 37982 57384
rect 4706 57264 4712 57316
rect 4764 57304 4770 57316
rect 15930 57304 15936 57316
rect 4764 57276 15936 57304
rect 4764 57264 4770 57276
rect 15930 57264 15936 57276
rect 15988 57264 15994 57316
rect 1762 57236 1768 57248
rect 1723 57208 1768 57236
rect 1762 57196 1768 57208
rect 1820 57196 1826 57248
rect 5534 57196 5540 57248
rect 5592 57236 5598 57248
rect 31478 57236 31484 57248
rect 5592 57208 31484 57236
rect 5592 57196 5598 57208
rect 31478 57196 31484 57208
rect 31536 57196 31542 57248
rect 1104 57146 58880 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 58880 57146
rect 1104 57072 58880 57094
rect 29362 56992 29368 57044
rect 29420 57032 29426 57044
rect 30650 57032 30656 57044
rect 29420 57004 30656 57032
rect 29420 56992 29426 57004
rect 30650 56992 30656 57004
rect 30708 56992 30714 57044
rect 17034 56856 17040 56908
rect 17092 56896 17098 56908
rect 22094 56896 22100 56908
rect 17092 56868 22100 56896
rect 17092 56856 17098 56868
rect 22094 56856 22100 56868
rect 22152 56856 22158 56908
rect 26878 56856 26884 56908
rect 26936 56896 26942 56908
rect 32861 56899 32919 56905
rect 32861 56896 32873 56899
rect 26936 56868 32873 56896
rect 26936 56856 26942 56868
rect 32861 56865 32873 56868
rect 32907 56865 32919 56899
rect 32861 56859 32919 56865
rect 32950 56856 32956 56908
rect 33008 56896 33014 56908
rect 33321 56899 33379 56905
rect 33321 56896 33333 56899
rect 33008 56868 33333 56896
rect 33008 56856 33014 56868
rect 33321 56865 33333 56868
rect 33367 56896 33379 56899
rect 33367 56868 35894 56896
rect 33367 56865 33379 56868
rect 33321 56859 33379 56865
rect 33042 56828 33048 56840
rect 33003 56800 33048 56828
rect 33042 56788 33048 56800
rect 33100 56788 33106 56840
rect 33413 56831 33471 56837
rect 33413 56797 33425 56831
rect 33459 56797 33471 56831
rect 35866 56828 35894 56868
rect 36262 56828 36268 56840
rect 35866 56800 36268 56828
rect 33413 56791 33471 56797
rect 1670 56760 1676 56772
rect 1631 56732 1676 56760
rect 1670 56720 1676 56732
rect 1728 56720 1734 56772
rect 2038 56760 2044 56772
rect 1999 56732 2044 56760
rect 2038 56720 2044 56732
rect 2096 56720 2102 56772
rect 33428 56760 33456 56791
rect 36262 56788 36268 56800
rect 36320 56788 36326 56840
rect 41322 56788 41328 56840
rect 41380 56828 41386 56840
rect 43990 56828 43996 56840
rect 41380 56800 43996 56828
rect 41380 56788 41386 56800
rect 43990 56788 43996 56800
rect 44048 56788 44054 56840
rect 57882 56828 57888 56840
rect 57843 56800 57888 56828
rect 57882 56788 57888 56800
rect 57940 56788 57946 56840
rect 49602 56760 49608 56772
rect 33428 56732 49608 56760
rect 49602 56720 49608 56732
rect 49660 56720 49666 56772
rect 51718 56720 51724 56772
rect 51776 56760 51782 56772
rect 58161 56763 58219 56769
rect 58161 56760 58173 56763
rect 51776 56732 58173 56760
rect 51776 56720 51782 56732
rect 58161 56729 58173 56732
rect 58207 56729 58219 56763
rect 58161 56723 58219 56729
rect 32490 56692 32496 56704
rect 32451 56664 32496 56692
rect 32490 56652 32496 56664
rect 32548 56652 32554 56704
rect 1104 56602 58880 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 58880 56602
rect 1104 56528 58880 56550
rect 1762 56448 1768 56500
rect 1820 56488 1826 56500
rect 1820 56460 29868 56488
rect 1820 56448 1826 56460
rect 2038 56380 2044 56432
rect 2096 56420 2102 56432
rect 2096 56392 22094 56420
rect 2096 56380 2102 56392
rect 22066 56216 22094 56392
rect 23566 56380 23572 56432
rect 23624 56420 23630 56432
rect 24210 56420 24216 56432
rect 23624 56392 24216 56420
rect 23624 56380 23630 56392
rect 24210 56380 24216 56392
rect 24268 56420 24274 56432
rect 24268 56392 24900 56420
rect 24268 56380 24274 56392
rect 24394 56352 24400 56364
rect 24355 56324 24400 56352
rect 24394 56312 24400 56324
rect 24452 56312 24458 56364
rect 24762 56352 24768 56364
rect 24723 56324 24768 56352
rect 24762 56312 24768 56324
rect 24820 56312 24826 56364
rect 24872 56361 24900 56392
rect 24857 56355 24915 56361
rect 24857 56321 24869 56355
rect 24903 56321 24915 56355
rect 24857 56315 24915 56321
rect 25314 56312 25320 56364
rect 25372 56352 25378 56364
rect 25372 56324 28994 56352
rect 25372 56312 25378 56324
rect 24026 56244 24032 56296
rect 24084 56284 24090 56296
rect 24305 56287 24363 56293
rect 24305 56284 24317 56287
rect 24084 56256 24317 56284
rect 24084 56244 24090 56256
rect 24305 56253 24317 56256
rect 24351 56253 24363 56287
rect 28966 56284 28994 56324
rect 29362 56312 29368 56364
rect 29420 56352 29426 56364
rect 29840 56361 29868 56460
rect 41230 56380 41236 56432
rect 41288 56420 41294 56432
rect 58158 56420 58164 56432
rect 41288 56392 41552 56420
rect 58119 56392 58164 56420
rect 41288 56380 41294 56392
rect 41524 56361 41552 56392
rect 58158 56380 58164 56392
rect 58216 56380 58222 56432
rect 29457 56355 29515 56361
rect 29457 56352 29469 56355
rect 29420 56324 29469 56352
rect 29420 56312 29426 56324
rect 29457 56321 29469 56324
rect 29503 56321 29515 56355
rect 29457 56315 29515 56321
rect 29825 56355 29883 56361
rect 29825 56321 29837 56355
rect 29871 56321 29883 56355
rect 41325 56355 41383 56361
rect 41325 56352 41337 56355
rect 29825 56315 29883 56321
rect 35866 56324 41337 56352
rect 29549 56287 29607 56293
rect 29549 56284 29561 56287
rect 28966 56256 29561 56284
rect 24305 56247 24363 56253
rect 29549 56253 29561 56256
rect 29595 56253 29607 56287
rect 29549 56247 29607 56253
rect 29730 56244 29736 56296
rect 29788 56284 29794 56296
rect 29917 56287 29975 56293
rect 29917 56284 29929 56287
rect 29788 56256 29929 56284
rect 29788 56244 29794 56256
rect 29917 56253 29929 56256
rect 29963 56253 29975 56287
rect 29917 56247 29975 56253
rect 35866 56216 35894 56324
rect 41325 56321 41337 56324
rect 41371 56321 41383 56355
rect 41325 56315 41383 56321
rect 41509 56355 41567 56361
rect 41509 56321 41521 56355
rect 41555 56321 41567 56355
rect 41509 56315 41567 56321
rect 41877 56355 41935 56361
rect 41877 56321 41889 56355
rect 41923 56352 41935 56355
rect 46842 56352 46848 56364
rect 41923 56324 46848 56352
rect 41923 56321 41935 56324
rect 41877 56315 41935 56321
rect 46842 56312 46848 56324
rect 46900 56312 46906 56364
rect 40954 56244 40960 56296
rect 41012 56284 41018 56296
rect 41785 56287 41843 56293
rect 41785 56284 41797 56287
rect 41012 56256 41797 56284
rect 41012 56244 41018 56256
rect 41785 56253 41797 56256
rect 41831 56253 41843 56287
rect 41785 56247 41843 56253
rect 22066 56188 35894 56216
rect 23842 56148 23848 56160
rect 23803 56120 23848 56148
rect 23842 56108 23848 56120
rect 23900 56108 23906 56160
rect 28905 56151 28963 56157
rect 28905 56117 28917 56151
rect 28951 56148 28963 56151
rect 28994 56148 29000 56160
rect 28951 56120 29000 56148
rect 28951 56117 28963 56120
rect 28905 56111 28963 56117
rect 28994 56108 29000 56120
rect 29052 56108 29058 56160
rect 41141 56151 41199 56157
rect 41141 56117 41153 56151
rect 41187 56148 41199 56151
rect 41322 56148 41328 56160
rect 41187 56120 41328 56148
rect 41187 56117 41199 56120
rect 41141 56111 41199 56117
rect 41322 56108 41328 56120
rect 41380 56108 41386 56160
rect 49602 56108 49608 56160
rect 49660 56148 49666 56160
rect 58253 56151 58311 56157
rect 58253 56148 58265 56151
rect 49660 56120 58265 56148
rect 49660 56108 49666 56120
rect 58253 56117 58265 56120
rect 58299 56117 58311 56151
rect 58253 56111 58311 56117
rect 1104 56058 58880 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 58880 56058
rect 1104 55984 58880 56006
rect 58342 55944 58348 55956
rect 58303 55916 58348 55944
rect 58342 55904 58348 55916
rect 58400 55904 58406 55956
rect 1762 55836 1768 55888
rect 1820 55876 1826 55888
rect 40862 55876 40868 55888
rect 1820 55848 40868 55876
rect 1820 55836 1826 55848
rect 40862 55836 40868 55848
rect 40920 55836 40926 55888
rect 31018 55808 31024 55820
rect 25240 55780 31024 55808
rect 25240 55749 25268 55780
rect 31018 55768 31024 55780
rect 31076 55768 31082 55820
rect 25225 55743 25283 55749
rect 25225 55709 25237 55743
rect 25271 55709 25283 55743
rect 25225 55703 25283 55709
rect 25314 55700 25320 55752
rect 25372 55740 25378 55752
rect 25593 55743 25651 55749
rect 25372 55712 25417 55740
rect 25372 55700 25378 55712
rect 25593 55709 25605 55743
rect 25639 55709 25651 55743
rect 25593 55703 25651 55709
rect 1670 55672 1676 55684
rect 1631 55644 1676 55672
rect 1670 55632 1676 55644
rect 1728 55632 1734 55684
rect 24302 55632 24308 55684
rect 24360 55672 24366 55684
rect 24581 55675 24639 55681
rect 24581 55672 24593 55675
rect 24360 55644 24593 55672
rect 24360 55632 24366 55644
rect 24581 55641 24593 55644
rect 24627 55641 24639 55675
rect 24581 55635 24639 55641
rect 1765 55607 1823 55613
rect 1765 55573 1777 55607
rect 1811 55604 1823 55607
rect 25608 55604 25636 55703
rect 25682 55700 25688 55752
rect 25740 55740 25746 55752
rect 29730 55740 29736 55752
rect 25740 55712 29736 55740
rect 25740 55700 25746 55712
rect 29730 55700 29736 55712
rect 29788 55740 29794 55752
rect 29788 55712 31754 55740
rect 29788 55700 29794 55712
rect 31726 55672 31754 55712
rect 35342 55672 35348 55684
rect 31726 55644 35348 55672
rect 35342 55632 35348 55644
rect 35400 55632 35406 55684
rect 1811 55576 25636 55604
rect 1811 55573 1823 55576
rect 1765 55567 1823 55573
rect 1104 55514 58880 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 58880 55514
rect 1104 55440 58880 55462
rect 1762 55400 1768 55412
rect 1723 55372 1768 55400
rect 1762 55360 1768 55372
rect 1820 55360 1826 55412
rect 41230 55400 41236 55412
rect 41064 55372 41236 55400
rect 40494 55292 40500 55344
rect 40552 55332 40558 55344
rect 41064 55341 41092 55372
rect 41230 55360 41236 55372
rect 41288 55360 41294 55412
rect 41049 55335 41107 55341
rect 41049 55332 41061 55335
rect 40552 55304 41061 55332
rect 40552 55292 40558 55304
rect 41049 55301 41061 55304
rect 41095 55301 41107 55335
rect 41049 55295 41107 55301
rect 41141 55335 41199 55341
rect 41141 55301 41153 55335
rect 41187 55332 41199 55335
rect 44174 55332 44180 55344
rect 41187 55304 44180 55332
rect 41187 55301 41199 55304
rect 41141 55295 41199 55301
rect 44174 55292 44180 55304
rect 44232 55292 44238 55344
rect 1578 55264 1584 55276
rect 1539 55236 1584 55264
rect 1578 55224 1584 55236
rect 1636 55224 1642 55276
rect 40862 55264 40868 55276
rect 40823 55236 40868 55264
rect 40862 55224 40868 55236
rect 40920 55224 40926 55276
rect 40954 55224 40960 55276
rect 41012 55264 41018 55276
rect 41230 55264 41236 55276
rect 41288 55273 41294 55276
rect 41012 55236 41236 55264
rect 41012 55224 41018 55236
rect 41230 55224 41236 55236
rect 41288 55227 41296 55273
rect 41434 55267 41492 55273
rect 41434 55233 41446 55267
rect 41480 55264 41492 55267
rect 42058 55264 42064 55276
rect 41480 55236 42064 55264
rect 41480 55233 41492 55236
rect 41434 55227 41492 55233
rect 41288 55224 41294 55227
rect 42058 55224 42064 55236
rect 42116 55224 42122 55276
rect 1104 54970 58880 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 58880 54970
rect 1104 54896 58880 54918
rect 24854 54788 24860 54800
rect 23400 54760 24860 54788
rect 23400 54729 23428 54760
rect 24854 54748 24860 54760
rect 24912 54788 24918 54800
rect 25314 54788 25320 54800
rect 24912 54760 25320 54788
rect 24912 54748 24918 54760
rect 25314 54748 25320 54760
rect 25372 54748 25378 54800
rect 23385 54723 23443 54729
rect 23385 54689 23397 54723
rect 23431 54689 23443 54723
rect 28718 54720 28724 54732
rect 23385 54683 23443 54689
rect 23492 54692 28724 54720
rect 23492 54661 23520 54692
rect 28718 54680 28724 54692
rect 28776 54680 28782 54732
rect 23477 54655 23535 54661
rect 23477 54621 23489 54655
rect 23523 54621 23535 54655
rect 23477 54615 23535 54621
rect 23845 54655 23903 54661
rect 23845 54621 23857 54655
rect 23891 54621 23903 54655
rect 23845 54615 23903 54621
rect 24029 54655 24087 54661
rect 24029 54621 24041 54655
rect 24075 54652 24087 54655
rect 25682 54652 25688 54664
rect 24075 54624 25688 54652
rect 24075 54621 24087 54624
rect 24029 54615 24087 54621
rect 1670 54584 1676 54596
rect 1631 54556 1676 54584
rect 1670 54544 1676 54556
rect 1728 54544 1734 54596
rect 22830 54584 22836 54596
rect 22791 54556 22836 54584
rect 22830 54544 22836 54556
rect 22888 54544 22894 54596
rect 1765 54519 1823 54525
rect 1765 54485 1777 54519
rect 1811 54516 1823 54519
rect 23860 54516 23888 54615
rect 25682 54612 25688 54624
rect 25740 54612 25746 54664
rect 58342 54652 58348 54664
rect 58303 54624 58348 54652
rect 58342 54612 58348 54624
rect 58400 54612 58406 54664
rect 1811 54488 23888 54516
rect 1811 54485 1823 54488
rect 1765 54479 1823 54485
rect 28074 54476 28080 54528
rect 28132 54516 28138 54528
rect 39390 54516 39396 54528
rect 28132 54488 39396 54516
rect 28132 54476 28138 54488
rect 39390 54476 39396 54488
rect 39448 54476 39454 54528
rect 1104 54426 58880 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 58880 54426
rect 1104 54352 58880 54374
rect 1578 54176 1584 54188
rect 1539 54148 1584 54176
rect 1578 54136 1584 54148
rect 1636 54136 1642 54188
rect 1762 53972 1768 53984
rect 1723 53944 1768 53972
rect 1762 53932 1768 53944
rect 1820 53932 1826 53984
rect 1104 53882 58880 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 58880 53882
rect 1104 53808 58880 53830
rect 40862 53700 40868 53712
rect 40823 53672 40868 53700
rect 40862 53660 40868 53672
rect 40920 53660 40926 53712
rect 41325 53635 41383 53641
rect 41325 53632 41337 53635
rect 40328 53604 41337 53632
rect 1762 53524 1768 53576
rect 1820 53564 1826 53576
rect 40328 53573 40356 53604
rect 41325 53601 41337 53604
rect 41371 53601 41383 53635
rect 41325 53595 41383 53601
rect 40313 53567 40371 53573
rect 40313 53564 40325 53567
rect 1820 53536 40325 53564
rect 1820 53524 1826 53536
rect 40313 53533 40325 53536
rect 40359 53533 40371 53567
rect 40313 53527 40371 53533
rect 40733 53567 40791 53573
rect 40733 53533 40745 53567
rect 40779 53564 40791 53567
rect 41230 53564 41236 53576
rect 40779 53536 41236 53564
rect 40779 53533 40791 53536
rect 40733 53527 40791 53533
rect 41230 53524 41236 53536
rect 41288 53524 41294 53576
rect 24946 53456 24952 53508
rect 25004 53496 25010 53508
rect 40494 53496 40500 53508
rect 25004 53468 40500 53496
rect 25004 53456 25010 53468
rect 40494 53456 40500 53468
rect 40552 53456 40558 53508
rect 40589 53499 40647 53505
rect 40589 53465 40601 53499
rect 40635 53496 40647 53499
rect 46106 53496 46112 53508
rect 40635 53468 46112 53496
rect 40635 53465 40647 53468
rect 40589 53459 40647 53465
rect 46106 53456 46112 53468
rect 46164 53456 46170 53508
rect 23474 53388 23480 53440
rect 23532 53428 23538 53440
rect 24578 53428 24584 53440
rect 23532 53400 24584 53428
rect 23532 53388 23538 53400
rect 24578 53388 24584 53400
rect 24636 53388 24642 53440
rect 1104 53338 58880 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 58880 53338
rect 1104 53264 58880 53286
rect 24946 53224 24952 53236
rect 23768 53196 24952 53224
rect 23768 53165 23796 53196
rect 24946 53184 24952 53196
rect 25004 53184 25010 53236
rect 23753 53159 23811 53165
rect 23753 53125 23765 53159
rect 23799 53125 23811 53159
rect 23753 53119 23811 53125
rect 23845 53159 23903 53165
rect 23845 53125 23857 53159
rect 23891 53156 23903 53159
rect 45370 53156 45376 53168
rect 23891 53128 45376 53156
rect 23891 53125 23903 53128
rect 23845 53119 23903 53125
rect 45370 53116 45376 53128
rect 45428 53116 45434 53168
rect 1670 53088 1676 53100
rect 1631 53060 1676 53088
rect 1670 53048 1676 53060
rect 1728 53048 1734 53100
rect 23569 53091 23627 53097
rect 23569 53088 23581 53091
rect 6886 53060 23581 53088
rect 1765 52887 1823 52893
rect 1765 52853 1777 52887
rect 1811 52884 1823 52887
rect 6886 52884 6914 53060
rect 23569 53057 23581 53060
rect 23615 53057 23627 53091
rect 23934 53088 23940 53100
rect 23847 53060 23940 53088
rect 23569 53051 23627 53057
rect 23934 53048 23940 53060
rect 23992 53048 23998 53100
rect 24578 53048 24584 53100
rect 24636 53088 24642 53100
rect 24636 53060 24681 53088
rect 24636 53048 24642 53060
rect 23952 53020 23980 53048
rect 24765 53023 24823 53029
rect 24765 53020 24777 53023
rect 23952 52992 24777 53020
rect 24765 52989 24777 52992
rect 24811 52989 24823 53023
rect 24765 52983 24823 52989
rect 1811 52856 6914 52884
rect 1811 52853 1823 52856
rect 1765 52847 1823 52853
rect 23934 52844 23940 52896
rect 23992 52884 23998 52896
rect 24121 52887 24179 52893
rect 24121 52884 24133 52887
rect 23992 52856 24133 52884
rect 23992 52844 23998 52856
rect 24121 52853 24133 52856
rect 24167 52853 24179 52887
rect 58342 52884 58348 52896
rect 58303 52856 58348 52884
rect 24121 52847 24179 52853
rect 58342 52844 58348 52856
rect 58400 52844 58406 52896
rect 1104 52794 58880 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 58880 52794
rect 1104 52720 58880 52742
rect 24946 52680 24952 52692
rect 24907 52652 24952 52680
rect 24946 52640 24952 52652
rect 25004 52640 25010 52692
rect 1857 52547 1915 52553
rect 1857 52513 1869 52547
rect 1903 52544 1915 52547
rect 10778 52544 10784 52556
rect 1903 52516 10784 52544
rect 1903 52513 1915 52516
rect 1857 52507 1915 52513
rect 10778 52504 10784 52516
rect 10836 52504 10842 52556
rect 1578 52476 1584 52488
rect 1539 52448 1584 52476
rect 1578 52436 1584 52448
rect 1636 52436 1642 52488
rect 20714 52368 20720 52420
rect 20772 52408 20778 52420
rect 24673 52411 24731 52417
rect 24673 52408 24685 52411
rect 20772 52380 24685 52408
rect 20772 52368 20778 52380
rect 24673 52377 24685 52380
rect 24719 52377 24731 52411
rect 24673 52371 24731 52377
rect 1104 52250 58880 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 58880 52250
rect 1104 52176 58880 52198
rect 1857 52071 1915 52077
rect 1857 52037 1869 52071
rect 1903 52068 1915 52071
rect 8205 52071 8263 52077
rect 8205 52068 8217 52071
rect 1903 52040 8217 52068
rect 1903 52037 1915 52040
rect 1857 52031 1915 52037
rect 8205 52037 8217 52040
rect 8251 52037 8263 52071
rect 8205 52031 8263 52037
rect 1670 52000 1676 52012
rect 1631 51972 1676 52000
rect 1670 51960 1676 51972
rect 1728 51960 1734 52012
rect 8018 52000 8024 52012
rect 7979 51972 8024 52000
rect 8018 51960 8024 51972
rect 8076 51960 8082 52012
rect 8297 52003 8355 52009
rect 8297 51969 8309 52003
rect 8343 52000 8355 52003
rect 20714 52000 20720 52012
rect 8343 51972 20720 52000
rect 8343 51969 8355 51972
rect 8297 51963 8355 51969
rect 4062 51892 4068 51944
rect 4120 51932 4126 51944
rect 8312 51932 8340 51963
rect 20714 51960 20720 51972
rect 20772 51960 20778 52012
rect 4120 51904 8340 51932
rect 4120 51892 4126 51904
rect 7834 51796 7840 51808
rect 7795 51768 7840 51796
rect 7834 51756 7840 51768
rect 7892 51756 7898 51808
rect 1104 51706 58880 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 58880 51706
rect 1104 51632 58880 51654
rect 20809 51595 20867 51601
rect 20809 51561 20821 51595
rect 20855 51592 20867 51595
rect 24118 51592 24124 51604
rect 20855 51564 24124 51592
rect 20855 51561 20867 51564
rect 20809 51555 20867 51561
rect 24118 51552 24124 51564
rect 24176 51552 24182 51604
rect 17862 51484 17868 51536
rect 17920 51524 17926 51536
rect 20993 51527 21051 51533
rect 20993 51524 21005 51527
rect 17920 51496 21005 51524
rect 17920 51484 17926 51496
rect 20993 51493 21005 51496
rect 21039 51493 21051 51527
rect 20993 51487 21051 51493
rect 20901 51459 20959 51465
rect 20901 51425 20913 51459
rect 20947 51456 20959 51459
rect 41138 51456 41144 51468
rect 20947 51428 41144 51456
rect 20947 51425 20959 51428
rect 20901 51419 20959 51425
rect 41138 51416 41144 51428
rect 41196 51416 41202 51468
rect 21085 51391 21143 51397
rect 21085 51357 21097 51391
rect 21131 51357 21143 51391
rect 21085 51351 21143 51357
rect 1670 51320 1676 51332
rect 1631 51292 1676 51320
rect 1670 51280 1676 51292
rect 1728 51280 1734 51332
rect 1857 51323 1915 51329
rect 1857 51289 1869 51323
rect 1903 51320 1915 51323
rect 3970 51320 3976 51332
rect 1903 51292 3976 51320
rect 1903 51289 1915 51292
rect 1857 51283 1915 51289
rect 3970 51280 3976 51292
rect 4028 51280 4034 51332
rect 20254 51280 20260 51332
rect 20312 51320 20318 51332
rect 21100 51320 21128 51351
rect 21174 51348 21180 51400
rect 21232 51388 21238 51400
rect 21269 51391 21327 51397
rect 21269 51388 21281 51391
rect 21232 51360 21281 51388
rect 21232 51348 21238 51360
rect 21269 51357 21281 51360
rect 21315 51357 21327 51391
rect 58342 51388 58348 51400
rect 58303 51360 58348 51388
rect 21269 51351 21327 51357
rect 58342 51348 58348 51360
rect 58400 51348 58406 51400
rect 20312 51292 21128 51320
rect 20312 51280 20318 51292
rect 20438 51212 20444 51264
rect 20496 51252 20502 51264
rect 20533 51255 20591 51261
rect 20533 51252 20545 51255
rect 20496 51224 20545 51252
rect 20496 51212 20502 51224
rect 20533 51221 20545 51224
rect 20579 51221 20591 51255
rect 20533 51215 20591 51221
rect 1104 51162 58880 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 58880 51162
rect 1104 51088 58880 51110
rect 4614 51048 4620 51060
rect 3712 51020 4620 51048
rect 3712 50921 3740 51020
rect 4614 51008 4620 51020
rect 4672 51008 4678 51060
rect 3970 50980 3976 50992
rect 3931 50952 3976 50980
rect 3970 50940 3976 50952
rect 4028 50940 4034 50992
rect 3697 50915 3755 50921
rect 3697 50881 3709 50915
rect 3743 50881 3755 50915
rect 3697 50875 3755 50881
rect 3881 50915 3939 50921
rect 3881 50881 3893 50915
rect 3927 50881 3939 50915
rect 3881 50875 3939 50881
rect 2590 50804 2596 50856
rect 2648 50844 2654 50856
rect 3896 50844 3924 50875
rect 4062 50872 4068 50924
rect 4120 50921 4126 50924
rect 4120 50912 4128 50921
rect 4120 50884 4165 50912
rect 4120 50875 4128 50884
rect 4120 50872 4126 50875
rect 2648 50816 3924 50844
rect 2648 50804 2654 50816
rect 4249 50711 4307 50717
rect 4249 50677 4261 50711
rect 4295 50708 4307 50711
rect 6270 50708 6276 50720
rect 4295 50680 6276 50708
rect 4295 50677 4307 50680
rect 4249 50671 4307 50677
rect 6270 50668 6276 50680
rect 6328 50668 6334 50720
rect 1104 50618 58880 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 58880 50618
rect 1104 50544 58880 50566
rect 29914 50396 29920 50448
rect 29972 50436 29978 50448
rect 41782 50436 41788 50448
rect 29972 50408 41788 50436
rect 29972 50396 29978 50408
rect 41782 50396 41788 50408
rect 41840 50396 41846 50448
rect 10134 50328 10140 50380
rect 10192 50368 10198 50380
rect 29822 50368 29828 50380
rect 10192 50340 29828 50368
rect 10192 50328 10198 50340
rect 29822 50328 29828 50340
rect 29880 50328 29886 50380
rect 39482 50328 39488 50380
rect 39540 50368 39546 50380
rect 55766 50368 55772 50380
rect 39540 50340 55772 50368
rect 39540 50328 39546 50340
rect 55766 50328 55772 50340
rect 55824 50328 55830 50380
rect 57422 50260 57428 50312
rect 57480 50300 57486 50312
rect 57885 50303 57943 50309
rect 57885 50300 57897 50303
rect 57480 50272 57897 50300
rect 57480 50260 57486 50272
rect 57885 50269 57897 50272
rect 57931 50269 57943 50303
rect 57885 50263 57943 50269
rect 1670 50232 1676 50244
rect 1631 50204 1676 50232
rect 1670 50192 1676 50204
rect 1728 50192 1734 50244
rect 1857 50235 1915 50241
rect 1857 50201 1869 50235
rect 1903 50232 1915 50235
rect 2038 50232 2044 50244
rect 1903 50204 2044 50232
rect 1903 50201 1915 50204
rect 1857 50195 1915 50201
rect 2038 50192 2044 50204
rect 2096 50192 2102 50244
rect 58161 50235 58219 50241
rect 58161 50232 58173 50235
rect 57900 50204 58173 50232
rect 57900 50176 57928 50204
rect 58161 50201 58173 50204
rect 58207 50201 58219 50235
rect 58161 50195 58219 50201
rect 57882 50124 57888 50176
rect 57940 50124 57946 50176
rect 1104 50074 58880 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 58880 50074
rect 1104 50000 58880 50022
rect 1578 49824 1584 49836
rect 1539 49796 1584 49824
rect 1578 49784 1584 49796
rect 1636 49784 1642 49836
rect 13078 49756 13084 49768
rect 1780 49728 13084 49756
rect 1780 49697 1808 49728
rect 13078 49716 13084 49728
rect 13136 49716 13142 49768
rect 1765 49691 1823 49697
rect 1765 49657 1777 49691
rect 1811 49657 1823 49691
rect 1765 49651 1823 49657
rect 1104 49530 58880 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 58880 49530
rect 1104 49456 58880 49478
rect 1578 49212 1584 49224
rect 1539 49184 1584 49212
rect 1578 49172 1584 49184
rect 1636 49172 1642 49224
rect 57974 49144 57980 49156
rect 57935 49116 57980 49144
rect 57974 49104 57980 49116
rect 58032 49104 58038 49156
rect 58345 49147 58403 49153
rect 58345 49113 58357 49147
rect 58391 49144 58403 49147
rect 59078 49144 59084 49156
rect 58391 49116 59084 49144
rect 58391 49113 58403 49116
rect 58345 49107 58403 49113
rect 59078 49104 59084 49116
rect 59136 49104 59142 49156
rect 1765 49079 1823 49085
rect 1765 49045 1777 49079
rect 1811 49076 1823 49079
rect 18598 49076 18604 49088
rect 1811 49048 18604 49076
rect 1811 49045 1823 49048
rect 1765 49039 1823 49045
rect 18598 49036 18604 49048
rect 18656 49036 18662 49088
rect 1104 48986 58880 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 58880 48986
rect 1104 48912 58880 48934
rect 1670 48736 1676 48748
rect 1631 48708 1676 48736
rect 1670 48696 1676 48708
rect 1728 48696 1734 48748
rect 1857 48603 1915 48609
rect 1857 48569 1869 48603
rect 1903 48600 1915 48603
rect 1946 48600 1952 48612
rect 1903 48572 1952 48600
rect 1903 48569 1915 48572
rect 1857 48563 1915 48569
rect 1946 48560 1952 48572
rect 2004 48560 2010 48612
rect 1104 48442 58880 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 58880 48442
rect 1104 48368 58880 48390
rect 2593 48263 2651 48269
rect 2593 48229 2605 48263
rect 2639 48260 2651 48263
rect 17862 48260 17868 48272
rect 2639 48232 17868 48260
rect 2639 48229 2651 48232
rect 2593 48223 2651 48229
rect 17862 48220 17868 48232
rect 17920 48220 17926 48272
rect 2866 48192 2872 48204
rect 2240 48164 2872 48192
rect 2038 48124 2044 48136
rect 1999 48096 2044 48124
rect 2038 48084 2044 48096
rect 2096 48084 2102 48136
rect 2240 48133 2268 48164
rect 2866 48152 2872 48164
rect 2924 48192 2930 48204
rect 4062 48192 4068 48204
rect 2924 48164 4068 48192
rect 2924 48152 2930 48164
rect 4062 48152 4068 48164
rect 4120 48152 4126 48204
rect 2225 48127 2283 48133
rect 2225 48093 2237 48127
rect 2271 48093 2283 48127
rect 2406 48124 2412 48136
rect 2464 48133 2470 48136
rect 2372 48096 2412 48124
rect 2225 48087 2283 48093
rect 2406 48084 2412 48096
rect 2464 48087 2472 48133
rect 2464 48084 2470 48087
rect 57790 48084 57796 48136
rect 57848 48124 57854 48136
rect 57885 48127 57943 48133
rect 57885 48124 57897 48127
rect 57848 48096 57897 48124
rect 57848 48084 57854 48096
rect 57885 48093 57897 48096
rect 57931 48093 57943 48127
rect 57885 48087 57943 48093
rect 2317 48059 2375 48065
rect 2317 48025 2329 48059
rect 2363 48025 2375 48059
rect 58158 48056 58164 48068
rect 58119 48028 58164 48056
rect 2317 48019 2375 48025
rect 1854 47948 1860 48000
rect 1912 47988 1918 48000
rect 2332 47988 2360 48019
rect 58158 48016 58164 48028
rect 58216 48016 58222 48068
rect 1912 47960 2360 47988
rect 1912 47948 1918 47960
rect 1104 47898 58880 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 58880 47898
rect 1104 47824 58880 47846
rect 53374 47744 53380 47796
rect 53432 47784 53438 47796
rect 58066 47784 58072 47796
rect 53432 47756 58072 47784
rect 53432 47744 53438 47756
rect 58066 47744 58072 47756
rect 58124 47744 58130 47796
rect 1670 47648 1676 47660
rect 1631 47620 1676 47648
rect 1670 47608 1676 47620
rect 1728 47608 1734 47660
rect 25406 47608 25412 47660
rect 25464 47648 25470 47660
rect 40126 47648 40132 47660
rect 25464 47620 40132 47648
rect 25464 47608 25470 47620
rect 40126 47608 40132 47620
rect 40184 47608 40190 47660
rect 58066 47648 58072 47660
rect 58027 47620 58072 47648
rect 58066 47608 58072 47620
rect 58124 47608 58130 47660
rect 10778 47540 10784 47592
rect 10836 47580 10842 47592
rect 26234 47580 26240 47592
rect 10836 47552 26240 47580
rect 10836 47540 10842 47552
rect 26234 47540 26240 47552
rect 26292 47540 26298 47592
rect 35802 47540 35808 47592
rect 35860 47580 35866 47592
rect 53190 47580 53196 47592
rect 35860 47552 53196 47580
rect 35860 47540 35866 47552
rect 53190 47540 53196 47552
rect 53248 47540 53254 47592
rect 1857 47515 1915 47521
rect 1857 47481 1869 47515
rect 1903 47512 1915 47515
rect 6178 47512 6184 47524
rect 1903 47484 6184 47512
rect 1903 47481 1915 47484
rect 1857 47475 1915 47481
rect 6178 47472 6184 47484
rect 6236 47472 6242 47524
rect 58253 47447 58311 47453
rect 58253 47413 58265 47447
rect 58299 47444 58311 47447
rect 58802 47444 58808 47456
rect 58299 47416 58808 47444
rect 58299 47413 58311 47416
rect 58253 47407 58311 47413
rect 58802 47404 58808 47416
rect 58860 47404 58866 47456
rect 1104 47354 58880 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 58880 47354
rect 1104 47280 58880 47302
rect 1578 47036 1584 47048
rect 1539 47008 1584 47036
rect 1578 46996 1584 47008
rect 1636 46996 1642 47048
rect 10318 46968 10324 46980
rect 1780 46940 10324 46968
rect 1780 46909 1808 46940
rect 10318 46928 10324 46940
rect 10376 46928 10382 46980
rect 32582 46928 32588 46980
rect 32640 46968 32646 46980
rect 37918 46968 37924 46980
rect 32640 46940 37924 46968
rect 32640 46928 32646 46940
rect 37918 46928 37924 46940
rect 37976 46928 37982 46980
rect 1765 46903 1823 46909
rect 1765 46869 1777 46903
rect 1811 46869 1823 46903
rect 1765 46863 1823 46869
rect 1104 46810 58880 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 58880 46810
rect 1104 46736 58880 46758
rect 1578 46560 1584 46572
rect 1539 46532 1584 46560
rect 1578 46520 1584 46532
rect 1636 46520 1642 46572
rect 1765 46359 1823 46365
rect 1765 46325 1777 46359
rect 1811 46356 1823 46359
rect 36354 46356 36360 46368
rect 1811 46328 36360 46356
rect 1811 46325 1823 46328
rect 1765 46319 1823 46325
rect 36354 46316 36360 46328
rect 36412 46316 36418 46368
rect 1104 46266 58880 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 58880 46266
rect 1104 46192 58880 46214
rect 58158 46016 58164 46028
rect 58119 45988 58164 46016
rect 58158 45976 58164 45988
rect 58216 45976 58222 46028
rect 57698 45908 57704 45960
rect 57756 45948 57762 45960
rect 57885 45951 57943 45957
rect 57885 45948 57897 45951
rect 57756 45920 57897 45948
rect 57756 45908 57762 45920
rect 57885 45917 57897 45920
rect 57931 45917 57943 45951
rect 57885 45911 57943 45917
rect 1670 45880 1676 45892
rect 1631 45852 1676 45880
rect 1670 45840 1676 45852
rect 1728 45840 1734 45892
rect 1765 45815 1823 45821
rect 1765 45781 1777 45815
rect 1811 45812 1823 45815
rect 15194 45812 15200 45824
rect 1811 45784 15200 45812
rect 1811 45781 1823 45784
rect 1765 45775 1823 45781
rect 15194 45772 15200 45784
rect 15252 45772 15258 45824
rect 1104 45722 58880 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 58880 45722
rect 1104 45648 58880 45670
rect 15194 45500 15200 45552
rect 15252 45540 15258 45552
rect 20714 45540 20720 45552
rect 15252 45512 17172 45540
rect 15252 45500 15258 45512
rect 17144 45481 17172 45512
rect 17328 45512 20720 45540
rect 17328 45481 17356 45512
rect 20714 45500 20720 45512
rect 20772 45500 20778 45552
rect 35342 45500 35348 45552
rect 35400 45540 35406 45552
rect 36541 45543 36599 45549
rect 36541 45540 36553 45543
rect 35400 45512 36553 45540
rect 35400 45500 35406 45512
rect 36541 45509 36553 45512
rect 36587 45509 36599 45543
rect 38197 45543 38255 45549
rect 38197 45540 38209 45543
rect 36541 45503 36599 45509
rect 37476 45512 38209 45540
rect 37476 45484 37504 45512
rect 38197 45509 38209 45512
rect 38243 45509 38255 45543
rect 38197 45503 38255 45509
rect 38289 45543 38347 45549
rect 38289 45509 38301 45543
rect 38335 45540 38347 45543
rect 38335 45512 45554 45540
rect 38335 45509 38347 45512
rect 38289 45503 38347 45509
rect 17037 45475 17095 45481
rect 17037 45441 17049 45475
rect 17083 45441 17095 45475
rect 17037 45435 17095 45441
rect 17130 45475 17188 45481
rect 17130 45441 17142 45475
rect 17176 45441 17188 45475
rect 17130 45435 17188 45441
rect 17313 45475 17371 45481
rect 17313 45441 17325 45475
rect 17359 45441 17371 45475
rect 17313 45435 17371 45441
rect 17052 45268 17080 45435
rect 17402 45432 17408 45484
rect 17460 45472 17466 45484
rect 17543 45475 17601 45481
rect 17460 45444 17502 45472
rect 17460 45432 17466 45444
rect 17543 45441 17555 45475
rect 17589 45472 17601 45475
rect 23474 45472 23480 45484
rect 17589 45444 23480 45472
rect 17589 45441 17601 45444
rect 17543 45435 17601 45441
rect 23474 45432 23480 45444
rect 23532 45472 23538 45484
rect 24210 45472 24216 45484
rect 23532 45444 24216 45472
rect 23532 45432 23538 45444
rect 24210 45432 24216 45444
rect 24268 45432 24274 45484
rect 36354 45472 36360 45484
rect 36315 45444 36360 45472
rect 36354 45432 36360 45444
rect 36412 45432 36418 45484
rect 36630 45432 36636 45484
rect 36688 45472 36694 45484
rect 36771 45475 36829 45481
rect 36688 45444 36733 45472
rect 36688 45432 36694 45444
rect 36771 45441 36783 45475
rect 36817 45472 36829 45475
rect 37458 45472 37464 45484
rect 36817 45444 37464 45472
rect 36817 45441 36829 45444
rect 36771 45435 36829 45441
rect 37458 45432 37464 45444
rect 37516 45432 37522 45484
rect 37737 45475 37795 45481
rect 37737 45441 37749 45475
rect 37783 45472 37795 45475
rect 38010 45472 38016 45484
rect 37783 45444 38016 45472
rect 37783 45441 37795 45444
rect 37737 45435 37795 45441
rect 38010 45432 38016 45444
rect 38068 45432 38074 45484
rect 38386 45475 38444 45481
rect 38386 45472 38398 45475
rect 38120 45444 38398 45472
rect 35986 45364 35992 45416
rect 36044 45404 36050 45416
rect 37182 45404 37188 45416
rect 36044 45376 37188 45404
rect 36044 45364 36050 45376
rect 37182 45364 37188 45376
rect 37240 45404 37246 45416
rect 38120 45404 38148 45444
rect 38386 45441 38398 45444
rect 38432 45441 38444 45475
rect 45526 45472 45554 45512
rect 57054 45472 57060 45484
rect 45526 45444 57060 45472
rect 38386 45435 38444 45441
rect 57054 45432 57060 45444
rect 57112 45432 57118 45484
rect 58066 45472 58072 45484
rect 58027 45444 58072 45472
rect 58066 45432 58072 45444
rect 58124 45432 58130 45484
rect 37240 45376 38148 45404
rect 37240 45364 37246 45376
rect 36906 45336 36912 45348
rect 17512 45308 26234 45336
rect 36867 45308 36912 45336
rect 17512 45268 17540 45308
rect 17678 45268 17684 45280
rect 17052 45240 17540 45268
rect 17639 45240 17684 45268
rect 17678 45228 17684 45240
rect 17736 45228 17742 45280
rect 26206 45268 26234 45308
rect 36906 45296 36912 45308
rect 36964 45296 36970 45348
rect 38565 45339 38623 45345
rect 38565 45336 38577 45339
rect 37016 45308 38577 45336
rect 37016 45268 37044 45308
rect 38565 45305 38577 45308
rect 38611 45305 38623 45339
rect 38565 45299 38623 45305
rect 26206 45240 37044 45268
rect 58253 45271 58311 45277
rect 58253 45237 58265 45271
rect 58299 45268 58311 45271
rect 58618 45268 58624 45280
rect 58299 45240 58624 45268
rect 58299 45237 58311 45240
rect 58253 45231 58311 45237
rect 58618 45228 58624 45240
rect 58676 45228 58682 45280
rect 1104 45178 58880 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 58880 45178
rect 1104 45104 58880 45126
rect 1578 44860 1584 44872
rect 1539 44832 1584 44860
rect 1578 44820 1584 44832
rect 1636 44820 1642 44872
rect 56778 44820 56784 44872
rect 56836 44860 56842 44872
rect 56965 44863 57023 44869
rect 56965 44860 56977 44863
rect 56836 44832 56977 44860
rect 56836 44820 56842 44832
rect 56965 44829 56977 44832
rect 57011 44829 57023 44863
rect 56965 44823 57023 44829
rect 1857 44795 1915 44801
rect 1857 44761 1869 44795
rect 1903 44792 1915 44795
rect 36814 44792 36820 44804
rect 1903 44764 36820 44792
rect 1903 44761 1915 44764
rect 1857 44755 1915 44761
rect 36814 44752 36820 44764
rect 36872 44752 36878 44804
rect 57238 44792 57244 44804
rect 57199 44764 57244 44792
rect 57238 44752 57244 44764
rect 57296 44752 57302 44804
rect 57882 44752 57888 44804
rect 57940 44792 57946 44804
rect 57977 44795 58035 44801
rect 57977 44792 57989 44795
rect 57940 44764 57989 44792
rect 57940 44752 57946 44764
rect 57977 44761 57989 44764
rect 58023 44761 58035 44795
rect 57977 44755 58035 44761
rect 58345 44795 58403 44801
rect 58345 44761 58357 44795
rect 58391 44792 58403 44795
rect 58710 44792 58716 44804
rect 58391 44764 58716 44792
rect 58391 44761 58403 44764
rect 58345 44755 58403 44761
rect 58710 44752 58716 44764
rect 58768 44752 58774 44804
rect 1104 44634 58880 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 58880 44634
rect 1104 44560 58880 44582
rect 34054 44480 34060 44532
rect 34112 44520 34118 44532
rect 34112 44492 41414 44520
rect 34112 44480 34118 44492
rect 9214 44412 9220 44464
rect 9272 44452 9278 44464
rect 34333 44455 34391 44461
rect 34333 44452 34345 44455
rect 9272 44424 34345 44452
rect 9272 44412 9278 44424
rect 34333 44421 34345 44424
rect 34379 44421 34391 44455
rect 34333 44415 34391 44421
rect 1670 44384 1676 44396
rect 1631 44356 1676 44384
rect 1670 44344 1676 44356
rect 1728 44344 1734 44396
rect 34054 44384 34060 44396
rect 34015 44356 34060 44384
rect 34054 44344 34060 44356
rect 34112 44344 34118 44396
rect 34146 44344 34152 44396
rect 34204 44384 34210 44396
rect 34241 44387 34299 44393
rect 34241 44384 34253 44387
rect 34204 44356 34253 44384
rect 34204 44344 34210 44356
rect 34241 44353 34253 44356
rect 34287 44353 34299 44387
rect 34430 44387 34488 44393
rect 34430 44384 34442 44387
rect 34241 44347 34299 44353
rect 34348 44356 34442 44384
rect 21450 44276 21456 44328
rect 21508 44316 21514 44328
rect 34348 44316 34376 44356
rect 34430 44353 34442 44356
rect 34476 44353 34488 44387
rect 41386 44384 41414 44492
rect 45738 44384 45744 44396
rect 41386 44356 45744 44384
rect 34430 44347 34488 44353
rect 45738 44344 45744 44356
rect 45796 44344 45802 44396
rect 21508 44288 34376 44316
rect 21508 44276 21514 44288
rect 1857 44251 1915 44257
rect 1857 44217 1869 44251
rect 1903 44248 1915 44251
rect 9582 44248 9588 44260
rect 1903 44220 9588 44248
rect 1903 44217 1915 44220
rect 1857 44211 1915 44217
rect 9582 44208 9588 44220
rect 9640 44208 9646 44260
rect 34606 44248 34612 44260
rect 34567 44220 34612 44248
rect 34606 44208 34612 44220
rect 34664 44208 34670 44260
rect 1104 44090 58880 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 58880 44090
rect 1104 44016 58880 44038
rect 34238 43908 34244 43920
rect 34199 43880 34244 43908
rect 34238 43868 34244 43880
rect 34296 43868 34302 43920
rect 9582 43800 9588 43852
rect 9640 43840 9646 43852
rect 9640 43812 26234 43840
rect 9640 43800 9646 43812
rect 26206 43772 26234 43812
rect 33689 43775 33747 43781
rect 33689 43772 33701 43775
rect 26206 43744 33701 43772
rect 33689 43741 33701 43744
rect 33735 43741 33747 43775
rect 34062 43775 34120 43781
rect 34062 43772 34074 43775
rect 33689 43735 33747 43741
rect 33796 43744 34074 43772
rect 1670 43704 1676 43716
rect 1631 43676 1676 43704
rect 1670 43664 1676 43676
rect 1728 43664 1734 43716
rect 33042 43664 33048 43716
rect 33100 43704 33106 43716
rect 33796 43704 33824 43744
rect 34062 43741 34074 43744
rect 34108 43741 34120 43775
rect 34062 43735 34120 43741
rect 57606 43732 57612 43784
rect 57664 43772 57670 43784
rect 57885 43775 57943 43781
rect 57885 43772 57897 43775
rect 57664 43744 57897 43772
rect 57664 43732 57670 43744
rect 57885 43741 57897 43744
rect 57931 43741 57943 43775
rect 57885 43735 57943 43741
rect 33100 43676 33824 43704
rect 33873 43707 33931 43713
rect 33100 43664 33106 43676
rect 33873 43673 33885 43707
rect 33919 43673 33931 43707
rect 33873 43667 33931 43673
rect 33965 43707 34023 43713
rect 33965 43673 33977 43707
rect 34011 43704 34023 43707
rect 35894 43704 35900 43716
rect 34011 43676 35900 43704
rect 34011 43673 34023 43676
rect 33965 43667 34023 43673
rect 1765 43639 1823 43645
rect 1765 43605 1777 43639
rect 1811 43636 1823 43639
rect 32306 43636 32312 43648
rect 1811 43608 32312 43636
rect 1811 43605 1823 43608
rect 1765 43599 1823 43605
rect 32306 43596 32312 43608
rect 32364 43596 32370 43648
rect 33686 43596 33692 43648
rect 33744 43636 33750 43648
rect 33888 43636 33916 43667
rect 35894 43664 35900 43676
rect 35952 43664 35958 43716
rect 58158 43704 58164 43716
rect 58119 43676 58164 43704
rect 58158 43664 58164 43676
rect 58216 43664 58222 43716
rect 35342 43636 35348 43648
rect 33744 43608 35348 43636
rect 33744 43596 33750 43608
rect 35342 43596 35348 43608
rect 35400 43596 35406 43648
rect 1104 43546 58880 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 58880 43546
rect 1104 43472 58880 43494
rect 33226 43432 33232 43444
rect 32508 43404 33232 43432
rect 32508 43373 32536 43404
rect 33226 43392 33232 43404
rect 33284 43432 33290 43444
rect 33686 43432 33692 43444
rect 33284 43404 33692 43432
rect 33284 43392 33290 43404
rect 33686 43392 33692 43404
rect 33744 43392 33750 43444
rect 32493 43367 32551 43373
rect 32493 43333 32505 43367
rect 32539 43333 32551 43367
rect 32493 43327 32551 43333
rect 32585 43367 32643 43373
rect 32585 43333 32597 43367
rect 32631 43364 32643 43367
rect 54846 43364 54852 43376
rect 32631 43336 54852 43364
rect 32631 43333 32643 43336
rect 32585 43327 32643 43333
rect 54846 43324 54852 43336
rect 54904 43324 54910 43376
rect 1578 43296 1584 43308
rect 1539 43268 1584 43296
rect 1578 43256 1584 43268
rect 1636 43256 1642 43308
rect 32306 43296 32312 43308
rect 32267 43268 32312 43296
rect 32306 43256 32312 43268
rect 32364 43256 32370 43308
rect 32766 43305 32772 43308
rect 32729 43299 32772 43305
rect 32729 43265 32741 43299
rect 32729 43259 32772 43265
rect 32766 43256 32772 43259
rect 32824 43256 32830 43308
rect 1762 43092 1768 43104
rect 1723 43064 1768 43092
rect 1762 43052 1768 43064
rect 1820 43052 1826 43104
rect 32861 43095 32919 43101
rect 32861 43061 32873 43095
rect 32907 43092 32919 43095
rect 32950 43092 32956 43104
rect 32907 43064 32956 43092
rect 32907 43061 32919 43064
rect 32861 43055 32919 43061
rect 32950 43052 32956 43064
rect 33008 43052 33014 43104
rect 1104 43002 58880 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 58880 43002
rect 1104 42928 58880 42950
rect 32766 42712 32772 42764
rect 32824 42752 32830 42764
rect 32824 42724 37688 42752
rect 32824 42712 32830 42724
rect 33042 42684 33048 42696
rect 33003 42656 33048 42684
rect 33042 42644 33048 42656
rect 33100 42644 33106 42696
rect 33134 42644 33140 42696
rect 33192 42684 33198 42696
rect 33413 42687 33471 42693
rect 33192 42656 33237 42684
rect 33192 42644 33198 42656
rect 33413 42653 33425 42687
rect 33459 42653 33471 42687
rect 33686 42684 33692 42696
rect 33647 42656 33692 42684
rect 33413 42647 33471 42653
rect 32677 42551 32735 42557
rect 32677 42517 32689 42551
rect 32723 42548 32735 42551
rect 32766 42548 32772 42560
rect 32723 42520 32772 42548
rect 32723 42517 32735 42520
rect 32677 42511 32735 42517
rect 32766 42508 32772 42520
rect 32824 42508 32830 42560
rect 33428 42548 33456 42647
rect 33686 42644 33692 42656
rect 33744 42644 33750 42696
rect 33870 42684 33876 42696
rect 33831 42656 33876 42684
rect 33870 42644 33876 42656
rect 33928 42644 33934 42696
rect 34238 42644 34244 42696
rect 34296 42684 34302 42696
rect 34790 42684 34796 42696
rect 34296 42656 34796 42684
rect 34296 42644 34302 42656
rect 34790 42644 34796 42656
rect 34848 42644 34854 42696
rect 37274 42684 37280 42696
rect 37235 42656 37280 42684
rect 37274 42644 37280 42656
rect 37332 42644 37338 42696
rect 37660 42693 37688 42724
rect 37645 42687 37703 42693
rect 37645 42653 37657 42687
rect 37691 42653 37703 42687
rect 37645 42647 37703 42653
rect 37458 42616 37464 42628
rect 37419 42588 37464 42616
rect 37458 42576 37464 42588
rect 37516 42576 37522 42628
rect 37553 42619 37611 42625
rect 37553 42585 37565 42619
rect 37599 42616 37611 42619
rect 54294 42616 54300 42628
rect 37599 42588 54300 42616
rect 37599 42585 37611 42588
rect 37553 42579 37611 42585
rect 54294 42576 54300 42588
rect 54352 42576 54358 42628
rect 57054 42616 57060 42628
rect 57015 42588 57060 42616
rect 57054 42576 57060 42588
rect 57112 42576 57118 42628
rect 57974 42616 57980 42628
rect 57935 42588 57980 42616
rect 57974 42576 57980 42588
rect 58032 42576 58038 42628
rect 58342 42616 58348 42628
rect 58303 42588 58348 42616
rect 58342 42576 58348 42588
rect 58400 42576 58406 42628
rect 37829 42551 37887 42557
rect 37829 42548 37841 42551
rect 33428 42520 37841 42548
rect 37829 42517 37841 42520
rect 37875 42517 37887 42551
rect 57330 42548 57336 42560
rect 57291 42520 57336 42548
rect 37829 42511 37887 42517
rect 57330 42508 57336 42520
rect 57388 42508 57394 42560
rect 1104 42458 58880 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 58880 42458
rect 1104 42384 58880 42406
rect 1762 42304 1768 42356
rect 1820 42344 1826 42356
rect 33870 42344 33876 42356
rect 1820 42316 33876 42344
rect 1820 42304 1826 42316
rect 33870 42304 33876 42316
rect 33928 42304 33934 42356
rect 1578 42208 1584 42220
rect 1539 42180 1584 42208
rect 1578 42168 1584 42180
rect 1636 42168 1642 42220
rect 1765 42007 1823 42013
rect 1765 41973 1777 42007
rect 1811 42004 1823 42007
rect 2130 42004 2136 42016
rect 1811 41976 2136 42004
rect 1811 41973 1823 41976
rect 1765 41967 1823 41973
rect 2130 41964 2136 41976
rect 2188 41964 2194 42016
rect 1104 41914 58880 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 58880 41914
rect 1104 41840 58880 41862
rect 54662 41556 54668 41608
rect 54720 41596 54726 41608
rect 56965 41599 57023 41605
rect 56965 41596 56977 41599
rect 54720 41568 56977 41596
rect 54720 41556 54726 41568
rect 56965 41565 56977 41568
rect 57011 41565 57023 41599
rect 56965 41559 57023 41565
rect 1670 41528 1676 41540
rect 1631 41500 1676 41528
rect 1670 41488 1676 41500
rect 1728 41488 1734 41540
rect 57238 41528 57244 41540
rect 57199 41500 57244 41528
rect 57238 41488 57244 41500
rect 57296 41488 57302 41540
rect 57882 41488 57888 41540
rect 57940 41528 57946 41540
rect 57977 41531 58035 41537
rect 57977 41528 57989 41531
rect 57940 41500 57989 41528
rect 57940 41488 57946 41500
rect 57977 41497 57989 41500
rect 58023 41497 58035 41531
rect 57977 41491 58035 41497
rect 58345 41531 58403 41537
rect 58345 41497 58357 41531
rect 58391 41528 58403 41531
rect 58434 41528 58440 41540
rect 58391 41500 58440 41528
rect 58391 41497 58403 41500
rect 58345 41491 58403 41497
rect 58434 41488 58440 41500
rect 58492 41488 58498 41540
rect 1949 41463 2007 41469
rect 1949 41429 1961 41463
rect 1995 41460 2007 41463
rect 26878 41460 26884 41472
rect 1995 41432 26884 41460
rect 1995 41429 2007 41432
rect 1949 41423 2007 41429
rect 26878 41420 26884 41432
rect 26936 41420 26942 41472
rect 1104 41370 58880 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 58880 41370
rect 1104 41296 58880 41318
rect 1670 41120 1676 41132
rect 1631 41092 1676 41120
rect 1670 41080 1676 41092
rect 1728 41080 1734 41132
rect 1765 40919 1823 40925
rect 1765 40885 1777 40919
rect 1811 40916 1823 40919
rect 21174 40916 21180 40928
rect 1811 40888 21180 40916
rect 1811 40885 1823 40888
rect 1765 40879 1823 40885
rect 21174 40876 21180 40888
rect 21232 40876 21238 40928
rect 1104 40826 58880 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 58880 40826
rect 1104 40752 58880 40774
rect 57514 40468 57520 40520
rect 57572 40508 57578 40520
rect 57885 40511 57943 40517
rect 57885 40508 57897 40511
rect 57572 40480 57897 40508
rect 57572 40468 57578 40480
rect 57885 40477 57897 40480
rect 57931 40477 57943 40511
rect 57885 40471 57943 40477
rect 1670 40440 1676 40452
rect 1631 40412 1676 40440
rect 1670 40400 1676 40412
rect 1728 40400 1734 40452
rect 18598 40400 18604 40452
rect 18656 40440 18662 40452
rect 22462 40440 22468 40452
rect 18656 40412 22468 40440
rect 18656 40400 18662 40412
rect 22462 40400 22468 40412
rect 22520 40400 22526 40452
rect 36630 40400 36636 40452
rect 36688 40440 36694 40452
rect 45094 40440 45100 40452
rect 36688 40412 45100 40440
rect 36688 40400 36694 40412
rect 45094 40400 45100 40412
rect 45152 40400 45158 40452
rect 57054 40440 57060 40452
rect 57015 40412 57060 40440
rect 57054 40400 57060 40412
rect 57112 40400 57118 40452
rect 58161 40443 58219 40449
rect 58161 40440 58173 40443
rect 57900 40412 58173 40440
rect 57900 40384 57928 40412
rect 58161 40409 58173 40412
rect 58207 40409 58219 40443
rect 58161 40403 58219 40409
rect 1765 40375 1823 40381
rect 1765 40341 1777 40375
rect 1811 40372 1823 40375
rect 23290 40372 23296 40384
rect 1811 40344 23296 40372
rect 1811 40341 1823 40344
rect 1765 40335 1823 40341
rect 23290 40332 23296 40344
rect 23348 40332 23354 40384
rect 47578 40332 47584 40384
rect 47636 40372 47642 40384
rect 57149 40375 57207 40381
rect 57149 40372 57161 40375
rect 47636 40344 57161 40372
rect 47636 40332 47642 40344
rect 57149 40341 57161 40344
rect 57195 40341 57207 40375
rect 57149 40335 57207 40341
rect 57882 40332 57888 40384
rect 57940 40332 57946 40384
rect 1104 40282 58880 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 58880 40282
rect 1104 40208 58880 40230
rect 20898 40128 20904 40180
rect 20956 40128 20962 40180
rect 23474 40168 23480 40180
rect 21008 40140 23480 40168
rect 20916 40041 20944 40128
rect 21008 40044 21036 40140
rect 23474 40128 23480 40140
rect 23532 40168 23538 40180
rect 25314 40168 25320 40180
rect 23532 40140 25320 40168
rect 23532 40128 23538 40140
rect 25314 40128 25320 40140
rect 25372 40128 25378 40180
rect 21174 40100 21180 40112
rect 21135 40072 21180 40100
rect 21174 40060 21180 40072
rect 21232 40060 21238 40112
rect 20901 40035 20959 40041
rect 20901 40001 20913 40035
rect 20947 40001 20959 40035
rect 20901 39995 20959 40001
rect 20990 39992 20996 40044
rect 21048 40032 21054 40044
rect 21085 40035 21143 40041
rect 21085 40032 21097 40035
rect 21048 40004 21097 40032
rect 21048 39992 21054 40004
rect 21085 40001 21097 40004
rect 21131 40001 21143 40035
rect 21085 39995 21143 40001
rect 21269 40035 21327 40041
rect 21269 40001 21281 40035
rect 21315 40032 21327 40035
rect 23750 40032 23756 40044
rect 21315 40004 23756 40032
rect 21315 40001 21327 40004
rect 21269 39995 21327 40001
rect 2774 39924 2780 39976
rect 2832 39964 2838 39976
rect 21284 39964 21312 39995
rect 23750 39992 23756 40004
rect 23808 39992 23814 40044
rect 2832 39936 21312 39964
rect 2832 39924 2838 39936
rect 21453 39831 21511 39837
rect 21453 39797 21465 39831
rect 21499 39828 21511 39831
rect 21726 39828 21732 39840
rect 21499 39800 21732 39828
rect 21499 39797 21511 39800
rect 21453 39791 21511 39797
rect 21726 39788 21732 39800
rect 21784 39788 21790 39840
rect 1104 39738 58880 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 58880 39738
rect 1104 39664 58880 39686
rect 2222 39516 2228 39568
rect 2280 39556 2286 39568
rect 2406 39556 2412 39568
rect 2280 39528 2412 39556
rect 2280 39516 2286 39528
rect 2406 39516 2412 39528
rect 2464 39516 2470 39568
rect 2869 39559 2927 39565
rect 2869 39525 2881 39559
rect 2915 39556 2927 39559
rect 22278 39556 22284 39568
rect 2915 39528 22284 39556
rect 2915 39525 2927 39528
rect 2869 39519 2927 39525
rect 22278 39516 22284 39528
rect 22336 39516 22342 39568
rect 1857 39491 1915 39497
rect 1857 39457 1869 39491
rect 1903 39488 1915 39491
rect 1903 39460 2636 39488
rect 1903 39457 1915 39460
rect 1857 39451 1915 39457
rect 2314 39420 2320 39432
rect 2275 39392 2320 39420
rect 2314 39380 2320 39392
rect 2372 39380 2378 39432
rect 2608 39429 2636 39460
rect 2774 39429 2780 39432
rect 2593 39423 2651 39429
rect 2593 39389 2605 39423
rect 2639 39389 2651 39423
rect 2593 39383 2651 39389
rect 2737 39423 2780 39429
rect 2737 39389 2749 39423
rect 2737 39383 2780 39389
rect 2774 39380 2780 39383
rect 2832 39380 2838 39432
rect 1670 39352 1676 39364
rect 1631 39324 1676 39352
rect 1670 39312 1676 39324
rect 1728 39312 1734 39364
rect 2501 39355 2559 39361
rect 2501 39321 2513 39355
rect 2547 39321 2559 39355
rect 2501 39315 2559 39321
rect 2406 39244 2412 39296
rect 2464 39284 2470 39296
rect 2516 39284 2544 39315
rect 13078 39312 13084 39364
rect 13136 39352 13142 39364
rect 23566 39352 23572 39364
rect 13136 39324 23572 39352
rect 13136 39312 13142 39324
rect 23566 39312 23572 39324
rect 23624 39312 23630 39364
rect 57054 39352 57060 39364
rect 57015 39324 57060 39352
rect 57054 39312 57060 39324
rect 57112 39312 57118 39364
rect 57974 39352 57980 39364
rect 57935 39324 57980 39352
rect 57974 39312 57980 39324
rect 58032 39312 58038 39364
rect 2590 39284 2596 39296
rect 2464 39256 2596 39284
rect 2464 39244 2470 39256
rect 2590 39244 2596 39256
rect 2648 39244 2654 39296
rect 33778 39244 33784 39296
rect 33836 39284 33842 39296
rect 57149 39287 57207 39293
rect 57149 39284 57161 39287
rect 33836 39256 57161 39284
rect 33836 39244 33842 39256
rect 57149 39253 57161 39256
rect 57195 39253 57207 39287
rect 58066 39284 58072 39296
rect 58027 39256 58072 39284
rect 57149 39247 57207 39253
rect 58066 39244 58072 39256
rect 58124 39244 58130 39296
rect 1104 39194 58880 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 58880 39194
rect 1104 39120 58880 39142
rect 23124 39052 26234 39080
rect 1670 38944 1676 38956
rect 1631 38916 1676 38944
rect 1670 38904 1676 38916
rect 1728 38904 1734 38956
rect 22922 38944 22928 38956
rect 22883 38916 22928 38944
rect 22922 38904 22928 38916
rect 22980 38904 22986 38956
rect 23124 38953 23152 39052
rect 23290 38972 23296 39024
rect 23348 39012 23354 39024
rect 23348 38984 23390 39012
rect 23348 38972 23354 38984
rect 23073 38947 23152 38953
rect 23073 38913 23085 38947
rect 23119 38916 23152 38947
rect 23119 38913 23131 38916
rect 23073 38907 23131 38913
rect 23198 38904 23204 38956
rect 23256 38944 23262 38956
rect 23390 38947 23448 38953
rect 23256 38916 23301 38944
rect 23256 38904 23262 38916
rect 23390 38913 23402 38947
rect 23436 38913 23448 38947
rect 23390 38907 23448 38913
rect 23400 38876 23428 38907
rect 23124 38848 23428 38876
rect 26206 38876 26234 39052
rect 50706 39040 50712 39092
rect 50764 39080 50770 39092
rect 58066 39080 58072 39092
rect 50764 39052 58072 39080
rect 50764 39040 50770 39052
rect 58066 39040 58072 39052
rect 58124 39040 58130 39092
rect 36998 38876 37004 38888
rect 26206 38848 37004 38876
rect 23124 38820 23152 38848
rect 36998 38836 37004 38848
rect 37056 38836 37062 38888
rect 1854 38808 1860 38820
rect 1815 38780 1860 38808
rect 1854 38768 1860 38780
rect 1912 38768 1918 38820
rect 23106 38768 23112 38820
rect 23164 38768 23170 38820
rect 23569 38743 23627 38749
rect 23569 38709 23581 38743
rect 23615 38740 23627 38743
rect 24762 38740 24768 38752
rect 23615 38712 24768 38740
rect 23615 38709 23627 38712
rect 23569 38703 23627 38709
rect 24762 38700 24768 38712
rect 24820 38700 24826 38752
rect 1104 38650 58880 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 58880 38650
rect 1104 38576 58880 38598
rect 1765 38539 1823 38545
rect 1765 38505 1777 38539
rect 1811 38536 1823 38539
rect 1811 38508 2774 38536
rect 1811 38505 1823 38508
rect 1765 38499 1823 38505
rect 1854 38360 1860 38412
rect 1912 38400 1918 38412
rect 2593 38403 2651 38409
rect 2593 38400 2605 38403
rect 1912 38372 2605 38400
rect 1912 38360 1918 38372
rect 2593 38369 2605 38372
rect 2639 38369 2651 38403
rect 2746 38400 2774 38508
rect 16298 38496 16304 38548
rect 16356 38536 16362 38548
rect 20165 38539 20223 38545
rect 20165 38536 20177 38539
rect 16356 38508 20177 38536
rect 16356 38496 16362 38508
rect 20165 38505 20177 38508
rect 20211 38505 20223 38539
rect 23014 38536 23020 38548
rect 20165 38499 20223 38505
rect 22066 38508 23020 38536
rect 19150 38428 19156 38480
rect 19208 38468 19214 38480
rect 22066 38468 22094 38508
rect 23014 38496 23020 38508
rect 23072 38496 23078 38548
rect 19208 38440 22094 38468
rect 19208 38428 19214 38440
rect 19426 38400 19432 38412
rect 2746 38372 19432 38400
rect 2593 38363 2651 38369
rect 19426 38360 19432 38372
rect 19484 38360 19490 38412
rect 19978 38360 19984 38412
rect 20036 38400 20042 38412
rect 20622 38400 20628 38412
rect 20036 38372 20628 38400
rect 20036 38360 20042 38372
rect 20622 38360 20628 38372
rect 20680 38360 20686 38412
rect 21177 38403 21235 38409
rect 21177 38369 21189 38403
rect 21223 38400 21235 38403
rect 21545 38403 21603 38409
rect 21545 38400 21557 38403
rect 21223 38372 21557 38400
rect 21223 38369 21235 38372
rect 21177 38363 21235 38369
rect 21545 38369 21557 38372
rect 21591 38400 21603 38403
rect 39574 38400 39580 38412
rect 21591 38372 39580 38400
rect 21591 38369 21603 38372
rect 21545 38363 21603 38369
rect 39574 38360 39580 38372
rect 39632 38360 39638 38412
rect 2774 38292 2780 38344
rect 2832 38332 2838 38344
rect 20162 38332 20168 38344
rect 2832 38304 2877 38332
rect 20123 38304 20168 38332
rect 2832 38292 2838 38304
rect 20162 38292 20168 38304
rect 20220 38292 20226 38344
rect 20349 38335 20407 38341
rect 20349 38301 20361 38335
rect 20395 38301 20407 38335
rect 20349 38295 20407 38301
rect 20441 38335 20499 38341
rect 20441 38301 20453 38335
rect 20487 38301 20499 38335
rect 20441 38295 20499 38301
rect 1670 38264 1676 38276
rect 1631 38236 1676 38264
rect 1670 38224 1676 38236
rect 1728 38224 1734 38276
rect 2961 38267 3019 38273
rect 2961 38233 2973 38267
rect 3007 38264 3019 38267
rect 20364 38264 20392 38295
rect 3007 38236 20392 38264
rect 3007 38233 3019 38236
rect 2961 38227 3019 38233
rect 20162 38156 20168 38208
rect 20220 38196 20226 38208
rect 20456 38196 20484 38295
rect 20530 38292 20536 38344
rect 20588 38332 20594 38344
rect 21453 38335 21511 38341
rect 21453 38332 21465 38335
rect 20588 38304 21465 38332
rect 20588 38292 20594 38304
rect 21453 38301 21465 38304
rect 21499 38301 21511 38335
rect 21726 38332 21732 38344
rect 21687 38304 21732 38332
rect 21453 38295 21511 38301
rect 21726 38292 21732 38304
rect 21784 38292 21790 38344
rect 22922 38292 22928 38344
rect 22980 38332 22986 38344
rect 23109 38335 23167 38341
rect 23109 38332 23121 38335
rect 22980 38304 23121 38332
rect 22980 38292 22986 38304
rect 23109 38301 23121 38304
rect 23155 38301 23167 38335
rect 23109 38295 23167 38301
rect 46842 38292 46848 38344
rect 46900 38332 46906 38344
rect 57885 38335 57943 38341
rect 57885 38332 57897 38335
rect 46900 38304 57897 38332
rect 46900 38292 46906 38304
rect 57885 38301 57897 38304
rect 57931 38301 57943 38335
rect 57885 38295 57943 38301
rect 21082 38224 21088 38276
rect 21140 38264 21146 38276
rect 23477 38267 23535 38273
rect 23477 38264 23489 38267
rect 21140 38236 23489 38264
rect 21140 38224 21146 38236
rect 23477 38233 23489 38236
rect 23523 38233 23535 38267
rect 58158 38264 58164 38276
rect 58119 38236 58164 38264
rect 23477 38227 23535 38233
rect 58158 38224 58164 38236
rect 58216 38224 58222 38276
rect 20220 38168 20484 38196
rect 20625 38199 20683 38205
rect 20220 38156 20226 38168
rect 20625 38165 20637 38199
rect 20671 38196 20683 38199
rect 21818 38196 21824 38208
rect 20671 38168 21824 38196
rect 20671 38165 20683 38168
rect 20625 38159 20683 38165
rect 21818 38156 21824 38168
rect 21876 38156 21882 38208
rect 21913 38199 21971 38205
rect 21913 38165 21925 38199
rect 21959 38196 21971 38199
rect 22002 38196 22008 38208
rect 21959 38168 22008 38196
rect 21959 38165 21971 38168
rect 21913 38159 21971 38165
rect 22002 38156 22008 38168
rect 22060 38156 22066 38208
rect 23014 38156 23020 38208
rect 23072 38196 23078 38208
rect 26142 38196 26148 38208
rect 23072 38168 26148 38196
rect 23072 38156 23078 38168
rect 26142 38156 26148 38168
rect 26200 38156 26206 38208
rect 1104 38106 58880 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 58880 38106
rect 1104 38032 58880 38054
rect 5902 37952 5908 38004
rect 5960 37992 5966 38004
rect 5960 37964 22784 37992
rect 5960 37952 5966 37964
rect 2225 37927 2283 37933
rect 2225 37893 2237 37927
rect 2271 37924 2283 37927
rect 2866 37924 2872 37936
rect 2271 37896 2872 37924
rect 2271 37893 2283 37896
rect 2225 37887 2283 37893
rect 2866 37884 2872 37896
rect 2924 37884 2930 37936
rect 6178 37884 6184 37936
rect 6236 37924 6242 37936
rect 20993 37927 21051 37933
rect 20993 37924 21005 37927
rect 6236 37896 21005 37924
rect 6236 37884 6242 37896
rect 20993 37893 21005 37896
rect 21039 37893 21051 37927
rect 20993 37887 21051 37893
rect 1946 37816 1952 37868
rect 2004 37856 2010 37868
rect 2041 37859 2099 37865
rect 2041 37856 2053 37859
rect 2004 37828 2053 37856
rect 2004 37816 2010 37828
rect 2041 37825 2053 37828
rect 2087 37825 2099 37859
rect 2317 37859 2375 37865
rect 2317 37856 2329 37859
rect 2041 37819 2099 37825
rect 2148 37828 2329 37856
rect 2148 37720 2176 37828
rect 2317 37825 2329 37828
rect 2363 37825 2375 37859
rect 2317 37819 2375 37825
rect 2409 37859 2467 37865
rect 2409 37825 2421 37859
rect 2455 37856 2467 37859
rect 3050 37856 3056 37868
rect 2455 37828 3056 37856
rect 2455 37825 2467 37828
rect 2409 37819 2467 37825
rect 2222 37748 2228 37800
rect 2280 37788 2286 37800
rect 2424 37788 2452 37819
rect 3050 37816 3056 37828
rect 3108 37816 3114 37868
rect 19334 37856 19340 37868
rect 19295 37828 19340 37856
rect 19334 37816 19340 37828
rect 19392 37816 19398 37868
rect 19485 37859 19543 37865
rect 19485 37825 19497 37859
rect 19531 37856 19543 37859
rect 19613 37859 19671 37865
rect 19531 37825 19564 37856
rect 19485 37819 19564 37825
rect 19613 37825 19625 37859
rect 19659 37825 19671 37859
rect 19613 37819 19671 37825
rect 2280 37760 2452 37788
rect 2280 37748 2286 37760
rect 2314 37720 2320 37732
rect 2148 37692 2320 37720
rect 2314 37680 2320 37692
rect 2372 37680 2378 37732
rect 2590 37652 2596 37664
rect 2551 37624 2596 37652
rect 2590 37612 2596 37624
rect 2648 37612 2654 37664
rect 19536 37652 19564 37819
rect 19628 37788 19656 37819
rect 19702 37816 19708 37868
rect 19760 37856 19766 37868
rect 19843 37859 19901 37865
rect 19760 37828 19805 37856
rect 19760 37816 19766 37828
rect 19843 37825 19855 37859
rect 19889 37856 19901 37859
rect 20254 37856 20260 37868
rect 19889 37828 20260 37856
rect 19889 37825 19901 37828
rect 19843 37819 19901 37825
rect 20254 37816 20260 37828
rect 20312 37816 20318 37868
rect 20349 37859 20407 37865
rect 20349 37825 20361 37859
rect 20395 37856 20407 37859
rect 20806 37856 20812 37868
rect 20395 37828 20812 37856
rect 20395 37825 20407 37828
rect 20349 37819 20407 37825
rect 20806 37816 20812 37828
rect 20864 37816 20870 37868
rect 20898 37816 20904 37868
rect 20956 37856 20962 37868
rect 21082 37856 21088 37868
rect 20956 37828 21088 37856
rect 20956 37816 20962 37828
rect 21082 37816 21088 37828
rect 21140 37816 21146 37868
rect 22756 37865 22784 37964
rect 23014 37952 23020 38004
rect 23072 37992 23078 38004
rect 23293 37995 23351 38001
rect 23072 37964 23152 37992
rect 23072 37952 23078 37964
rect 22922 37924 22928 37936
rect 22883 37896 22928 37924
rect 22922 37884 22928 37896
rect 22980 37884 22986 37936
rect 22741 37859 22799 37865
rect 22741 37825 22753 37859
rect 22787 37825 22799 37859
rect 23014 37856 23020 37868
rect 22975 37828 23020 37856
rect 22741 37819 22799 37825
rect 23014 37816 23020 37828
rect 23072 37816 23078 37868
rect 23124 37865 23152 37964
rect 23293 37961 23305 37995
rect 23339 37992 23351 37995
rect 23339 37964 23796 37992
rect 23339 37961 23351 37964
rect 23293 37955 23351 37961
rect 23768 37933 23796 37964
rect 25102 37964 25452 37992
rect 23753 37927 23811 37933
rect 23753 37893 23765 37927
rect 23799 37893 23811 37927
rect 25102 37924 25130 37964
rect 25222 37924 25228 37936
rect 23753 37887 23811 37893
rect 23860 37896 25130 37924
rect 25183 37896 25228 37924
rect 23109 37859 23167 37865
rect 23109 37825 23121 37859
rect 23155 37825 23167 37859
rect 23109 37819 23167 37825
rect 22465 37791 22523 37797
rect 19628 37760 21312 37788
rect 21284 37732 21312 37760
rect 22465 37757 22477 37791
rect 22511 37788 22523 37791
rect 22554 37788 22560 37800
rect 22511 37760 22560 37788
rect 22511 37757 22523 37760
rect 22465 37751 22523 37757
rect 22554 37748 22560 37760
rect 22612 37748 22618 37800
rect 19981 37723 20039 37729
rect 19981 37689 19993 37723
rect 20027 37720 20039 37723
rect 20438 37720 20444 37732
rect 20027 37692 20444 37720
rect 20027 37689 20039 37692
rect 19981 37683 20039 37689
rect 20438 37680 20444 37692
rect 20496 37680 20502 37732
rect 21266 37680 21272 37732
rect 21324 37720 21330 37732
rect 23860 37720 23888 37896
rect 25102 37865 25130 37896
rect 25222 37884 25228 37896
rect 25280 37884 25286 37936
rect 24949 37859 25007 37865
rect 24949 37825 24961 37859
rect 24995 37825 25007 37859
rect 24949 37819 25007 37825
rect 25087 37859 25145 37865
rect 25087 37825 25099 37859
rect 25133 37825 25145 37859
rect 25314 37856 25320 37868
rect 25275 37828 25320 37856
rect 25087 37819 25145 37825
rect 23934 37748 23940 37800
rect 23992 37748 23998 37800
rect 24118 37788 24124 37800
rect 24079 37760 24124 37788
rect 24118 37748 24124 37760
rect 24176 37748 24182 37800
rect 24964 37788 24992 37819
rect 25314 37816 25320 37828
rect 25372 37816 25378 37868
rect 25424 37856 25452 37964
rect 26142 37952 26148 38004
rect 26200 37992 26206 38004
rect 26200 37952 26234 37992
rect 26206 37924 26234 37952
rect 37458 37924 37464 37936
rect 26206 37896 37464 37924
rect 37458 37884 37464 37896
rect 37516 37884 37522 37936
rect 29730 37856 29736 37868
rect 25424 37828 29736 37856
rect 29730 37816 29736 37828
rect 29788 37816 29794 37868
rect 58066 37856 58072 37868
rect 58027 37828 58072 37856
rect 58066 37816 58072 37828
rect 58124 37816 58130 37868
rect 44174 37788 44180 37800
rect 24964 37760 44180 37788
rect 44174 37748 44180 37760
rect 44232 37748 44238 37800
rect 21324 37692 23888 37720
rect 23952 37720 23980 37748
rect 24029 37723 24087 37729
rect 24029 37720 24041 37723
rect 23952 37692 24041 37720
rect 21324 37680 21330 37692
rect 24029 37689 24041 37692
rect 24075 37689 24087 37723
rect 25501 37723 25559 37729
rect 25501 37720 25513 37723
rect 24029 37683 24087 37689
rect 24136 37692 25513 37720
rect 20346 37652 20352 37664
rect 19536 37624 20352 37652
rect 20346 37612 20352 37624
rect 20404 37612 20410 37664
rect 20622 37652 20628 37664
rect 20583 37624 20628 37652
rect 20622 37612 20628 37624
rect 20680 37612 20686 37664
rect 23918 37655 23976 37661
rect 23918 37621 23930 37655
rect 23964 37652 23976 37655
rect 24136 37652 24164 37692
rect 25501 37689 25513 37692
rect 25547 37689 25559 37723
rect 25501 37683 25559 37689
rect 24394 37652 24400 37664
rect 23964 37624 24164 37652
rect 24355 37624 24400 37652
rect 23964 37621 23976 37624
rect 23918 37615 23976 37621
rect 24394 37612 24400 37624
rect 24452 37612 24458 37664
rect 58253 37655 58311 37661
rect 58253 37621 58265 37655
rect 58299 37652 58311 37655
rect 58526 37652 58532 37664
rect 58299 37624 58532 37652
rect 58299 37621 58311 37624
rect 58253 37615 58311 37621
rect 58526 37612 58532 37624
rect 58584 37612 58590 37664
rect 1104 37562 58880 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 58880 37562
rect 1104 37488 58880 37510
rect 2590 37408 2596 37460
rect 2648 37448 2654 37460
rect 16298 37448 16304 37460
rect 2648 37420 16304 37448
rect 2648 37408 2654 37420
rect 16298 37408 16304 37420
rect 16356 37408 16362 37460
rect 16482 37408 16488 37460
rect 16540 37448 16546 37460
rect 20714 37448 20720 37460
rect 16540 37420 20720 37448
rect 16540 37408 16546 37420
rect 20714 37408 20720 37420
rect 20772 37408 20778 37460
rect 20806 37408 20812 37460
rect 20864 37448 20870 37460
rect 54202 37448 54208 37460
rect 20864 37420 54208 37448
rect 20864 37408 20870 37420
rect 54202 37408 54208 37420
rect 54260 37408 54266 37460
rect 20254 37340 20260 37392
rect 20312 37380 20318 37392
rect 23106 37380 23112 37392
rect 20312 37352 23112 37380
rect 20312 37340 20318 37352
rect 23106 37340 23112 37352
rect 23164 37340 23170 37392
rect 1857 37315 1915 37321
rect 1857 37281 1869 37315
rect 1903 37312 1915 37315
rect 2682 37312 2688 37324
rect 1903 37284 2688 37312
rect 1903 37281 1915 37284
rect 1857 37275 1915 37281
rect 2682 37272 2688 37284
rect 2740 37272 2746 37324
rect 3050 37272 3056 37324
rect 3108 37312 3114 37324
rect 9030 37312 9036 37324
rect 3108 37284 9036 37312
rect 3108 37272 3114 37284
rect 1670 37244 1676 37256
rect 1631 37216 1676 37244
rect 1670 37204 1676 37216
rect 1728 37204 1734 37256
rect 5905 37247 5963 37253
rect 5905 37244 5917 37247
rect 5736 37216 5917 37244
rect 5534 37108 5540 37120
rect 5495 37080 5540 37108
rect 5534 37068 5540 37080
rect 5592 37068 5598 37120
rect 5736 37108 5764 37216
rect 5905 37213 5917 37216
rect 5951 37213 5963 37247
rect 5905 37207 5963 37213
rect 5994 37204 6000 37256
rect 6052 37244 6058 37256
rect 6270 37244 6276 37256
rect 6052 37216 6097 37244
rect 6231 37216 6276 37244
rect 6052 37204 6058 37216
rect 6270 37204 6276 37216
rect 6328 37204 6334 37256
rect 6564 37253 6592 37284
rect 9030 37272 9036 37284
rect 9088 37272 9094 37324
rect 21082 37312 21088 37324
rect 21043 37284 21088 37312
rect 21082 37272 21088 37284
rect 21140 37272 21146 37324
rect 6549 37247 6607 37253
rect 6549 37213 6561 37247
rect 6595 37213 6607 37247
rect 6730 37244 6736 37256
rect 6691 37216 6736 37244
rect 6549 37207 6607 37213
rect 6730 37204 6736 37216
rect 6788 37204 6794 37256
rect 19334 37244 19340 37256
rect 9646 37216 19340 37244
rect 9646 37176 9674 37216
rect 19334 37204 19340 37216
rect 19392 37204 19398 37256
rect 19613 37247 19671 37253
rect 19613 37213 19625 37247
rect 19659 37244 19671 37247
rect 20530 37244 20536 37256
rect 19659 37216 20536 37244
rect 19659 37213 19671 37216
rect 19613 37207 19671 37213
rect 20530 37204 20536 37216
rect 20588 37204 20594 37256
rect 20901 37247 20959 37253
rect 20901 37213 20913 37247
rect 20947 37244 20959 37247
rect 21910 37244 21916 37256
rect 20947 37216 21916 37244
rect 20947 37213 20959 37216
rect 20901 37207 20959 37213
rect 21910 37204 21916 37216
rect 21968 37204 21974 37256
rect 53834 37244 53840 37256
rect 53795 37216 53840 37244
rect 53834 37204 53840 37216
rect 53892 37204 53898 37256
rect 54110 37244 54116 37256
rect 54071 37216 54116 37244
rect 54110 37204 54116 37216
rect 54168 37204 54174 37256
rect 54294 37253 54300 37256
rect 54257 37247 54300 37253
rect 54257 37213 54269 37247
rect 54257 37207 54300 37213
rect 54294 37204 54300 37207
rect 54352 37204 54358 37256
rect 54478 37204 54484 37256
rect 54536 37244 54542 37256
rect 57885 37247 57943 37253
rect 57885 37244 57897 37247
rect 54536 37216 57897 37244
rect 54536 37204 54542 37216
rect 57885 37213 57897 37216
rect 57931 37213 57943 37247
rect 57885 37207 57943 37213
rect 8956 37148 9674 37176
rect 8956 37108 8984 37148
rect 18782 37136 18788 37188
rect 18840 37176 18846 37188
rect 19981 37179 20039 37185
rect 19981 37176 19993 37179
rect 18840 37148 19993 37176
rect 18840 37136 18846 37148
rect 19981 37145 19993 37148
rect 20027 37176 20039 37179
rect 20990 37176 20996 37188
rect 20027 37148 20996 37176
rect 20027 37145 20039 37148
rect 19981 37139 20039 37145
rect 20990 37136 20996 37148
rect 21048 37136 21054 37188
rect 54018 37176 54024 37188
rect 53979 37148 54024 37176
rect 54018 37136 54024 37148
rect 54076 37136 54082 37188
rect 58158 37176 58164 37188
rect 58119 37148 58164 37176
rect 58158 37136 58164 37148
rect 58216 37136 58222 37188
rect 5736 37080 8984 37108
rect 9030 37068 9036 37120
rect 9088 37108 9094 37120
rect 19242 37108 19248 37120
rect 9088 37080 19248 37108
rect 9088 37068 9094 37080
rect 19242 37068 19248 37080
rect 19300 37068 19306 37120
rect 49970 37068 49976 37120
rect 50028 37108 50034 37120
rect 54397 37111 54455 37117
rect 54397 37108 54409 37111
rect 50028 37080 54409 37108
rect 50028 37068 50034 37080
rect 54397 37077 54409 37080
rect 54443 37077 54455 37111
rect 54397 37071 54455 37077
rect 1104 37018 58880 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 58880 37018
rect 1104 36944 58880 36966
rect 5994 36864 6000 36916
rect 6052 36904 6058 36916
rect 42886 36904 42892 36916
rect 6052 36876 42892 36904
rect 6052 36864 6058 36876
rect 42886 36864 42892 36876
rect 42944 36864 42950 36916
rect 45526 36876 54064 36904
rect 18693 36839 18751 36845
rect 18693 36805 18705 36839
rect 18739 36836 18751 36839
rect 18874 36836 18880 36848
rect 18739 36808 18880 36836
rect 18739 36805 18751 36808
rect 18693 36799 18751 36805
rect 18874 36796 18880 36808
rect 18932 36796 18938 36848
rect 20070 36796 20076 36848
rect 20128 36836 20134 36848
rect 20254 36836 20260 36848
rect 20128 36808 20260 36836
rect 20128 36796 20134 36808
rect 20254 36796 20260 36808
rect 20312 36796 20318 36848
rect 20530 36796 20536 36848
rect 20588 36836 20594 36848
rect 28442 36836 28448 36848
rect 20588 36808 28448 36836
rect 20588 36796 20594 36808
rect 28442 36796 28448 36808
rect 28500 36796 28506 36848
rect 36262 36796 36268 36848
rect 36320 36836 36326 36848
rect 45526 36836 45554 36876
rect 53926 36836 53932 36848
rect 36320 36808 45554 36836
rect 53887 36808 53932 36836
rect 36320 36796 36326 36808
rect 53926 36796 53932 36808
rect 53984 36796 53990 36848
rect 1578 36768 1584 36780
rect 1539 36740 1584 36768
rect 1578 36728 1584 36740
rect 1636 36728 1642 36780
rect 18414 36768 18420 36780
rect 18375 36740 18420 36768
rect 18414 36728 18420 36740
rect 18472 36728 18478 36780
rect 18601 36771 18659 36777
rect 18601 36737 18613 36771
rect 18647 36737 18659 36771
rect 18782 36768 18788 36780
rect 18743 36740 18788 36768
rect 18601 36731 18659 36737
rect 18616 36700 18644 36731
rect 18782 36728 18788 36740
rect 18840 36728 18846 36780
rect 19426 36768 19432 36780
rect 19387 36740 19432 36768
rect 19426 36728 19432 36740
rect 19484 36728 19490 36780
rect 20990 36768 20996 36780
rect 20088 36740 20996 36768
rect 20088 36700 20116 36740
rect 20990 36728 20996 36740
rect 21048 36728 21054 36780
rect 23477 36771 23535 36777
rect 23477 36737 23489 36771
rect 23523 36768 23535 36771
rect 23753 36771 23811 36777
rect 23753 36768 23765 36771
rect 23523 36740 23765 36768
rect 23523 36737 23535 36740
rect 23477 36731 23535 36737
rect 23753 36737 23765 36740
rect 23799 36768 23811 36771
rect 23799 36740 23980 36768
rect 23799 36737 23811 36740
rect 23753 36731 23811 36737
rect 18616 36672 20116 36700
rect 20162 36660 20168 36712
rect 20220 36700 20226 36712
rect 23842 36700 23848 36712
rect 20220 36672 23336 36700
rect 23803 36672 23848 36700
rect 20220 36660 20226 36672
rect 19334 36592 19340 36644
rect 19392 36632 19398 36644
rect 20717 36635 20775 36641
rect 20717 36632 20729 36635
rect 19392 36604 20729 36632
rect 19392 36592 19398 36604
rect 20717 36601 20729 36604
rect 20763 36601 20775 36635
rect 23308 36632 23336 36672
rect 23842 36660 23848 36672
rect 23900 36660 23906 36712
rect 23952 36700 23980 36740
rect 24026 36728 24032 36780
rect 24084 36768 24090 36780
rect 25498 36768 25504 36780
rect 24084 36740 25504 36768
rect 24084 36728 24090 36740
rect 25498 36728 25504 36740
rect 25556 36728 25562 36780
rect 53650 36768 53656 36780
rect 53611 36740 53656 36768
rect 53650 36728 53656 36740
rect 53708 36728 53714 36780
rect 54036 36777 54064 36876
rect 53837 36771 53895 36777
rect 53837 36737 53849 36771
rect 53883 36737 53895 36771
rect 53837 36731 53895 36737
rect 54026 36771 54084 36777
rect 54026 36737 54038 36771
rect 54072 36737 54084 36771
rect 54026 36731 54084 36737
rect 37274 36700 37280 36712
rect 23952 36672 37280 36700
rect 37274 36660 37280 36672
rect 37332 36660 37338 36712
rect 53852 36700 53880 36731
rect 53852 36672 54064 36700
rect 54036 36644 54064 36672
rect 49970 36632 49976 36644
rect 23308 36604 49976 36632
rect 20717 36595 20775 36601
rect 49970 36592 49976 36604
rect 50028 36592 50034 36644
rect 54018 36592 54024 36644
rect 54076 36592 54082 36644
rect 54202 36632 54208 36644
rect 54163 36604 54208 36632
rect 54202 36592 54208 36604
rect 54260 36592 54266 36644
rect 1765 36567 1823 36573
rect 1765 36533 1777 36567
rect 1811 36564 1823 36567
rect 2590 36564 2596 36576
rect 1811 36536 2596 36564
rect 1811 36533 1823 36536
rect 1765 36527 1823 36533
rect 2590 36524 2596 36536
rect 2648 36524 2654 36576
rect 18969 36567 19027 36573
rect 18969 36533 18981 36567
rect 19015 36564 19027 36567
rect 20070 36564 20076 36576
rect 19015 36536 20076 36564
rect 19015 36533 19027 36536
rect 18969 36527 19027 36533
rect 20070 36524 20076 36536
rect 20128 36524 20134 36576
rect 23474 36524 23480 36576
rect 23532 36564 23538 36576
rect 23753 36567 23811 36573
rect 23753 36564 23765 36567
rect 23532 36536 23765 36564
rect 23532 36524 23538 36536
rect 23753 36533 23765 36536
rect 23799 36533 23811 36567
rect 23753 36527 23811 36533
rect 24213 36567 24271 36573
rect 24213 36533 24225 36567
rect 24259 36564 24271 36567
rect 24578 36564 24584 36576
rect 24259 36536 24584 36564
rect 24259 36533 24271 36536
rect 24213 36527 24271 36533
rect 24578 36524 24584 36536
rect 24636 36524 24642 36576
rect 53834 36524 53840 36576
rect 53892 36564 53898 36576
rect 55030 36564 55036 36576
rect 53892 36536 55036 36564
rect 53892 36524 53898 36536
rect 55030 36524 55036 36536
rect 55088 36524 55094 36576
rect 1104 36474 58880 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 58880 36474
rect 1104 36400 58880 36422
rect 1765 36363 1823 36369
rect 1765 36329 1777 36363
rect 1811 36360 1823 36363
rect 3053 36363 3111 36369
rect 1811 36332 2774 36360
rect 1811 36329 1823 36332
rect 1765 36323 1823 36329
rect 2746 36292 2774 36332
rect 3053 36329 3065 36363
rect 3099 36360 3111 36363
rect 23474 36360 23480 36372
rect 3099 36332 23480 36360
rect 3099 36329 3111 36332
rect 3053 36323 3111 36329
rect 23474 36320 23480 36332
rect 23532 36320 23538 36372
rect 23842 36360 23848 36372
rect 23803 36332 23848 36360
rect 23842 36320 23848 36332
rect 23900 36320 23906 36372
rect 6730 36292 6736 36304
rect 2746 36264 6736 36292
rect 6730 36252 6736 36264
rect 6788 36252 6794 36304
rect 20257 36295 20315 36301
rect 20257 36261 20269 36295
rect 20303 36292 20315 36295
rect 20622 36292 20628 36304
rect 20303 36264 20628 36292
rect 20303 36261 20315 36264
rect 20257 36255 20315 36261
rect 20622 36252 20628 36264
rect 20680 36252 20686 36304
rect 20990 36252 20996 36304
rect 21048 36292 21054 36304
rect 23198 36292 23204 36304
rect 21048 36264 23204 36292
rect 21048 36252 21054 36264
rect 23198 36252 23204 36264
rect 23256 36252 23262 36304
rect 20714 36224 20720 36236
rect 20675 36196 20720 36224
rect 20714 36184 20720 36196
rect 20772 36184 20778 36236
rect 33226 36224 33232 36236
rect 22572 36196 23428 36224
rect 2498 36156 2504 36168
rect 2459 36128 2504 36156
rect 2498 36116 2504 36128
rect 2556 36116 2562 36168
rect 2866 36116 2872 36168
rect 2924 36165 2930 36168
rect 2924 36156 2932 36165
rect 3050 36156 3056 36168
rect 2924 36128 3056 36156
rect 2924 36119 2932 36128
rect 2924 36116 2930 36119
rect 3050 36116 3056 36128
rect 3108 36116 3114 36168
rect 20162 36156 20168 36168
rect 20123 36128 20168 36156
rect 20162 36116 20168 36128
rect 20220 36116 20226 36168
rect 20438 36156 20444 36168
rect 20399 36128 20444 36156
rect 20438 36116 20444 36128
rect 20496 36116 20502 36168
rect 22186 36156 22192 36168
rect 22147 36128 22192 36156
rect 22186 36116 22192 36128
rect 22244 36116 22250 36168
rect 22462 36156 22468 36168
rect 22423 36128 22468 36156
rect 22462 36116 22468 36128
rect 22520 36116 22526 36168
rect 22572 36165 22600 36196
rect 23400 36168 23428 36196
rect 23676 36196 33232 36224
rect 22557 36159 22615 36165
rect 22557 36125 22569 36159
rect 22603 36125 22615 36159
rect 23290 36156 23296 36168
rect 23251 36128 23296 36156
rect 22557 36119 22615 36125
rect 23290 36116 23296 36128
rect 23348 36116 23354 36168
rect 23382 36116 23388 36168
rect 23440 36156 23446 36168
rect 23676 36165 23704 36196
rect 33226 36184 33232 36196
rect 33284 36184 33290 36236
rect 23661 36159 23719 36165
rect 23661 36156 23673 36159
rect 23440 36128 23673 36156
rect 23440 36116 23446 36128
rect 23661 36125 23673 36128
rect 23707 36125 23719 36159
rect 24578 36156 24584 36168
rect 24539 36128 24584 36156
rect 23661 36119 23719 36125
rect 24578 36116 24584 36128
rect 24636 36116 24642 36168
rect 24762 36156 24768 36168
rect 24723 36128 24768 36156
rect 24762 36116 24768 36128
rect 24820 36116 24826 36168
rect 1670 36088 1676 36100
rect 1631 36060 1676 36088
rect 1670 36048 1676 36060
rect 1728 36048 1734 36100
rect 2406 36048 2412 36100
rect 2464 36088 2470 36100
rect 2685 36091 2743 36097
rect 2685 36088 2697 36091
rect 2464 36060 2697 36088
rect 2464 36048 2470 36060
rect 2685 36057 2697 36060
rect 2731 36057 2743 36091
rect 2685 36051 2743 36057
rect 2700 36020 2728 36051
rect 2774 36048 2780 36100
rect 2832 36088 2838 36100
rect 22373 36091 22431 36097
rect 2832 36060 2877 36088
rect 2832 36048 2838 36060
rect 22373 36057 22385 36091
rect 22419 36057 22431 36091
rect 23477 36091 23535 36097
rect 23477 36088 23489 36091
rect 22373 36051 22431 36057
rect 22572 36060 23489 36088
rect 15746 36020 15752 36032
rect 2700 35992 15752 36020
rect 15746 35980 15752 35992
rect 15804 36020 15810 36032
rect 16482 36020 16488 36032
rect 15804 35992 16488 36020
rect 15804 35980 15810 35992
rect 16482 35980 16488 35992
rect 16540 35980 16546 36032
rect 22388 36020 22416 36051
rect 22572 36020 22600 36060
rect 23477 36057 23489 36060
rect 23523 36057 23535 36091
rect 23477 36051 23535 36057
rect 22738 36020 22744 36032
rect 22388 35992 22600 36020
rect 22699 35992 22744 36020
rect 22738 35980 22744 35992
rect 22796 35980 22802 36032
rect 23492 36020 23520 36051
rect 23566 36048 23572 36100
rect 23624 36088 23630 36100
rect 25133 36091 25191 36097
rect 23624 36060 23669 36088
rect 23624 36048 23630 36060
rect 25133 36057 25145 36091
rect 25179 36088 25191 36091
rect 25406 36088 25412 36100
rect 25179 36060 25412 36088
rect 25179 36057 25191 36060
rect 25133 36051 25191 36057
rect 25406 36048 25412 36060
rect 25464 36048 25470 36100
rect 57974 36088 57980 36100
rect 57935 36060 57980 36088
rect 57974 36048 57980 36060
rect 58032 36048 58038 36100
rect 58345 36091 58403 36097
rect 58345 36057 58357 36091
rect 58391 36088 58403 36091
rect 58894 36088 58900 36100
rect 58391 36060 58900 36088
rect 58391 36057 58403 36060
rect 58345 36051 58403 36057
rect 58894 36048 58900 36060
rect 58952 36048 58958 36100
rect 24946 36020 24952 36032
rect 23492 35992 24952 36020
rect 24946 35980 24952 35992
rect 25004 35980 25010 36032
rect 1104 35930 58880 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 58880 35930
rect 1104 35856 58880 35878
rect 1762 35816 1768 35828
rect 1723 35788 1768 35816
rect 1762 35776 1768 35788
rect 1820 35776 1826 35828
rect 19334 35776 19340 35828
rect 19392 35816 19398 35828
rect 19392 35788 19564 35816
rect 19392 35776 19398 35788
rect 19242 35748 19248 35760
rect 19203 35720 19248 35748
rect 19242 35708 19248 35720
rect 19300 35708 19306 35760
rect 19536 35748 19564 35788
rect 20162 35776 20168 35828
rect 20220 35816 20226 35828
rect 20441 35819 20499 35825
rect 20441 35816 20453 35819
rect 20220 35788 20453 35816
rect 20220 35776 20226 35788
rect 20441 35785 20453 35788
rect 20487 35785 20499 35819
rect 33042 35816 33048 35828
rect 20441 35779 20499 35785
rect 24688 35788 33048 35816
rect 24688 35760 24716 35788
rect 33042 35776 33048 35788
rect 33100 35776 33106 35828
rect 37274 35776 37280 35828
rect 37332 35816 37338 35828
rect 40773 35819 40831 35825
rect 40773 35816 40785 35819
rect 37332 35788 40785 35816
rect 37332 35776 37338 35788
rect 40773 35785 40785 35788
rect 40819 35785 40831 35819
rect 40773 35779 40831 35785
rect 24670 35748 24676 35760
rect 19536 35720 24676 35748
rect 1670 35680 1676 35692
rect 1631 35652 1676 35680
rect 1670 35640 1676 35652
rect 1728 35640 1734 35692
rect 16574 35640 16580 35692
rect 16632 35680 16638 35692
rect 19061 35683 19119 35689
rect 19061 35680 19073 35683
rect 16632 35652 19073 35680
rect 16632 35640 16638 35652
rect 19061 35649 19073 35652
rect 19107 35649 19119 35683
rect 19061 35643 19119 35649
rect 19337 35683 19395 35689
rect 19337 35649 19349 35683
rect 19383 35649 19395 35683
rect 19337 35643 19395 35649
rect 19429 35683 19487 35689
rect 19429 35649 19441 35683
rect 19475 35680 19487 35683
rect 19536 35680 19564 35720
rect 24670 35708 24676 35720
rect 24728 35708 24734 35760
rect 29730 35708 29736 35760
rect 29788 35748 29794 35760
rect 40405 35751 40463 35757
rect 40405 35748 40417 35751
rect 29788 35720 40417 35748
rect 29788 35708 29794 35720
rect 40405 35717 40417 35720
rect 40451 35717 40463 35751
rect 40405 35711 40463 35717
rect 40512 35720 41414 35748
rect 20073 35683 20131 35689
rect 20073 35680 20085 35683
rect 19475 35652 19564 35680
rect 19628 35652 20085 35680
rect 19475 35649 19487 35652
rect 19429 35643 19487 35649
rect 19352 35556 19380 35643
rect 19334 35504 19340 35556
rect 19392 35504 19398 35556
rect 19628 35553 19656 35652
rect 20073 35649 20085 35652
rect 20119 35649 20131 35683
rect 20073 35643 20131 35649
rect 21082 35640 21088 35692
rect 21140 35680 21146 35692
rect 22649 35683 22707 35689
rect 22649 35680 22661 35683
rect 21140 35652 22661 35680
rect 21140 35640 21146 35652
rect 22649 35649 22661 35652
rect 22695 35649 22707 35683
rect 24118 35680 24124 35692
rect 22649 35643 22707 35649
rect 22756 35652 24124 35680
rect 20165 35615 20223 35621
rect 20165 35581 20177 35615
rect 20211 35612 20223 35615
rect 22756 35612 22784 35652
rect 24118 35640 24124 35652
rect 24176 35640 24182 35692
rect 40512 35689 40540 35720
rect 40221 35683 40279 35689
rect 40221 35649 40233 35683
rect 40267 35680 40279 35683
rect 40497 35683 40555 35689
rect 40267 35652 40448 35680
rect 40267 35649 40279 35652
rect 40221 35643 40279 35649
rect 40420 35624 40448 35652
rect 40497 35649 40509 35683
rect 40543 35649 40555 35683
rect 40497 35643 40555 35649
rect 40586 35640 40592 35692
rect 40644 35680 40650 35692
rect 40644 35652 40689 35680
rect 40644 35640 40650 35652
rect 23382 35612 23388 35624
rect 20211 35584 22784 35612
rect 23343 35584 23388 35612
rect 20211 35581 20223 35584
rect 20165 35575 20223 35581
rect 23382 35572 23388 35584
rect 23440 35572 23446 35624
rect 40402 35572 40408 35624
rect 40460 35572 40466 35624
rect 41386 35612 41414 35720
rect 41690 35612 41696 35624
rect 40512 35584 40816 35612
rect 41386 35584 41696 35612
rect 19613 35547 19671 35553
rect 19613 35513 19625 35547
rect 19659 35513 19671 35547
rect 19613 35507 19671 35513
rect 22186 35504 22192 35556
rect 22244 35544 22250 35556
rect 40512 35544 40540 35584
rect 22244 35516 40540 35544
rect 22244 35504 22250 35516
rect 40586 35504 40592 35556
rect 40644 35504 40650 35556
rect 40788 35544 40816 35584
rect 41690 35572 41696 35584
rect 41748 35572 41754 35624
rect 48958 35544 48964 35556
rect 40788 35516 48964 35544
rect 48958 35504 48964 35516
rect 49016 35504 49022 35556
rect 20070 35476 20076 35488
rect 20031 35448 20076 35476
rect 20070 35436 20076 35448
rect 20128 35436 20134 35488
rect 33042 35436 33048 35488
rect 33100 35476 33106 35488
rect 40604 35476 40632 35504
rect 33100 35448 40632 35476
rect 33100 35436 33106 35448
rect 1104 35386 58880 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 58880 35386
rect 1104 35312 58880 35334
rect 2682 35232 2688 35284
rect 2740 35272 2746 35284
rect 13814 35272 13820 35284
rect 2740 35244 13820 35272
rect 2740 35232 2746 35244
rect 13814 35232 13820 35244
rect 13872 35232 13878 35284
rect 22738 35272 22744 35284
rect 22699 35244 22744 35272
rect 22738 35232 22744 35244
rect 22796 35232 22802 35284
rect 40589 35275 40647 35281
rect 40589 35272 40601 35275
rect 36096 35244 40601 35272
rect 1857 35207 1915 35213
rect 1857 35173 1869 35207
rect 1903 35204 1915 35207
rect 2774 35204 2780 35216
rect 1903 35176 2780 35204
rect 1903 35173 1915 35176
rect 1857 35167 1915 35173
rect 2774 35164 2780 35176
rect 2832 35164 2838 35216
rect 23290 35164 23296 35216
rect 23348 35204 23354 35216
rect 31754 35204 31760 35216
rect 23348 35176 31760 35204
rect 23348 35164 23354 35176
rect 31754 35164 31760 35176
rect 31812 35164 31818 35216
rect 22741 35139 22799 35145
rect 22741 35105 22753 35139
rect 22787 35136 22799 35139
rect 36096 35136 36124 35244
rect 40589 35241 40601 35244
rect 40635 35241 40647 35275
rect 40589 35235 40647 35241
rect 40678 35232 40684 35284
rect 40736 35272 40742 35284
rect 47670 35272 47676 35284
rect 40736 35244 47676 35272
rect 40736 35232 40742 35244
rect 47670 35232 47676 35244
rect 47728 35232 47734 35284
rect 53190 35204 53196 35216
rect 22787 35108 36124 35136
rect 36280 35176 53196 35204
rect 22787 35105 22799 35108
rect 22741 35099 22799 35105
rect 22278 35028 22284 35080
rect 22336 35068 22342 35080
rect 22557 35071 22615 35077
rect 22557 35068 22569 35071
rect 22336 35040 22569 35068
rect 22336 35028 22342 35040
rect 22557 35037 22569 35040
rect 22603 35037 22615 35071
rect 22557 35031 22615 35037
rect 22833 35071 22891 35077
rect 22833 35037 22845 35071
rect 22879 35068 22891 35071
rect 24854 35068 24860 35080
rect 22879 35040 24860 35068
rect 22879 35037 22891 35040
rect 22833 35031 22891 35037
rect 24854 35028 24860 35040
rect 24912 35028 24918 35080
rect 31754 35028 31760 35080
rect 31812 35068 31818 35080
rect 36280 35068 36308 35176
rect 53190 35164 53196 35176
rect 53248 35164 53254 35216
rect 40494 35136 40500 35148
rect 40052 35108 40500 35136
rect 40052 35077 40080 35108
rect 40494 35096 40500 35108
rect 40552 35096 40558 35148
rect 31812 35040 36308 35068
rect 40037 35071 40095 35077
rect 31812 35028 31818 35040
rect 40037 35037 40049 35071
rect 40083 35037 40095 35071
rect 40310 35068 40316 35080
rect 40271 35040 40316 35068
rect 40037 35031 40095 35037
rect 40310 35028 40316 35040
rect 40368 35028 40374 35080
rect 40402 35028 40408 35080
rect 40460 35068 40466 35080
rect 40460 35040 40505 35068
rect 40460 35028 40466 35040
rect 51626 35028 51632 35080
rect 51684 35068 51690 35080
rect 57885 35071 57943 35077
rect 57885 35068 57897 35071
rect 51684 35040 57897 35068
rect 51684 35028 51690 35040
rect 57885 35037 57897 35040
rect 57931 35037 57943 35071
rect 57885 35031 57943 35037
rect 1670 35000 1676 35012
rect 1631 34972 1676 35000
rect 1670 34960 1676 34972
rect 1728 34960 1734 35012
rect 23198 34960 23204 35012
rect 23256 35000 23262 35012
rect 40221 35003 40279 35009
rect 40221 35000 40233 35003
rect 23256 34972 40233 35000
rect 23256 34960 23262 34972
rect 40221 34969 40233 34972
rect 40267 34969 40279 35003
rect 58158 35000 58164 35012
rect 58119 34972 58164 35000
rect 40221 34963 40279 34969
rect 58158 34960 58164 34972
rect 58216 34960 58222 35012
rect 23014 34932 23020 34944
rect 22975 34904 23020 34932
rect 23014 34892 23020 34904
rect 23072 34892 23078 34944
rect 1104 34842 58880 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 58880 34842
rect 1104 34768 58880 34790
rect 19334 34688 19340 34740
rect 19392 34728 19398 34740
rect 39114 34728 39120 34740
rect 19392 34700 39120 34728
rect 19392 34688 19398 34700
rect 39114 34688 39120 34700
rect 39172 34688 39178 34740
rect 58253 34731 58311 34737
rect 58253 34697 58265 34731
rect 58299 34728 58311 34731
rect 58986 34728 58992 34740
rect 58299 34700 58992 34728
rect 58299 34697 58311 34700
rect 58253 34691 58311 34697
rect 58986 34688 58992 34700
rect 59044 34688 59050 34740
rect 19978 34620 19984 34672
rect 20036 34660 20042 34672
rect 22370 34660 22376 34672
rect 20036 34632 22376 34660
rect 20036 34620 20042 34632
rect 22370 34620 22376 34632
rect 22428 34620 22434 34672
rect 19426 34552 19432 34604
rect 19484 34592 19490 34604
rect 22830 34592 22836 34604
rect 19484 34564 22836 34592
rect 19484 34552 19490 34564
rect 22830 34552 22836 34564
rect 22888 34552 22894 34604
rect 57882 34552 57888 34604
rect 57940 34592 57946 34604
rect 58069 34595 58127 34601
rect 58069 34592 58081 34595
rect 57940 34564 58081 34592
rect 57940 34552 57946 34564
rect 58069 34561 58081 34564
rect 58115 34561 58127 34595
rect 58069 34555 58127 34561
rect 20990 34416 20996 34468
rect 21048 34456 21054 34468
rect 23198 34456 23204 34468
rect 21048 34428 23204 34456
rect 21048 34416 21054 34428
rect 23198 34416 23204 34428
rect 23256 34456 23262 34468
rect 23566 34456 23572 34468
rect 23256 34428 23572 34456
rect 23256 34416 23262 34428
rect 23566 34416 23572 34428
rect 23624 34416 23630 34468
rect 40402 34416 40408 34468
rect 40460 34456 40466 34468
rect 43254 34456 43260 34468
rect 40460 34428 43260 34456
rect 40460 34416 40466 34428
rect 43254 34416 43260 34428
rect 43312 34416 43318 34468
rect 1104 34298 58880 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 58880 34298
rect 1104 34224 58880 34246
rect 21726 34144 21732 34196
rect 21784 34184 21790 34196
rect 21784 34156 21869 34184
rect 21784 34144 21790 34156
rect 17310 34076 17316 34128
rect 17368 34116 17374 34128
rect 21542 34116 21548 34128
rect 17368 34088 21548 34116
rect 17368 34076 17374 34088
rect 21542 34076 21548 34088
rect 21600 34076 21606 34128
rect 21358 33980 21364 33992
rect 21319 33952 21364 33980
rect 21358 33940 21364 33952
rect 21416 33940 21422 33992
rect 21542 33989 21548 33992
rect 21509 33983 21548 33989
rect 21509 33949 21521 33983
rect 21509 33943 21548 33949
rect 21542 33940 21548 33943
rect 21600 33940 21606 33992
rect 21841 33989 21869 34156
rect 22186 34076 22192 34128
rect 22244 34116 22250 34128
rect 22244 34088 26234 34116
rect 22244 34076 22250 34088
rect 26206 34048 26234 34088
rect 46290 34048 46296 34060
rect 24964 34020 25544 34048
rect 26206 34020 46296 34048
rect 21826 33983 21884 33989
rect 21826 33949 21838 33983
rect 21872 33949 21884 33983
rect 21826 33943 21884 33949
rect 22557 33983 22615 33989
rect 22557 33949 22569 33983
rect 22603 33949 22615 33983
rect 23014 33980 23020 33992
rect 22975 33952 23020 33980
rect 22557 33943 22615 33949
rect 1670 33912 1676 33924
rect 1631 33884 1676 33912
rect 1670 33872 1676 33884
rect 1728 33872 1734 33924
rect 21266 33872 21272 33924
rect 21324 33912 21330 33924
rect 21637 33915 21695 33921
rect 21637 33912 21649 33915
rect 21324 33884 21649 33912
rect 21324 33872 21330 33884
rect 21637 33881 21649 33884
rect 21683 33881 21695 33915
rect 21637 33875 21695 33881
rect 21749 33915 21807 33921
rect 21749 33881 21761 33915
rect 21795 33912 21807 33915
rect 21795 33884 21864 33912
rect 21795 33881 21807 33884
rect 21749 33875 21807 33881
rect 1762 33844 1768 33856
rect 1723 33816 1768 33844
rect 1762 33804 1768 33816
rect 1820 33804 1826 33856
rect 17126 33804 17132 33856
rect 17184 33844 17190 33856
rect 21836 33844 21864 33884
rect 17184 33816 21864 33844
rect 22005 33847 22063 33853
rect 17184 33804 17190 33816
rect 22005 33813 22017 33847
rect 22051 33844 22063 33847
rect 22572 33844 22600 33943
rect 23014 33940 23020 33952
rect 23072 33940 23078 33992
rect 24486 33940 24492 33992
rect 24544 33980 24550 33992
rect 24581 33983 24639 33989
rect 24581 33980 24593 33983
rect 24544 33952 24593 33980
rect 24544 33940 24550 33952
rect 24581 33949 24593 33952
rect 24627 33949 24639 33983
rect 24581 33943 24639 33949
rect 24729 33983 24787 33989
rect 24729 33949 24741 33983
rect 24775 33980 24787 33983
rect 24964 33980 24992 34020
rect 24775 33952 24992 33980
rect 25087 33983 25145 33989
rect 24775 33949 24787 33952
rect 24729 33943 24787 33949
rect 25087 33949 25099 33983
rect 25133 33980 25145 33983
rect 25314 33980 25320 33992
rect 25133 33952 25320 33980
rect 25133 33949 25145 33952
rect 25087 33943 25145 33949
rect 25314 33940 25320 33952
rect 25372 33940 25378 33992
rect 23293 33915 23351 33921
rect 23293 33881 23305 33915
rect 23339 33912 23351 33915
rect 24026 33912 24032 33924
rect 23339 33884 24032 33912
rect 23339 33881 23351 33884
rect 23293 33875 23351 33881
rect 24026 33872 24032 33884
rect 24084 33872 24090 33924
rect 24854 33912 24860 33924
rect 24815 33884 24860 33912
rect 24854 33872 24860 33884
rect 24912 33872 24918 33924
rect 24949 33915 25007 33921
rect 24949 33881 24961 33915
rect 24995 33881 25007 33915
rect 25516 33912 25544 34020
rect 46290 34008 46296 34020
rect 46348 34008 46354 34060
rect 26970 33912 26976 33924
rect 25516 33884 26976 33912
rect 24949 33875 25007 33881
rect 22051 33816 22600 33844
rect 22051 33813 22063 33816
rect 22005 33807 22063 33813
rect 22738 33804 22744 33856
rect 22796 33844 22802 33856
rect 24964 33844 24992 33875
rect 26970 33872 26976 33884
rect 27028 33872 27034 33924
rect 25222 33844 25228 33856
rect 22796 33816 24992 33844
rect 25183 33816 25228 33844
rect 22796 33804 22802 33816
rect 25222 33804 25228 33816
rect 25280 33804 25286 33856
rect 1104 33754 58880 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 58880 33754
rect 1104 33680 58880 33702
rect 1762 33600 1768 33652
rect 1820 33640 1826 33652
rect 17126 33640 17132 33652
rect 1820 33612 17132 33640
rect 1820 33600 1826 33612
rect 17126 33600 17132 33612
rect 17184 33600 17190 33652
rect 22278 33600 22284 33652
rect 22336 33640 22342 33652
rect 34146 33640 34152 33652
rect 22336 33612 34152 33640
rect 22336 33600 22342 33612
rect 34146 33600 34152 33612
rect 34204 33600 34210 33652
rect 40402 33640 40408 33652
rect 35912 33612 40408 33640
rect 1857 33575 1915 33581
rect 1857 33541 1869 33575
rect 1903 33572 1915 33575
rect 2314 33572 2320 33584
rect 1903 33544 2320 33572
rect 1903 33541 1915 33544
rect 1857 33535 1915 33541
rect 2314 33532 2320 33544
rect 2372 33532 2378 33584
rect 12158 33532 12164 33584
rect 12216 33572 12222 33584
rect 21177 33575 21235 33581
rect 21177 33572 21189 33575
rect 12216 33544 21189 33572
rect 12216 33532 12222 33544
rect 21177 33541 21189 33544
rect 21223 33541 21235 33575
rect 21450 33572 21456 33584
rect 21177 33535 21235 33541
rect 21284 33544 21456 33572
rect 1670 33504 1676 33516
rect 1631 33476 1676 33504
rect 1670 33464 1676 33476
rect 1728 33464 1734 33516
rect 20625 33507 20683 33513
rect 20625 33473 20637 33507
rect 20671 33504 20683 33507
rect 20901 33507 20959 33513
rect 20901 33504 20913 33507
rect 20671 33476 20913 33504
rect 20671 33473 20683 33476
rect 20625 33467 20683 33473
rect 20901 33473 20913 33476
rect 20947 33504 20959 33507
rect 20947 33476 21036 33504
rect 20947 33473 20959 33476
rect 20901 33467 20959 33473
rect 16942 33260 16948 33312
rect 17000 33300 17006 33312
rect 20898 33300 20904 33312
rect 17000 33272 20904 33300
rect 17000 33260 17006 33272
rect 20898 33260 20904 33272
rect 20956 33260 20962 33312
rect 21008 33300 21036 33476
rect 21082 33464 21088 33516
rect 21140 33504 21146 33516
rect 21284 33513 21312 33544
rect 21450 33532 21456 33544
rect 21508 33532 21514 33584
rect 22186 33513 22192 33516
rect 21269 33507 21327 33513
rect 21140 33476 21185 33504
rect 21140 33464 21146 33476
rect 21269 33473 21281 33507
rect 21315 33473 21327 33507
rect 22005 33507 22063 33513
rect 22005 33504 22017 33507
rect 21269 33467 21327 33473
rect 21468 33476 22017 33504
rect 21468 33377 21496 33476
rect 22005 33473 22017 33476
rect 22051 33473 22063 33507
rect 22005 33467 22063 33473
rect 22153 33507 22192 33513
rect 22153 33473 22165 33507
rect 22153 33467 22192 33473
rect 22186 33464 22192 33467
rect 22244 33464 22250 33516
rect 22296 33513 22324 33600
rect 35912 33572 35940 33612
rect 36078 33572 36084 33584
rect 26206 33544 35940 33572
rect 36039 33544 36084 33572
rect 22281 33507 22339 33513
rect 22281 33473 22293 33507
rect 22327 33473 22339 33507
rect 22281 33467 22339 33473
rect 22370 33464 22376 33516
rect 22428 33504 22434 33516
rect 22554 33513 22560 33516
rect 22511 33507 22560 33513
rect 22428 33476 22473 33504
rect 22428 33464 22434 33476
rect 22511 33473 22523 33507
rect 22557 33473 22560 33507
rect 22511 33467 22560 33473
rect 22554 33464 22560 33467
rect 22612 33464 22618 33516
rect 22830 33464 22836 33516
rect 22888 33504 22894 33516
rect 26206 33504 26234 33544
rect 36078 33532 36084 33544
rect 36136 33532 36142 33584
rect 22888 33476 26234 33504
rect 22888 33464 22894 33476
rect 32214 33464 32220 33516
rect 32272 33504 32278 33516
rect 35713 33507 35771 33513
rect 35713 33504 35725 33507
rect 32272 33476 35725 33504
rect 32272 33464 32278 33476
rect 35713 33473 35725 33476
rect 35759 33473 35771 33507
rect 35713 33467 35771 33473
rect 35802 33464 35808 33516
rect 35860 33504 35866 33516
rect 35860 33476 35905 33504
rect 35860 33464 35866 33476
rect 35986 33464 35992 33516
rect 36044 33504 36050 33516
rect 36188 33513 36216 33612
rect 40402 33600 40408 33612
rect 40460 33600 40466 33652
rect 36178 33507 36236 33513
rect 36044 33476 36089 33504
rect 36044 33464 36050 33476
rect 36178 33473 36190 33507
rect 36224 33473 36236 33507
rect 36178 33467 36236 33473
rect 40402 33436 40408 33448
rect 22480 33408 40408 33436
rect 21453 33371 21511 33377
rect 21453 33337 21465 33371
rect 21499 33337 21511 33371
rect 22480 33368 22508 33408
rect 40402 33396 40408 33408
rect 40460 33396 40466 33448
rect 21453 33331 21511 33337
rect 22066 33340 22508 33368
rect 22066 33300 22094 33340
rect 23290 33328 23296 33380
rect 23348 33368 23354 33380
rect 35986 33368 35992 33380
rect 23348 33340 35992 33368
rect 23348 33328 23354 33340
rect 35986 33328 35992 33340
rect 36044 33328 36050 33380
rect 22646 33300 22652 33312
rect 21008 33272 22094 33300
rect 22607 33272 22652 33300
rect 22646 33260 22652 33272
rect 22704 33260 22710 33312
rect 36357 33303 36415 33309
rect 36357 33269 36369 33303
rect 36403 33300 36415 33303
rect 37642 33300 37648 33312
rect 36403 33272 37648 33300
rect 36403 33269 36415 33272
rect 36357 33263 36415 33269
rect 37642 33260 37648 33272
rect 37700 33260 37706 33312
rect 1104 33210 58880 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 58880 33210
rect 1104 33136 58880 33158
rect 20898 33056 20904 33108
rect 20956 33096 20962 33108
rect 21726 33096 21732 33108
rect 20956 33068 21732 33096
rect 20956 33056 20962 33068
rect 21726 33056 21732 33068
rect 21784 33056 21790 33108
rect 21913 33031 21971 33037
rect 21913 32997 21925 33031
rect 21959 33028 21971 33031
rect 22646 33028 22652 33040
rect 21959 33000 22652 33028
rect 21959 32997 21971 33000
rect 21913 32991 21971 32997
rect 22646 32988 22652 33000
rect 22704 32988 22710 33040
rect 24857 33031 24915 33037
rect 24857 32997 24869 33031
rect 24903 33028 24915 33031
rect 25222 33028 25228 33040
rect 24903 33000 25228 33028
rect 24903 32997 24915 33000
rect 24857 32991 24915 32997
rect 25222 32988 25228 33000
rect 25280 32988 25286 33040
rect 58158 32960 58164 32972
rect 58119 32932 58164 32960
rect 58158 32920 58164 32932
rect 58216 32920 58222 32972
rect 21818 32892 21824 32904
rect 21779 32864 21824 32892
rect 21818 32852 21824 32864
rect 21876 32852 21882 32904
rect 22097 32895 22155 32901
rect 22097 32861 22109 32895
rect 22143 32892 22155 32895
rect 23198 32892 23204 32904
rect 22143 32864 23204 32892
rect 22143 32861 22155 32864
rect 22097 32855 22155 32861
rect 23198 32852 23204 32864
rect 23256 32852 23262 32904
rect 24762 32892 24768 32904
rect 24723 32864 24768 32892
rect 24762 32852 24768 32864
rect 24820 32852 24826 32904
rect 25041 32895 25099 32901
rect 25041 32861 25053 32895
rect 25087 32892 25099 32895
rect 37550 32892 37556 32904
rect 25087 32864 37556 32892
rect 25087 32861 25099 32864
rect 25041 32855 25099 32861
rect 37550 32852 37556 32864
rect 37608 32852 37614 32904
rect 56134 32852 56140 32904
rect 56192 32892 56198 32904
rect 57885 32895 57943 32901
rect 57885 32892 57897 32895
rect 56192 32864 57897 32892
rect 56192 32852 56198 32864
rect 57885 32861 57897 32864
rect 57931 32861 57943 32895
rect 57885 32855 57943 32861
rect 1670 32824 1676 32836
rect 1631 32796 1676 32824
rect 1670 32784 1676 32796
rect 1728 32784 1734 32836
rect 22186 32784 22192 32836
rect 22244 32824 22250 32836
rect 57054 32824 57060 32836
rect 22244 32796 25268 32824
rect 57015 32796 57060 32824
rect 22244 32784 22250 32796
rect 1765 32759 1823 32765
rect 1765 32725 1777 32759
rect 1811 32756 1823 32759
rect 16574 32756 16580 32768
rect 1811 32728 16580 32756
rect 1811 32725 1823 32728
rect 1765 32719 1823 32725
rect 16574 32716 16580 32728
rect 16632 32716 16638 32768
rect 22094 32716 22100 32768
rect 22152 32756 22158 32768
rect 25240 32765 25268 32796
rect 57054 32784 57060 32796
rect 57112 32784 57118 32836
rect 22281 32759 22339 32765
rect 22281 32756 22293 32759
rect 22152 32728 22293 32756
rect 22152 32716 22158 32728
rect 22281 32725 22293 32728
rect 22327 32725 22339 32759
rect 22281 32719 22339 32725
rect 25225 32759 25283 32765
rect 25225 32725 25237 32759
rect 25271 32725 25283 32759
rect 25225 32719 25283 32725
rect 55858 32716 55864 32768
rect 55916 32756 55922 32768
rect 57149 32759 57207 32765
rect 57149 32756 57161 32759
rect 55916 32728 57161 32756
rect 55916 32716 55922 32728
rect 57149 32725 57161 32728
rect 57195 32725 57207 32759
rect 57149 32719 57207 32725
rect 1104 32666 58880 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 58880 32666
rect 1104 32592 58880 32614
rect 16482 32444 16488 32496
rect 16540 32484 16546 32496
rect 22278 32484 22284 32496
rect 16540 32456 22284 32484
rect 16540 32444 16546 32456
rect 22278 32444 22284 32456
rect 22336 32444 22342 32496
rect 1670 32416 1676 32428
rect 1631 32388 1676 32416
rect 1670 32376 1676 32388
rect 1728 32376 1734 32428
rect 22002 32376 22008 32428
rect 22060 32416 22066 32428
rect 29178 32416 29184 32428
rect 22060 32388 29184 32416
rect 22060 32376 22066 32388
rect 29178 32376 29184 32388
rect 29236 32376 29242 32428
rect 1765 32215 1823 32221
rect 1765 32181 1777 32215
rect 1811 32212 1823 32215
rect 22738 32212 22744 32224
rect 1811 32184 22744 32212
rect 1811 32181 1823 32184
rect 1765 32175 1823 32181
rect 22738 32172 22744 32184
rect 22796 32172 22802 32224
rect 1104 32122 58880 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 58880 32122
rect 1104 32048 58880 32070
rect 20254 31900 20260 31952
rect 20312 31940 20318 31952
rect 22922 31940 22928 31952
rect 20312 31912 22928 31940
rect 20312 31900 20318 31912
rect 22922 31900 22928 31912
rect 22980 31940 22986 31952
rect 23290 31940 23296 31952
rect 22980 31912 23296 31940
rect 22980 31900 22986 31912
rect 22465 31875 22523 31881
rect 22465 31841 22477 31875
rect 22511 31872 22523 31875
rect 22511 31844 23060 31872
rect 22511 31841 22523 31844
rect 22465 31835 22523 31841
rect 22738 31804 22744 31816
rect 22699 31776 22744 31804
rect 22738 31764 22744 31776
rect 22796 31764 22802 31816
rect 23032 31813 23060 31844
rect 23124 31813 23152 31912
rect 23290 31900 23296 31912
rect 23348 31900 23354 31952
rect 58250 31940 58256 31952
rect 26206 31912 58256 31940
rect 26206 31872 26234 31912
rect 58250 31900 58256 31912
rect 58308 31900 58314 31952
rect 23216 31844 26234 31872
rect 23017 31807 23075 31813
rect 23017 31773 23029 31807
rect 23063 31773 23075 31807
rect 23017 31767 23075 31773
rect 23109 31807 23167 31813
rect 23109 31773 23121 31807
rect 23155 31773 23167 31807
rect 23109 31767 23167 31773
rect 21726 31696 21732 31748
rect 21784 31736 21790 31748
rect 22925 31739 22983 31745
rect 22925 31736 22937 31739
rect 21784 31708 22937 31736
rect 21784 31696 21790 31708
rect 22925 31705 22937 31708
rect 22971 31705 22983 31739
rect 23032 31736 23060 31767
rect 23216 31736 23244 31844
rect 49142 31764 49148 31816
rect 49200 31804 49206 31816
rect 57885 31807 57943 31813
rect 57885 31804 57897 31807
rect 49200 31776 57897 31804
rect 49200 31764 49206 31776
rect 57885 31773 57897 31776
rect 57931 31773 57943 31807
rect 58158 31804 58164 31816
rect 58119 31776 58164 31804
rect 57885 31767 57943 31773
rect 58158 31764 58164 31776
rect 58216 31764 58222 31816
rect 23032 31708 23244 31736
rect 22925 31699 22983 31705
rect 23290 31668 23296 31680
rect 23251 31640 23296 31668
rect 23290 31628 23296 31640
rect 23348 31628 23354 31680
rect 1104 31578 58880 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 58880 31578
rect 1104 31504 58880 31526
rect 19242 31424 19248 31476
rect 19300 31464 19306 31476
rect 24578 31464 24584 31476
rect 19300 31436 24584 31464
rect 19300 31424 19306 31436
rect 24578 31424 24584 31436
rect 24636 31424 24642 31476
rect 1670 31328 1676 31340
rect 1631 31300 1676 31328
rect 1670 31288 1676 31300
rect 1728 31288 1734 31340
rect 24118 31328 24124 31340
rect 24079 31300 24124 31328
rect 24118 31288 24124 31300
rect 24176 31288 24182 31340
rect 24210 31288 24216 31340
rect 24268 31328 24274 31340
rect 24397 31331 24455 31337
rect 24268 31300 24313 31328
rect 24268 31288 24274 31300
rect 24397 31297 24409 31331
rect 24443 31297 24455 31331
rect 24397 31291 24455 31297
rect 24489 31331 24547 31337
rect 24489 31297 24501 31331
rect 24535 31297 24547 31331
rect 24489 31291 24547 31297
rect 21266 31220 21272 31272
rect 21324 31260 21330 31272
rect 22738 31260 22744 31272
rect 21324 31232 22744 31260
rect 21324 31220 21330 31232
rect 22738 31220 22744 31232
rect 22796 31260 22802 31272
rect 24412 31260 24440 31291
rect 22796 31232 24440 31260
rect 22796 31220 22802 31232
rect 10318 31152 10324 31204
rect 10376 31192 10382 31204
rect 21818 31192 21824 31204
rect 10376 31164 21824 31192
rect 10376 31152 10382 31164
rect 21818 31152 21824 31164
rect 21876 31152 21882 31204
rect 1765 31127 1823 31133
rect 1765 31093 1777 31127
rect 1811 31124 1823 31127
rect 24504 31124 24532 31291
rect 24578 31288 24584 31340
rect 24636 31337 24642 31340
rect 24636 31331 24663 31337
rect 24651 31297 24663 31331
rect 58066 31328 58072 31340
rect 58027 31300 58072 31328
rect 24636 31291 24663 31297
rect 24636 31288 24642 31291
rect 58066 31288 58072 31300
rect 58124 31288 58130 31340
rect 24762 31192 24768 31204
rect 24723 31164 24768 31192
rect 24762 31152 24768 31164
rect 24820 31152 24826 31204
rect 1811 31096 24532 31124
rect 1811 31093 1823 31096
rect 1765 31087 1823 31093
rect 44174 31084 44180 31136
rect 44232 31124 44238 31136
rect 49786 31124 49792 31136
rect 44232 31096 49792 31124
rect 44232 31084 44238 31096
rect 49786 31084 49792 31096
rect 49844 31084 49850 31136
rect 58253 31127 58311 31133
rect 58253 31093 58265 31127
rect 58299 31124 58311 31127
rect 59170 31124 59176 31136
rect 58299 31096 59176 31124
rect 58299 31093 58311 31096
rect 58253 31087 58311 31093
rect 59170 31084 59176 31096
rect 59228 31084 59234 31136
rect 1104 31034 58880 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 58880 31034
rect 1104 30960 58880 30982
rect 23201 30923 23259 30929
rect 23201 30889 23213 30923
rect 23247 30920 23259 30923
rect 23290 30920 23296 30932
rect 23247 30892 23296 30920
rect 23247 30889 23259 30892
rect 23201 30883 23259 30889
rect 23290 30880 23296 30892
rect 23348 30880 23354 30932
rect 24210 30880 24216 30932
rect 24268 30920 24274 30932
rect 29086 30920 29092 30932
rect 24268 30892 29092 30920
rect 24268 30880 24274 30892
rect 29086 30880 29092 30892
rect 29144 30880 29150 30932
rect 19334 30744 19340 30796
rect 19392 30784 19398 30796
rect 19521 30787 19579 30793
rect 19521 30784 19533 30787
rect 19392 30756 19533 30784
rect 19392 30744 19398 30756
rect 19521 30753 19533 30756
rect 19567 30753 19579 30787
rect 34698 30784 34704 30796
rect 19521 30747 19579 30753
rect 19628 30756 34704 30784
rect 19429 30719 19487 30725
rect 19429 30685 19441 30719
rect 19475 30716 19487 30719
rect 19628 30716 19656 30756
rect 34698 30744 34704 30756
rect 34756 30744 34762 30796
rect 19475 30688 19656 30716
rect 19705 30719 19763 30725
rect 19475 30685 19487 30688
rect 19429 30679 19487 30685
rect 19705 30685 19717 30719
rect 19751 30685 19763 30719
rect 23106 30716 23112 30728
rect 23067 30688 23112 30716
rect 19705 30679 19763 30685
rect 1670 30648 1676 30660
rect 1631 30620 1676 30648
rect 1670 30608 1676 30620
rect 1728 30608 1734 30660
rect 17678 30608 17684 30660
rect 17736 30648 17742 30660
rect 19720 30648 19748 30679
rect 23106 30676 23112 30688
rect 23164 30676 23170 30728
rect 23198 30676 23204 30728
rect 23256 30716 23262 30728
rect 23293 30719 23351 30725
rect 23293 30716 23305 30719
rect 23256 30688 23305 30716
rect 23256 30676 23262 30688
rect 23293 30685 23305 30688
rect 23339 30685 23351 30719
rect 23566 30716 23572 30728
rect 23527 30688 23572 30716
rect 23293 30679 23351 30685
rect 17736 30620 19748 30648
rect 20165 30651 20223 30657
rect 17736 30608 17742 30620
rect 20165 30617 20177 30651
rect 20211 30648 20223 30651
rect 20346 30648 20352 30660
rect 20211 30620 20352 30648
rect 20211 30617 20223 30620
rect 20165 30611 20223 30617
rect 20346 30608 20352 30620
rect 20404 30608 20410 30660
rect 22278 30608 22284 30660
rect 22336 30648 22342 30660
rect 22833 30651 22891 30657
rect 22833 30648 22845 30651
rect 22336 30620 22845 30648
rect 22336 30608 22342 30620
rect 22833 30617 22845 30620
rect 22879 30617 22891 30651
rect 23308 30648 23336 30679
rect 23566 30676 23572 30688
rect 23624 30676 23630 30728
rect 32214 30648 32220 30660
rect 23308 30620 32220 30648
rect 22833 30611 22891 30617
rect 32214 30608 32220 30620
rect 32272 30608 32278 30660
rect 1765 30583 1823 30589
rect 1765 30549 1777 30583
rect 1811 30580 1823 30583
rect 17954 30580 17960 30592
rect 1811 30552 17960 30580
rect 1811 30549 1823 30552
rect 1765 30543 1823 30549
rect 17954 30540 17960 30552
rect 18012 30540 18018 30592
rect 22557 30583 22615 30589
rect 22557 30549 22569 30583
rect 22603 30580 22615 30583
rect 23477 30583 23535 30589
rect 23477 30580 23489 30583
rect 22603 30552 23489 30580
rect 22603 30549 22615 30552
rect 22557 30543 22615 30549
rect 23477 30549 23489 30552
rect 23523 30580 23535 30583
rect 24854 30580 24860 30592
rect 23523 30552 24860 30580
rect 23523 30549 23535 30552
rect 23477 30543 23535 30549
rect 24854 30540 24860 30552
rect 24912 30540 24918 30592
rect 1104 30490 58880 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 58880 30490
rect 1104 30416 58880 30438
rect 17954 30336 17960 30388
rect 18012 30376 18018 30388
rect 19334 30376 19340 30388
rect 18012 30348 19104 30376
rect 19295 30348 19340 30376
rect 18012 30336 18018 30348
rect 15102 30268 15108 30320
rect 15160 30308 15166 30320
rect 19076 30317 19104 30348
rect 19334 30336 19340 30348
rect 19392 30336 19398 30388
rect 19061 30311 19119 30317
rect 15160 30280 19012 30308
rect 15160 30268 15166 30280
rect 18984 30252 19012 30280
rect 19061 30277 19073 30311
rect 19107 30277 19119 30311
rect 19061 30271 19119 30277
rect 1578 30240 1584 30252
rect 1539 30212 1584 30240
rect 1578 30200 1584 30212
rect 1636 30200 1642 30252
rect 18874 30249 18880 30252
rect 18693 30243 18751 30249
rect 18693 30209 18705 30243
rect 18739 30209 18751 30243
rect 18693 30203 18751 30209
rect 18841 30243 18880 30249
rect 18841 30209 18853 30243
rect 18841 30203 18880 30209
rect 1762 30172 1768 30184
rect 1723 30144 1768 30172
rect 1762 30132 1768 30144
rect 1820 30132 1826 30184
rect 18708 30104 18736 30203
rect 18874 30200 18880 30203
rect 18932 30200 18938 30252
rect 18966 30200 18972 30252
rect 19024 30240 19030 30252
rect 19242 30249 19248 30252
rect 19199 30243 19248 30249
rect 19024 30212 19117 30240
rect 19024 30200 19030 30212
rect 19199 30209 19211 30243
rect 19245 30209 19248 30243
rect 19199 30203 19248 30209
rect 19242 30200 19248 30203
rect 19300 30200 19306 30252
rect 22278 30240 22284 30252
rect 22239 30212 22284 30240
rect 22278 30200 22284 30212
rect 22336 30200 22342 30252
rect 22554 30240 22560 30252
rect 22515 30212 22560 30240
rect 22554 30200 22560 30212
rect 22612 30200 22618 30252
rect 21634 30132 21640 30184
rect 21692 30172 21698 30184
rect 22373 30175 22431 30181
rect 22373 30172 22385 30175
rect 21692 30144 22385 30172
rect 21692 30132 21698 30144
rect 22373 30141 22385 30144
rect 22419 30141 22431 30175
rect 22373 30135 22431 30141
rect 22462 30132 22468 30184
rect 22520 30172 22526 30184
rect 22741 30175 22799 30181
rect 22741 30172 22753 30175
rect 22520 30144 22753 30172
rect 22520 30132 22526 30144
rect 22741 30141 22753 30144
rect 22787 30141 22799 30175
rect 22741 30135 22799 30141
rect 24118 30104 24124 30116
rect 18708 30076 24124 30104
rect 24118 30064 24124 30076
rect 24176 30064 24182 30116
rect 1104 29946 58880 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 58880 29946
rect 1104 29872 58880 29894
rect 22097 29835 22155 29841
rect 22097 29801 22109 29835
rect 22143 29832 22155 29835
rect 22554 29832 22560 29844
rect 22143 29804 22560 29832
rect 22143 29801 22155 29804
rect 22097 29795 22155 29801
rect 22554 29792 22560 29804
rect 22612 29792 22618 29844
rect 23106 29832 23112 29844
rect 23067 29804 23112 29832
rect 23106 29792 23112 29804
rect 23164 29792 23170 29844
rect 13814 29656 13820 29708
rect 13872 29696 13878 29708
rect 33134 29696 33140 29708
rect 13872 29668 22094 29696
rect 13872 29656 13878 29668
rect 1581 29631 1639 29637
rect 1581 29597 1593 29631
rect 1627 29628 1639 29631
rect 1946 29628 1952 29640
rect 1627 29600 1952 29628
rect 1627 29597 1639 29600
rect 1581 29591 1639 29597
rect 1946 29588 1952 29600
rect 2004 29588 2010 29640
rect 2590 29588 2596 29640
rect 2648 29628 2654 29640
rect 9950 29628 9956 29640
rect 2648 29600 9956 29628
rect 2648 29588 2654 29600
rect 9950 29588 9956 29600
rect 10008 29588 10014 29640
rect 21542 29628 21548 29640
rect 21503 29600 21548 29628
rect 21542 29588 21548 29600
rect 21600 29588 21606 29640
rect 21910 29628 21916 29640
rect 21871 29600 21916 29628
rect 21910 29588 21916 29600
rect 21968 29588 21974 29640
rect 1854 29560 1860 29572
rect 1815 29532 1860 29560
rect 1854 29520 1860 29532
rect 1912 29520 1918 29572
rect 18966 29520 18972 29572
rect 19024 29560 19030 29572
rect 21729 29563 21787 29569
rect 21729 29560 21741 29563
rect 19024 29532 21741 29560
rect 19024 29520 19030 29532
rect 21729 29529 21741 29532
rect 21775 29529 21787 29563
rect 21729 29523 21787 29529
rect 21744 29492 21772 29523
rect 21818 29520 21824 29572
rect 21876 29560 21882 29572
rect 22066 29560 22094 29668
rect 22572 29668 33140 29696
rect 22572 29637 22600 29668
rect 33134 29656 33140 29668
rect 33192 29656 33198 29708
rect 35526 29656 35532 29708
rect 35584 29696 35590 29708
rect 51718 29696 51724 29708
rect 35584 29668 51724 29696
rect 35584 29656 35590 29668
rect 51718 29656 51724 29668
rect 51776 29656 51782 29708
rect 58158 29696 58164 29708
rect 58119 29668 58164 29696
rect 58158 29656 58164 29668
rect 58216 29656 58222 29708
rect 22557 29631 22615 29637
rect 22557 29597 22569 29631
rect 22603 29597 22615 29631
rect 22833 29631 22891 29637
rect 22833 29628 22845 29631
rect 22557 29591 22615 29597
rect 22664 29600 22845 29628
rect 22664 29560 22692 29600
rect 22833 29597 22845 29600
rect 22879 29597 22891 29631
rect 22833 29591 22891 29597
rect 22925 29631 22983 29637
rect 22925 29597 22937 29631
rect 22971 29628 22983 29631
rect 23014 29628 23020 29640
rect 22971 29600 23020 29628
rect 22971 29597 22983 29600
rect 22925 29591 22983 29597
rect 23014 29588 23020 29600
rect 23072 29588 23078 29640
rect 57146 29588 57152 29640
rect 57204 29628 57210 29640
rect 57885 29631 57943 29637
rect 57885 29628 57897 29631
rect 57204 29600 57897 29628
rect 57204 29588 57210 29600
rect 57885 29597 57897 29600
rect 57931 29597 57943 29631
rect 57885 29591 57943 29597
rect 21876 29532 21921 29560
rect 22066 29532 22692 29560
rect 21876 29520 21882 29532
rect 22738 29520 22744 29572
rect 22796 29560 22802 29572
rect 23382 29560 23388 29572
rect 22796 29532 23388 29560
rect 22796 29520 22802 29532
rect 23382 29520 23388 29532
rect 23440 29520 23446 29572
rect 57054 29560 57060 29572
rect 57015 29532 57060 29560
rect 57054 29520 57060 29532
rect 57112 29520 57118 29572
rect 24946 29492 24952 29504
rect 21744 29464 24952 29492
rect 24946 29452 24952 29464
rect 25004 29452 25010 29504
rect 44818 29452 44824 29504
rect 44876 29492 44882 29504
rect 57149 29495 57207 29501
rect 57149 29492 57161 29495
rect 44876 29464 57161 29492
rect 44876 29452 44882 29464
rect 57149 29461 57161 29464
rect 57195 29461 57207 29495
rect 57149 29455 57207 29461
rect 1104 29402 58880 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 58880 29402
rect 1104 29328 58880 29350
rect 1578 29248 1584 29300
rect 1636 29288 1642 29300
rect 9677 29291 9735 29297
rect 9677 29288 9689 29291
rect 1636 29260 9689 29288
rect 1636 29248 1642 29260
rect 9677 29257 9689 29260
rect 9723 29257 9735 29291
rect 9677 29251 9735 29257
rect 21542 29248 21548 29300
rect 21600 29288 21606 29300
rect 49050 29288 49056 29300
rect 21600 29260 49056 29288
rect 21600 29248 21606 29260
rect 49050 29248 49056 29260
rect 49108 29248 49114 29300
rect 9309 29155 9367 29161
rect 9309 29121 9321 29155
rect 9355 29121 9367 29155
rect 9309 29115 9367 29121
rect 9463 29155 9521 29161
rect 9463 29121 9475 29155
rect 9509 29152 9521 29155
rect 15102 29152 15108 29164
rect 9509 29124 15108 29152
rect 9509 29121 9521 29124
rect 9463 29115 9521 29121
rect 9324 29084 9352 29115
rect 15102 29112 15108 29124
rect 15160 29112 15166 29164
rect 21726 29112 21732 29164
rect 21784 29152 21790 29164
rect 23014 29152 23020 29164
rect 21784 29124 23020 29152
rect 21784 29112 21790 29124
rect 23014 29112 23020 29124
rect 23072 29112 23078 29164
rect 9674 29084 9680 29096
rect 9324 29056 9680 29084
rect 9674 29044 9680 29056
rect 9732 29044 9738 29096
rect 1104 28858 58880 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 58880 28858
rect 1104 28784 58880 28806
rect 2869 28611 2927 28617
rect 2869 28608 2881 28611
rect 1596 28580 2881 28608
rect 1596 28549 1624 28580
rect 2869 28577 2881 28580
rect 2915 28577 2927 28611
rect 2869 28571 2927 28577
rect 5534 28568 5540 28620
rect 5592 28608 5598 28620
rect 29270 28608 29276 28620
rect 5592 28580 29276 28608
rect 5592 28568 5598 28580
rect 29270 28568 29276 28580
rect 29328 28568 29334 28620
rect 1581 28543 1639 28549
rect 1581 28509 1593 28543
rect 1627 28509 1639 28543
rect 1581 28503 1639 28509
rect 2501 28543 2559 28549
rect 2501 28509 2513 28543
rect 2547 28509 2559 28543
rect 2501 28503 2559 28509
rect 2655 28543 2713 28549
rect 2655 28509 2667 28543
rect 2701 28540 2713 28543
rect 2958 28540 2964 28552
rect 2701 28512 2964 28540
rect 2701 28509 2713 28512
rect 2655 28503 2713 28509
rect 1854 28472 1860 28484
rect 1815 28444 1860 28472
rect 1854 28432 1860 28444
rect 1912 28432 1918 28484
rect 2516 28472 2544 28503
rect 2958 28500 2964 28512
rect 3016 28500 3022 28552
rect 8938 28500 8944 28552
rect 8996 28540 9002 28552
rect 8996 28512 9812 28540
rect 8996 28500 9002 28512
rect 9674 28472 9680 28484
rect 2516 28444 9680 28472
rect 9674 28432 9680 28444
rect 9732 28432 9738 28484
rect 9784 28472 9812 28512
rect 12802 28500 12808 28552
rect 12860 28540 12866 28552
rect 22646 28540 22652 28552
rect 12860 28512 22652 28540
rect 12860 28500 12866 28512
rect 22646 28500 22652 28512
rect 22704 28540 22710 28552
rect 23290 28540 23296 28552
rect 22704 28512 23296 28540
rect 22704 28500 22710 28512
rect 23290 28500 23296 28512
rect 23348 28500 23354 28552
rect 29086 28500 29092 28552
rect 29144 28540 29150 28552
rect 46474 28540 46480 28552
rect 29144 28512 46480 28540
rect 29144 28500 29150 28512
rect 46474 28500 46480 28512
rect 46532 28500 46538 28552
rect 55582 28500 55588 28552
rect 55640 28540 55646 28552
rect 57885 28543 57943 28549
rect 57885 28540 57897 28543
rect 55640 28512 57897 28540
rect 55640 28500 55646 28512
rect 57885 28509 57897 28512
rect 57931 28509 57943 28543
rect 57885 28503 57943 28509
rect 34054 28472 34060 28484
rect 9784 28444 34060 28472
rect 34054 28432 34060 28444
rect 34112 28432 34118 28484
rect 58158 28472 58164 28484
rect 58119 28444 58164 28472
rect 58158 28432 58164 28444
rect 58216 28432 58222 28484
rect 20438 28364 20444 28416
rect 20496 28404 20502 28416
rect 47302 28404 47308 28416
rect 20496 28376 47308 28404
rect 20496 28364 20502 28376
rect 47302 28364 47308 28376
rect 47360 28364 47366 28416
rect 1104 28314 58880 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 58880 28314
rect 1104 28240 58880 28262
rect 22830 28092 22836 28144
rect 22888 28132 22894 28144
rect 23293 28135 23351 28141
rect 22888 28104 23244 28132
rect 22888 28092 22894 28104
rect 1581 28067 1639 28073
rect 1581 28033 1593 28067
rect 1627 28064 1639 28067
rect 2222 28064 2228 28076
rect 1627 28036 2228 28064
rect 1627 28033 1639 28036
rect 1581 28027 1639 28033
rect 2222 28024 2228 28036
rect 2280 28024 2286 28076
rect 23106 28064 23112 28076
rect 23067 28036 23112 28064
rect 23106 28024 23112 28036
rect 23164 28024 23170 28076
rect 23216 28064 23244 28104
rect 23293 28101 23305 28135
rect 23339 28132 23351 28135
rect 23566 28132 23572 28144
rect 23339 28104 23572 28132
rect 23339 28101 23351 28104
rect 23293 28095 23351 28101
rect 23566 28092 23572 28104
rect 23624 28092 23630 28144
rect 23385 28067 23443 28073
rect 23385 28064 23397 28067
rect 23216 28036 23397 28064
rect 23385 28033 23397 28036
rect 23431 28033 23443 28067
rect 23385 28027 23443 28033
rect 23477 28067 23535 28073
rect 23477 28033 23489 28067
rect 23523 28064 23535 28067
rect 37274 28064 37280 28076
rect 23523 28036 37280 28064
rect 23523 28033 23535 28036
rect 23477 28027 23535 28033
rect 1762 27996 1768 28008
rect 1723 27968 1768 27996
rect 1762 27956 1768 27968
rect 1820 27956 1826 28008
rect 23290 27956 23296 28008
rect 23348 27996 23354 28008
rect 23492 27996 23520 28027
rect 37274 28024 37280 28036
rect 37332 28024 37338 28076
rect 23348 27968 23520 27996
rect 23348 27956 23354 27968
rect 23014 27820 23020 27872
rect 23072 27860 23078 27872
rect 23661 27863 23719 27869
rect 23661 27860 23673 27863
rect 23072 27832 23673 27860
rect 23072 27820 23078 27832
rect 23661 27829 23673 27832
rect 23707 27829 23719 27863
rect 23661 27823 23719 27829
rect 1104 27770 58880 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 58880 27770
rect 1104 27696 58880 27718
rect 23658 27616 23664 27668
rect 23716 27616 23722 27668
rect 6886 27560 23520 27588
rect 2130 27480 2136 27532
rect 2188 27520 2194 27532
rect 6886 27520 6914 27560
rect 2188 27492 6914 27520
rect 2188 27480 2194 27492
rect 1578 27452 1584 27464
rect 1539 27424 1584 27452
rect 1578 27412 1584 27424
rect 1636 27412 1642 27464
rect 23014 27412 23020 27464
rect 23072 27452 23078 27464
rect 23290 27461 23296 27464
rect 23109 27455 23167 27461
rect 23109 27452 23121 27455
rect 23072 27424 23121 27452
rect 23072 27412 23078 27424
rect 23109 27421 23121 27424
rect 23155 27421 23167 27455
rect 23109 27415 23167 27421
rect 23257 27455 23296 27461
rect 23257 27421 23269 27455
rect 23257 27415 23296 27421
rect 23290 27412 23296 27415
rect 23348 27412 23354 27464
rect 1854 27384 1860 27396
rect 1815 27356 1860 27384
rect 1854 27344 1860 27356
rect 1912 27344 1918 27396
rect 23382 27384 23388 27396
rect 23343 27356 23388 27384
rect 23382 27344 23388 27356
rect 23440 27344 23446 27396
rect 23492 27393 23520 27560
rect 23676 27520 23704 27616
rect 31110 27548 31116 27600
rect 31168 27588 31174 27600
rect 33778 27588 33784 27600
rect 31168 27560 33784 27588
rect 31168 27548 31174 27560
rect 33778 27548 33784 27560
rect 33836 27548 33842 27600
rect 23589 27492 23704 27520
rect 23589 27461 23617 27492
rect 23574 27455 23632 27461
rect 23574 27421 23586 27455
rect 23620 27421 23632 27455
rect 57974 27452 57980 27464
rect 57935 27424 57980 27452
rect 23574 27415 23632 27421
rect 57974 27412 57980 27424
rect 58032 27412 58038 27464
rect 23477 27387 23535 27393
rect 23477 27353 23489 27387
rect 23523 27353 23535 27387
rect 23477 27347 23535 27353
rect 22830 27276 22836 27328
rect 22888 27316 22894 27328
rect 23753 27319 23811 27325
rect 23753 27316 23765 27319
rect 22888 27288 23765 27316
rect 22888 27276 22894 27288
rect 23753 27285 23765 27288
rect 23799 27285 23811 27319
rect 58066 27316 58072 27328
rect 58027 27288 58072 27316
rect 23753 27279 23811 27285
rect 58066 27276 58072 27288
rect 58124 27276 58130 27328
rect 1104 27226 58880 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 58880 27226
rect 1104 27152 58880 27174
rect 1578 27072 1584 27124
rect 1636 27112 1642 27124
rect 2869 27115 2927 27121
rect 2869 27112 2881 27115
rect 1636 27084 2881 27112
rect 1636 27072 1642 27084
rect 2869 27081 2881 27084
rect 2915 27081 2927 27115
rect 2869 27075 2927 27081
rect 28350 27072 28356 27124
rect 28408 27112 28414 27124
rect 41690 27112 41696 27124
rect 28408 27084 41696 27112
rect 28408 27072 28414 27084
rect 41690 27072 41696 27084
rect 41748 27072 41754 27124
rect 18874 27004 18880 27056
rect 18932 27044 18938 27056
rect 50982 27044 50988 27056
rect 18932 27016 50988 27044
rect 18932 27004 18938 27016
rect 50982 27004 50988 27016
rect 51040 27004 51046 27056
rect 1578 26976 1584 26988
rect 1539 26948 1584 26976
rect 1578 26936 1584 26948
rect 1636 26936 1642 26988
rect 2498 26976 2504 26988
rect 2459 26948 2504 26976
rect 2498 26936 2504 26948
rect 2556 26936 2562 26988
rect 2590 26936 2596 26988
rect 2648 26976 2654 26988
rect 2648 26948 2693 26976
rect 2648 26936 2654 26948
rect 7834 26936 7840 26988
rect 7892 26976 7898 26988
rect 22741 26979 22799 26985
rect 22741 26976 22753 26979
rect 7892 26948 22753 26976
rect 7892 26936 7898 26948
rect 22741 26945 22753 26948
rect 22787 26945 22799 26979
rect 22741 26939 22799 26945
rect 22830 26936 22836 26988
rect 22888 26976 22894 26988
rect 23017 26979 23075 26985
rect 22888 26948 22933 26976
rect 22888 26936 22894 26948
rect 23017 26945 23029 26979
rect 23063 26976 23075 26979
rect 23198 26976 23204 26988
rect 23063 26948 23204 26976
rect 23063 26945 23075 26948
rect 23017 26939 23075 26945
rect 23198 26936 23204 26948
rect 23256 26936 23262 26988
rect 33134 26936 33140 26988
rect 33192 26976 33198 26988
rect 47486 26976 47492 26988
rect 33192 26948 47492 26976
rect 33192 26936 33198 26948
rect 47486 26936 47492 26948
rect 47544 26936 47550 26988
rect 1762 26908 1768 26920
rect 1723 26880 1768 26908
rect 1762 26868 1768 26880
rect 1820 26868 1826 26920
rect 20714 26868 20720 26920
rect 20772 26908 20778 26920
rect 23385 26911 23443 26917
rect 23385 26908 23397 26911
rect 20772 26880 23397 26908
rect 20772 26868 20778 26880
rect 23385 26877 23397 26880
rect 23431 26877 23443 26911
rect 23385 26871 23443 26877
rect 23400 26840 23428 26871
rect 26878 26868 26884 26920
rect 26936 26908 26942 26920
rect 27798 26908 27804 26920
rect 26936 26880 27804 26908
rect 26936 26868 26942 26880
rect 27798 26868 27804 26880
rect 27856 26868 27862 26920
rect 36630 26868 36636 26920
rect 36688 26908 36694 26920
rect 55858 26908 55864 26920
rect 36688 26880 55864 26908
rect 36688 26868 36694 26880
rect 55858 26868 55864 26880
rect 55916 26868 55922 26920
rect 27246 26840 27252 26852
rect 23400 26812 27252 26840
rect 27246 26800 27252 26812
rect 27304 26800 27310 26852
rect 1104 26682 58880 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 58880 26682
rect 1104 26608 58880 26630
rect 58158 26432 58164 26444
rect 58119 26404 58164 26432
rect 58158 26392 58164 26404
rect 58216 26392 58222 26444
rect 57882 26364 57888 26376
rect 57843 26336 57888 26364
rect 57882 26324 57888 26336
rect 57940 26324 57946 26376
rect 28442 26256 28448 26308
rect 28500 26296 28506 26308
rect 29638 26296 29644 26308
rect 28500 26268 29644 26296
rect 28500 26256 28506 26268
rect 29638 26256 29644 26268
rect 29696 26256 29702 26308
rect 1104 26138 58880 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 58880 26138
rect 1104 26064 58880 26086
rect 1581 25891 1639 25897
rect 1581 25857 1593 25891
rect 1627 25888 1639 25891
rect 1627 25860 6914 25888
rect 1627 25857 1639 25860
rect 1581 25851 1639 25857
rect 1762 25820 1768 25832
rect 1723 25792 1768 25820
rect 1762 25780 1768 25792
rect 1820 25780 1826 25832
rect 6886 25684 6914 25860
rect 9674 25848 9680 25900
rect 9732 25888 9738 25900
rect 10686 25888 10692 25900
rect 9732 25860 10692 25888
rect 9732 25848 9738 25860
rect 10686 25848 10692 25860
rect 10744 25848 10750 25900
rect 10843 25891 10901 25897
rect 10843 25857 10855 25891
rect 10889 25888 10901 25891
rect 17218 25888 17224 25900
rect 10889 25860 17224 25888
rect 10889 25857 10901 25860
rect 10843 25851 10901 25857
rect 17218 25848 17224 25860
rect 17276 25848 17282 25900
rect 58066 25888 58072 25900
rect 58027 25860 58072 25888
rect 58066 25848 58072 25860
rect 58124 25848 58130 25900
rect 18414 25780 18420 25832
rect 18472 25820 18478 25832
rect 34514 25820 34520 25832
rect 18472 25792 34520 25820
rect 18472 25780 18478 25792
rect 34514 25780 34520 25792
rect 34572 25780 34578 25832
rect 23106 25712 23112 25764
rect 23164 25752 23170 25764
rect 40310 25752 40316 25764
rect 23164 25724 40316 25752
rect 23164 25712 23170 25724
rect 40310 25712 40316 25724
rect 40368 25712 40374 25764
rect 10873 25687 10931 25693
rect 10873 25684 10885 25687
rect 6886 25656 10885 25684
rect 10873 25653 10885 25656
rect 10919 25653 10931 25687
rect 10873 25647 10931 25653
rect 23290 25644 23296 25696
rect 23348 25684 23354 25696
rect 48866 25684 48872 25696
rect 23348 25656 48872 25684
rect 23348 25644 23354 25656
rect 48866 25644 48872 25656
rect 48924 25644 48930 25696
rect 57974 25644 57980 25696
rect 58032 25684 58038 25696
rect 58253 25687 58311 25693
rect 58253 25684 58265 25687
rect 58032 25656 58265 25684
rect 58032 25644 58038 25656
rect 58253 25653 58265 25656
rect 58299 25653 58311 25687
rect 58253 25647 58311 25653
rect 1104 25594 58880 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 58880 25594
rect 1104 25520 58880 25542
rect 17218 25440 17224 25492
rect 17276 25480 17282 25492
rect 22554 25480 22560 25492
rect 17276 25452 22560 25480
rect 17276 25440 17282 25452
rect 22554 25440 22560 25452
rect 22612 25480 22618 25492
rect 27430 25480 27436 25492
rect 22612 25452 27436 25480
rect 22612 25440 22618 25452
rect 27430 25440 27436 25452
rect 27488 25440 27494 25492
rect 2869 25347 2927 25353
rect 2869 25344 2881 25347
rect 1596 25316 2881 25344
rect 1596 25285 1624 25316
rect 2869 25313 2881 25316
rect 2915 25313 2927 25347
rect 2869 25307 2927 25313
rect 1581 25279 1639 25285
rect 1581 25245 1593 25279
rect 1627 25245 1639 25279
rect 2498 25276 2504 25288
rect 2411 25248 2504 25276
rect 1581 25239 1639 25245
rect 2498 25236 2504 25248
rect 2556 25236 2562 25288
rect 2590 25236 2596 25288
rect 2648 25276 2654 25288
rect 2648 25248 2693 25276
rect 2648 25236 2654 25248
rect 44450 25236 44456 25288
rect 44508 25276 44514 25288
rect 57885 25279 57943 25285
rect 57885 25276 57897 25279
rect 44508 25248 57897 25276
rect 44508 25236 44514 25248
rect 57885 25245 57897 25248
rect 57931 25245 57943 25279
rect 57885 25239 57943 25245
rect 1854 25208 1860 25220
rect 1815 25180 1860 25208
rect 1854 25168 1860 25180
rect 1912 25168 1918 25220
rect 2516 25208 2544 25236
rect 2866 25208 2872 25220
rect 2516 25180 2872 25208
rect 2866 25168 2872 25180
rect 2924 25168 2930 25220
rect 58158 25208 58164 25220
rect 58119 25180 58164 25208
rect 58158 25168 58164 25180
rect 58216 25168 58222 25220
rect 1104 25050 58880 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 58880 25050
rect 1104 24976 58880 24998
rect 1581 24803 1639 24809
rect 1581 24769 1593 24803
rect 1627 24800 1639 24803
rect 3050 24800 3056 24812
rect 1627 24772 3056 24800
rect 1627 24769 1639 24772
rect 1581 24763 1639 24769
rect 3050 24760 3056 24772
rect 3108 24760 3114 24812
rect 58066 24800 58072 24812
rect 58027 24772 58072 24800
rect 58066 24760 58072 24772
rect 58124 24760 58130 24812
rect 1762 24732 1768 24744
rect 1723 24704 1768 24732
rect 1762 24692 1768 24704
rect 1820 24692 1826 24744
rect 58250 24596 58256 24608
rect 58211 24568 58256 24596
rect 58250 24556 58256 24568
rect 58308 24556 58314 24608
rect 1104 24506 58880 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 58880 24506
rect 1104 24432 58880 24454
rect 3050 24392 3056 24404
rect 3011 24364 3056 24392
rect 3050 24352 3056 24364
rect 3108 24352 3114 24404
rect 4798 24216 4804 24268
rect 4856 24256 4862 24268
rect 32398 24256 32404 24268
rect 4856 24228 32404 24256
rect 4856 24216 4862 24228
rect 32398 24216 32404 24228
rect 32456 24216 32462 24268
rect 1581 24191 1639 24197
rect 1581 24157 1593 24191
rect 1627 24188 1639 24191
rect 1627 24160 2820 24188
rect 1627 24157 1639 24160
rect 1581 24151 1639 24157
rect 1854 24120 1860 24132
rect 1815 24092 1860 24120
rect 1854 24080 1860 24092
rect 1912 24080 1918 24132
rect 2792 24120 2820 24160
rect 2866 24148 2872 24200
rect 2924 24188 2930 24200
rect 3023 24191 3081 24197
rect 2924 24160 2969 24188
rect 2924 24148 2930 24160
rect 3023 24157 3035 24191
rect 3069 24188 3081 24191
rect 30834 24188 30840 24200
rect 3069 24160 30840 24188
rect 3069 24157 3081 24160
rect 3023 24151 3081 24157
rect 30834 24148 30840 24160
rect 30892 24148 30898 24200
rect 12158 24120 12164 24132
rect 2792 24092 12164 24120
rect 12158 24080 12164 24092
rect 12216 24080 12222 24132
rect 13722 24080 13728 24132
rect 13780 24120 13786 24132
rect 26694 24120 26700 24132
rect 13780 24092 26700 24120
rect 13780 24080 13786 24092
rect 26694 24080 26700 24092
rect 26752 24080 26758 24132
rect 26970 24080 26976 24132
rect 27028 24120 27034 24132
rect 54938 24120 54944 24132
rect 27028 24092 54944 24120
rect 27028 24080 27034 24092
rect 54938 24080 54944 24092
rect 54996 24080 55002 24132
rect 1104 23962 58880 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 58880 23962
rect 1104 23888 58880 23910
rect 12802 23780 12808 23792
rect 12763 23752 12808 23780
rect 12802 23740 12808 23752
rect 12860 23740 12866 23792
rect 12253 23715 12311 23721
rect 12253 23681 12265 23715
rect 12299 23712 12311 23715
rect 13722 23712 13728 23724
rect 12299 23684 13728 23712
rect 12299 23681 12311 23684
rect 12253 23675 12311 23681
rect 13722 23672 13728 23684
rect 13780 23672 13786 23724
rect 46290 23536 46296 23588
rect 46348 23576 46354 23588
rect 47854 23576 47860 23588
rect 46348 23548 47860 23576
rect 46348 23536 46354 23548
rect 47854 23536 47860 23548
rect 47912 23536 47918 23588
rect 49510 23536 49516 23588
rect 49568 23576 49574 23588
rect 57514 23576 57520 23588
rect 49568 23548 57520 23576
rect 49568 23536 49574 23548
rect 57514 23536 57520 23548
rect 57572 23536 57578 23588
rect 32490 23468 32496 23520
rect 32548 23508 32554 23520
rect 33134 23508 33140 23520
rect 32548 23480 33140 23508
rect 32548 23468 32554 23480
rect 33134 23468 33140 23480
rect 33192 23468 33198 23520
rect 43622 23468 43628 23520
rect 43680 23508 43686 23520
rect 47578 23508 47584 23520
rect 43680 23480 47584 23508
rect 43680 23468 43686 23480
rect 47578 23468 47584 23480
rect 47636 23468 47642 23520
rect 47670 23468 47676 23520
rect 47728 23508 47734 23520
rect 48590 23508 48596 23520
rect 47728 23480 48596 23508
rect 47728 23468 47734 23480
rect 48590 23468 48596 23480
rect 48648 23468 48654 23520
rect 1104 23418 58880 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 58880 23418
rect 1104 23344 58880 23366
rect 12158 23304 12164 23316
rect 12119 23276 12164 23304
rect 12158 23264 12164 23276
rect 12216 23264 12222 23316
rect 26694 23264 26700 23316
rect 26752 23304 26758 23316
rect 29638 23304 29644 23316
rect 26752 23276 29644 23304
rect 26752 23264 26758 23276
rect 29638 23264 29644 23276
rect 29696 23264 29702 23316
rect 18233 23239 18291 23245
rect 18233 23205 18245 23239
rect 18279 23236 18291 23239
rect 18782 23236 18788 23248
rect 18279 23208 18788 23236
rect 18279 23205 18291 23208
rect 18233 23199 18291 23205
rect 18782 23196 18788 23208
rect 18840 23196 18846 23248
rect 23382 23168 23388 23180
rect 11900 23140 23388 23168
rect 1581 23103 1639 23109
rect 1581 23069 1593 23103
rect 1627 23100 1639 23103
rect 1627 23072 6914 23100
rect 1627 23069 1639 23072
rect 1581 23063 1639 23069
rect 1854 23032 1860 23044
rect 1815 23004 1860 23032
rect 1854 22992 1860 23004
rect 1912 22992 1918 23044
rect 6886 23032 6914 23072
rect 10134 23060 10140 23112
rect 10192 23100 10198 23112
rect 10686 23100 10692 23112
rect 10192 23072 10692 23100
rect 10192 23060 10198 23072
rect 10686 23060 10692 23072
rect 10744 23100 10750 23112
rect 10870 23100 10876 23112
rect 10744 23072 10876 23100
rect 10744 23060 10750 23072
rect 10870 23060 10876 23072
rect 10928 23060 10934 23112
rect 11027 23103 11085 23109
rect 11027 23069 11039 23103
rect 11073 23100 11085 23103
rect 11900 23100 11928 23140
rect 23382 23128 23388 23140
rect 23440 23168 23446 23180
rect 26602 23168 26608 23180
rect 23440 23140 26608 23168
rect 23440 23128 23446 23140
rect 26602 23128 26608 23140
rect 26660 23128 26666 23180
rect 58158 23168 58164 23180
rect 58119 23140 58164 23168
rect 58158 23128 58164 23140
rect 58216 23128 58222 23180
rect 11073 23072 11928 23100
rect 11977 23103 12035 23109
rect 11073 23069 11085 23072
rect 11027 23063 11085 23069
rect 11977 23069 11989 23103
rect 12023 23069 12035 23103
rect 11977 23063 12035 23069
rect 12131 23103 12189 23109
rect 12131 23069 12143 23103
rect 12177 23100 12189 23103
rect 12802 23100 12808 23112
rect 12177 23072 12808 23100
rect 12177 23069 12189 23072
rect 12131 23063 12189 23069
rect 11241 23035 11299 23041
rect 11241 23032 11253 23035
rect 6886 23004 11253 23032
rect 11241 23001 11253 23004
rect 11287 23001 11299 23035
rect 11241 22995 11299 23001
rect 10870 22924 10876 22976
rect 10928 22964 10934 22976
rect 11992 22964 12020 23063
rect 12802 23060 12808 23072
rect 12860 23060 12866 23112
rect 17862 23060 17868 23112
rect 17920 23100 17926 23112
rect 18509 23103 18567 23109
rect 18509 23100 18521 23103
rect 17920 23072 18521 23100
rect 17920 23060 17926 23072
rect 18509 23069 18521 23072
rect 18555 23069 18567 23103
rect 18509 23063 18567 23069
rect 44082 23060 44088 23112
rect 44140 23100 44146 23112
rect 57885 23103 57943 23109
rect 57885 23100 57897 23103
rect 44140 23072 57897 23100
rect 44140 23060 44146 23072
rect 57885 23069 57897 23072
rect 57931 23069 57943 23103
rect 57885 23063 57943 23069
rect 18230 23032 18236 23044
rect 18191 23004 18236 23032
rect 18230 22992 18236 23004
rect 18288 22992 18294 23044
rect 31294 22992 31300 23044
rect 31352 23032 31358 23044
rect 39666 23032 39672 23044
rect 31352 23004 39672 23032
rect 31352 22992 31358 23004
rect 39666 22992 39672 23004
rect 39724 22992 39730 23044
rect 10928 22936 12020 22964
rect 10928 22924 10934 22936
rect 17954 22924 17960 22976
rect 18012 22964 18018 22976
rect 18417 22967 18475 22973
rect 18417 22964 18429 22967
rect 18012 22936 18429 22964
rect 18012 22924 18018 22936
rect 18417 22933 18429 22936
rect 18463 22933 18475 22967
rect 18417 22927 18475 22933
rect 22554 22924 22560 22976
rect 22612 22964 22618 22976
rect 44818 22964 44824 22976
rect 22612 22936 44824 22964
rect 22612 22924 22618 22936
rect 44818 22924 44824 22936
rect 44876 22924 44882 22976
rect 1104 22874 58880 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 58880 22874
rect 1104 22800 58880 22822
rect 18230 22720 18236 22772
rect 18288 22760 18294 22772
rect 24946 22760 24952 22772
rect 18288 22732 24952 22760
rect 18288 22720 18294 22732
rect 17862 22692 17868 22704
rect 16960 22664 17868 22692
rect 1581 22627 1639 22633
rect 1581 22593 1593 22627
rect 1627 22624 1639 22627
rect 9674 22624 9680 22636
rect 1627 22596 9680 22624
rect 1627 22593 1639 22596
rect 1581 22587 1639 22593
rect 9674 22584 9680 22596
rect 9732 22584 9738 22636
rect 1762 22556 1768 22568
rect 1723 22528 1768 22556
rect 1762 22516 1768 22528
rect 1820 22516 1826 22568
rect 16666 22516 16672 22568
rect 16724 22556 16730 22568
rect 16960 22565 16988 22664
rect 17862 22652 17868 22664
rect 17920 22692 17926 22704
rect 19444 22701 19472 22732
rect 24946 22720 24952 22732
rect 25004 22720 25010 22772
rect 48682 22760 48688 22772
rect 31726 22732 48688 22760
rect 18417 22695 18475 22701
rect 18417 22692 18429 22695
rect 17920 22664 18429 22692
rect 17920 22652 17926 22664
rect 18417 22661 18429 22664
rect 18463 22661 18475 22695
rect 18417 22655 18475 22661
rect 19429 22695 19487 22701
rect 19429 22661 19441 22695
rect 19475 22661 19487 22695
rect 19629 22695 19687 22701
rect 19629 22692 19641 22695
rect 19429 22655 19487 22661
rect 19536 22664 19641 22692
rect 17037 22627 17095 22633
rect 17037 22593 17049 22627
rect 17083 22624 17095 22627
rect 17954 22624 17960 22636
rect 17083 22596 17960 22624
rect 17083 22593 17095 22596
rect 17037 22587 17095 22593
rect 17954 22584 17960 22596
rect 18012 22584 18018 22636
rect 18138 22624 18144 22636
rect 18099 22596 18144 22624
rect 18138 22584 18144 22596
rect 18196 22584 18202 22636
rect 18233 22627 18291 22633
rect 18233 22593 18245 22627
rect 18279 22624 18291 22627
rect 18322 22624 18328 22636
rect 18279 22596 18328 22624
rect 18279 22593 18291 22596
rect 18233 22587 18291 22593
rect 18322 22584 18328 22596
rect 18380 22584 18386 22636
rect 18432 22624 18460 22655
rect 19536 22624 19564 22664
rect 19629 22661 19641 22664
rect 19675 22661 19687 22695
rect 19629 22655 19687 22661
rect 21634 22652 21640 22704
rect 21692 22692 21698 22704
rect 31726 22692 31754 22732
rect 48682 22720 48688 22732
rect 48740 22720 48746 22772
rect 58158 22692 58164 22704
rect 21692 22664 31754 22692
rect 58119 22664 58164 22692
rect 21692 22652 21698 22664
rect 58158 22652 58164 22664
rect 58216 22652 58222 22704
rect 18432 22596 19564 22624
rect 24578 22584 24584 22636
rect 24636 22624 24642 22636
rect 25961 22627 26019 22633
rect 25961 22624 25973 22627
rect 24636 22596 25973 22624
rect 24636 22584 24642 22596
rect 25961 22593 25973 22596
rect 26007 22593 26019 22627
rect 25961 22587 26019 22593
rect 16945 22559 17003 22565
rect 16945 22556 16957 22559
rect 16724 22528 16957 22556
rect 16724 22516 16730 22528
rect 16945 22525 16957 22528
rect 16991 22525 17003 22559
rect 16945 22519 17003 22525
rect 16758 22380 16764 22432
rect 16816 22420 16822 22432
rect 17405 22423 17463 22429
rect 17405 22420 17417 22423
rect 16816 22392 17417 22420
rect 16816 22380 16822 22392
rect 17405 22389 17417 22392
rect 17451 22389 17463 22423
rect 17972 22420 18000 22584
rect 25590 22516 25596 22568
rect 25648 22556 25654 22568
rect 25777 22559 25835 22565
rect 25777 22556 25789 22559
rect 25648 22528 25789 22556
rect 25648 22516 25654 22528
rect 25777 22525 25789 22528
rect 25823 22525 25835 22559
rect 25777 22519 25835 22525
rect 19334 22448 19340 22500
rect 19392 22488 19398 22500
rect 19797 22491 19855 22497
rect 19797 22488 19809 22491
rect 19392 22460 19809 22488
rect 19392 22448 19398 22460
rect 19797 22457 19809 22460
rect 19843 22457 19855 22491
rect 19797 22451 19855 22457
rect 20806 22448 20812 22500
rect 20864 22488 20870 22500
rect 24670 22488 24676 22500
rect 20864 22460 24676 22488
rect 20864 22448 20870 22460
rect 24670 22448 24676 22460
rect 24728 22448 24734 22500
rect 19613 22423 19671 22429
rect 19613 22420 19625 22423
rect 17972 22392 19625 22420
rect 17405 22383 17463 22389
rect 19613 22389 19625 22392
rect 19659 22420 19671 22423
rect 20254 22420 20260 22432
rect 19659 22392 20260 22420
rect 19659 22389 19671 22392
rect 19613 22383 19671 22389
rect 20254 22380 20260 22392
rect 20312 22380 20318 22432
rect 24854 22380 24860 22432
rect 24912 22420 24918 22432
rect 26145 22423 26203 22429
rect 26145 22420 26157 22423
rect 24912 22392 26157 22420
rect 24912 22380 24918 22392
rect 26145 22389 26157 22392
rect 26191 22389 26203 22423
rect 26145 22383 26203 22389
rect 41966 22380 41972 22432
rect 42024 22420 42030 22432
rect 58253 22423 58311 22429
rect 58253 22420 58265 22423
rect 42024 22392 58265 22420
rect 42024 22380 42030 22392
rect 58253 22389 58265 22392
rect 58299 22389 58311 22423
rect 58253 22383 58311 22389
rect 1104 22330 58880 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 58880 22330
rect 1104 22256 58880 22278
rect 9674 22216 9680 22228
rect 9635 22188 9680 22216
rect 9674 22176 9680 22188
rect 9732 22176 9738 22228
rect 20990 22148 20996 22160
rect 19306 22120 20996 22148
rect 10134 22080 10140 22092
rect 9508 22052 10140 22080
rect 1581 22015 1639 22021
rect 1581 21981 1593 22015
rect 1627 22012 1639 22015
rect 7282 22012 7288 22024
rect 1627 21984 7288 22012
rect 1627 21981 1639 21984
rect 1581 21975 1639 21981
rect 7282 21972 7288 21984
rect 7340 21972 7346 22024
rect 9508 22021 9536 22052
rect 10134 22040 10140 22052
rect 10192 22040 10198 22092
rect 9493 22015 9551 22021
rect 9493 21981 9505 22015
rect 9539 21981 9551 22015
rect 9493 21975 9551 21981
rect 9647 22015 9705 22021
rect 9647 21981 9659 22015
rect 9693 22012 9705 22015
rect 11054 22012 11060 22024
rect 9693 21984 11060 22012
rect 9693 21981 9705 21984
rect 9647 21975 9705 21981
rect 11054 21972 11060 21984
rect 11112 21972 11118 22024
rect 15930 21972 15936 22024
rect 15988 22012 15994 22024
rect 16577 22015 16635 22021
rect 16577 22012 16589 22015
rect 15988 21984 16589 22012
rect 15988 21972 15994 21984
rect 16577 21981 16589 21984
rect 16623 21981 16635 22015
rect 16577 21975 16635 21981
rect 17126 21972 17132 22024
rect 17184 22012 17190 22024
rect 19306 22012 19334 22120
rect 20990 22108 20996 22120
rect 21048 22108 21054 22160
rect 37274 22108 37280 22160
rect 37332 22148 37338 22160
rect 42426 22148 42432 22160
rect 37332 22120 42432 22148
rect 37332 22108 37338 22120
rect 42426 22108 42432 22120
rect 42484 22108 42490 22160
rect 26142 22080 26148 22092
rect 26103 22052 26148 22080
rect 26142 22040 26148 22052
rect 26200 22080 26206 22092
rect 31202 22080 31208 22092
rect 26200 22052 31208 22080
rect 26200 22040 26206 22052
rect 31202 22040 31208 22052
rect 31260 22040 31266 22092
rect 57330 22040 57336 22092
rect 57388 22080 57394 22092
rect 57698 22080 57704 22092
rect 57388 22052 57704 22080
rect 57388 22040 57394 22052
rect 57698 22040 57704 22052
rect 57756 22040 57762 22092
rect 20990 22012 20996 22024
rect 17184 21984 19334 22012
rect 20951 21984 20996 22012
rect 17184 21972 17190 21984
rect 20990 21972 20996 21984
rect 21048 21972 21054 22024
rect 21177 22015 21235 22021
rect 21177 21981 21189 22015
rect 21223 22012 21235 22015
rect 22002 22012 22008 22024
rect 21223 21984 22008 22012
rect 21223 21981 21235 21984
rect 21177 21975 21235 21981
rect 22002 21972 22008 21984
rect 22060 21972 22066 22024
rect 22094 21972 22100 22024
rect 22152 22012 22158 22024
rect 22830 22012 22836 22024
rect 22152 21984 22836 22012
rect 22152 21972 22158 21984
rect 22830 21972 22836 21984
rect 22888 21972 22894 22024
rect 57054 21972 57060 22024
rect 57112 22012 57118 22024
rect 57885 22015 57943 22021
rect 57885 22012 57897 22015
rect 57112 21984 57897 22012
rect 57112 21972 57118 21984
rect 57885 21981 57897 21984
rect 57931 21981 57943 22015
rect 57885 21975 57943 21981
rect 1854 21944 1860 21956
rect 1815 21916 1860 21944
rect 1854 21904 1860 21916
rect 1912 21904 1918 21956
rect 16390 21904 16396 21956
rect 16448 21944 16454 21956
rect 18138 21944 18144 21956
rect 16448 21916 18144 21944
rect 16448 21904 16454 21916
rect 18138 21904 18144 21916
rect 18196 21904 18202 21956
rect 19426 21904 19432 21956
rect 19484 21944 19490 21956
rect 19613 21947 19671 21953
rect 19613 21944 19625 21947
rect 19484 21916 19625 21944
rect 19484 21904 19490 21916
rect 19613 21913 19625 21916
rect 19659 21913 19671 21947
rect 19613 21907 19671 21913
rect 19702 21904 19708 21956
rect 19760 21944 19766 21956
rect 19889 21947 19947 21953
rect 19889 21944 19901 21947
rect 19760 21916 19901 21944
rect 19760 21904 19766 21916
rect 19889 21913 19901 21916
rect 19935 21913 19947 21947
rect 19889 21907 19947 21913
rect 19981 21947 20039 21953
rect 19981 21913 19993 21947
rect 20027 21944 20039 21947
rect 20254 21944 20260 21956
rect 20027 21916 20260 21944
rect 20027 21913 20039 21916
rect 19981 21907 20039 21913
rect 20254 21904 20260 21916
rect 20312 21944 20318 21956
rect 25038 21944 25044 21956
rect 20312 21916 25044 21944
rect 20312 21904 20318 21916
rect 25038 21904 25044 21916
rect 25096 21904 25102 21956
rect 28626 21904 28632 21956
rect 28684 21944 28690 21956
rect 35986 21944 35992 21956
rect 28684 21916 35992 21944
rect 28684 21904 28690 21916
rect 35986 21904 35992 21916
rect 36044 21904 36050 21956
rect 58158 21944 58164 21956
rect 58119 21916 58164 21944
rect 58158 21904 58164 21916
rect 58216 21904 58222 21956
rect 15378 21836 15384 21888
rect 15436 21876 15442 21888
rect 17773 21879 17831 21885
rect 17773 21876 17785 21879
rect 15436 21848 17785 21876
rect 15436 21836 15442 21848
rect 17773 21845 17785 21848
rect 17819 21845 17831 21879
rect 19794 21876 19800 21888
rect 19755 21848 19800 21876
rect 17773 21839 17831 21845
rect 19794 21836 19800 21848
rect 19852 21836 19858 21888
rect 20162 21876 20168 21888
rect 20123 21848 20168 21876
rect 20162 21836 20168 21848
rect 20220 21836 20226 21888
rect 21361 21879 21419 21885
rect 21361 21845 21373 21879
rect 21407 21876 21419 21879
rect 22094 21876 22100 21888
rect 21407 21848 22100 21876
rect 21407 21845 21419 21848
rect 21361 21839 21419 21845
rect 22094 21836 22100 21848
rect 22152 21836 22158 21888
rect 23842 21836 23848 21888
rect 23900 21876 23906 21888
rect 25593 21879 25651 21885
rect 25593 21876 25605 21879
rect 23900 21848 25605 21876
rect 23900 21836 23906 21848
rect 25593 21845 25605 21848
rect 25639 21845 25651 21879
rect 25593 21839 25651 21845
rect 25866 21836 25872 21888
rect 25924 21876 25930 21888
rect 25961 21879 26019 21885
rect 25961 21876 25973 21879
rect 25924 21848 25973 21876
rect 25924 21836 25930 21848
rect 25961 21845 25973 21848
rect 26007 21845 26019 21879
rect 25961 21839 26019 21845
rect 26053 21879 26111 21885
rect 26053 21845 26065 21879
rect 26099 21876 26111 21879
rect 28534 21876 28540 21888
rect 26099 21848 28540 21876
rect 26099 21845 26111 21848
rect 26053 21839 26111 21845
rect 28534 21836 28540 21848
rect 28592 21836 28598 21888
rect 35802 21836 35808 21888
rect 35860 21876 35866 21888
rect 58986 21876 58992 21888
rect 35860 21848 58992 21876
rect 35860 21836 35866 21848
rect 58986 21836 58992 21848
rect 59044 21836 59050 21888
rect 1104 21786 58880 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 58880 21786
rect 1104 21712 58880 21734
rect 7282 21632 7288 21684
rect 7340 21672 7346 21684
rect 12069 21675 12127 21681
rect 12069 21672 12081 21675
rect 7340 21644 12081 21672
rect 7340 21632 7346 21644
rect 12069 21641 12081 21644
rect 12115 21641 12127 21675
rect 12069 21635 12127 21641
rect 15838 21632 15844 21684
rect 15896 21672 15902 21684
rect 18322 21672 18328 21684
rect 15896 21644 18328 21672
rect 15896 21632 15902 21644
rect 18322 21632 18328 21644
rect 18380 21672 18386 21684
rect 19702 21672 19708 21684
rect 18380 21644 19708 21672
rect 18380 21632 18386 21644
rect 19702 21632 19708 21644
rect 19760 21632 19766 21684
rect 19978 21632 19984 21684
rect 20036 21672 20042 21684
rect 21450 21672 21456 21684
rect 20036 21644 21456 21672
rect 20036 21632 20042 21644
rect 21450 21632 21456 21644
rect 21508 21632 21514 21684
rect 22002 21672 22008 21684
rect 21963 21644 22008 21672
rect 22002 21632 22008 21644
rect 22060 21632 22066 21684
rect 22278 21632 22284 21684
rect 22336 21672 22342 21684
rect 22373 21675 22431 21681
rect 22373 21672 22385 21675
rect 22336 21644 22385 21672
rect 22336 21632 22342 21644
rect 22373 21641 22385 21644
rect 22419 21641 22431 21675
rect 22373 21635 22431 21641
rect 22462 21632 22468 21684
rect 22520 21672 22526 21684
rect 22738 21672 22744 21684
rect 22520 21644 22744 21672
rect 22520 21632 22526 21644
rect 22738 21632 22744 21644
rect 22796 21632 22802 21684
rect 24946 21672 24952 21684
rect 24907 21644 24952 21672
rect 24946 21632 24952 21644
rect 25004 21632 25010 21684
rect 25038 21632 25044 21684
rect 25096 21672 25102 21684
rect 29825 21675 29883 21681
rect 29825 21672 29837 21675
rect 25096 21644 29837 21672
rect 25096 21632 25102 21644
rect 29825 21641 29837 21644
rect 29871 21641 29883 21675
rect 57974 21672 57980 21684
rect 29825 21635 29883 21641
rect 29932 21644 57980 21672
rect 12406 21576 18920 21604
rect 1673 21539 1731 21545
rect 1673 21505 1685 21539
rect 1719 21536 1731 21539
rect 6822 21536 6828 21548
rect 1719 21508 6828 21536
rect 1719 21505 1731 21508
rect 1673 21499 1731 21505
rect 6822 21496 6828 21508
rect 6880 21496 6886 21548
rect 10318 21496 10324 21548
rect 10376 21536 10382 21548
rect 11701 21539 11759 21545
rect 11701 21536 11713 21539
rect 10376 21508 11713 21536
rect 10376 21496 10382 21508
rect 11701 21505 11713 21508
rect 11747 21505 11759 21539
rect 11701 21499 11759 21505
rect 11855 21539 11913 21545
rect 11855 21505 11867 21539
rect 11901 21536 11913 21539
rect 12406 21536 12434 21576
rect 11901 21508 12434 21536
rect 11901 21505 11913 21508
rect 11855 21499 11913 21505
rect 12710 21496 12716 21548
rect 12768 21536 12774 21548
rect 12989 21539 13047 21545
rect 12989 21536 13001 21539
rect 12768 21508 13001 21536
rect 12768 21496 12774 21508
rect 12989 21505 13001 21508
rect 13035 21505 13047 21539
rect 12989 21499 13047 21505
rect 13081 21539 13139 21545
rect 13081 21505 13093 21539
rect 13127 21505 13139 21539
rect 13262 21536 13268 21548
rect 13223 21508 13268 21536
rect 13081 21499 13139 21505
rect 12894 21428 12900 21480
rect 12952 21468 12958 21480
rect 13096 21468 13124 21499
rect 13262 21496 13268 21508
rect 13320 21496 13326 21548
rect 15203 21539 15261 21545
rect 15203 21505 15215 21539
rect 15249 21505 15261 21539
rect 15203 21499 15261 21505
rect 15381 21539 15439 21545
rect 15381 21505 15393 21539
rect 15427 21536 15439 21539
rect 16022 21536 16028 21548
rect 15427 21508 16028 21536
rect 15427 21505 15439 21508
rect 15381 21499 15439 21505
rect 12952 21440 13124 21468
rect 12952 21428 12958 21440
rect 13170 21428 13176 21480
rect 13228 21468 13234 21480
rect 15212 21468 15240 21499
rect 16022 21496 16028 21508
rect 16080 21496 16086 21548
rect 16117 21539 16175 21545
rect 16117 21505 16129 21539
rect 16163 21505 16175 21539
rect 16298 21536 16304 21548
rect 16259 21508 16304 21536
rect 16117 21499 16175 21505
rect 16132 21468 16160 21499
rect 16298 21496 16304 21508
rect 16356 21496 16362 21548
rect 17212 21539 17270 21545
rect 17212 21505 17224 21539
rect 17258 21536 17270 21539
rect 18046 21536 18052 21548
rect 17258 21508 18052 21536
rect 17258 21505 17270 21508
rect 17212 21499 17270 21505
rect 18046 21496 18052 21508
rect 18104 21496 18110 21548
rect 18782 21536 18788 21548
rect 18743 21508 18788 21536
rect 18782 21496 18788 21508
rect 18840 21496 18846 21548
rect 18892 21536 18920 21576
rect 20070 21564 20076 21616
rect 20128 21604 20134 21616
rect 20806 21604 20812 21616
rect 20128 21576 20812 21604
rect 20128 21564 20134 21576
rect 20806 21564 20812 21576
rect 20864 21604 20870 21616
rect 20864 21576 23612 21604
rect 20864 21564 20870 21576
rect 23474 21536 23480 21548
rect 18892 21508 23480 21536
rect 23474 21496 23480 21508
rect 23532 21496 23538 21548
rect 23584 21545 23612 21576
rect 27522 21564 27528 21616
rect 27580 21604 27586 21616
rect 29932 21604 29960 21644
rect 57974 21632 57980 21644
rect 58032 21632 58038 21684
rect 27580 21576 29960 21604
rect 27580 21564 27586 21576
rect 30006 21564 30012 21616
rect 30064 21604 30070 21616
rect 38378 21604 38384 21616
rect 30064 21576 38384 21604
rect 30064 21564 30070 21576
rect 38378 21564 38384 21576
rect 38436 21564 38442 21616
rect 58250 21604 58256 21616
rect 38764 21576 58256 21604
rect 23569 21539 23627 21545
rect 23569 21505 23581 21539
rect 23615 21536 23627 21539
rect 27706 21536 27712 21548
rect 23615 21508 27712 21536
rect 23615 21505 23627 21508
rect 23569 21499 23627 21505
rect 27706 21496 27712 21508
rect 27764 21496 27770 21548
rect 27801 21539 27859 21545
rect 27801 21505 27813 21539
rect 27847 21536 27859 21539
rect 28626 21536 28632 21548
rect 27847 21508 28488 21536
rect 28587 21508 28632 21536
rect 27847 21505 27859 21508
rect 27801 21499 27859 21505
rect 16574 21468 16580 21480
rect 13228 21440 13273 21468
rect 15212 21440 15332 21468
rect 16132 21440 16580 21468
rect 13228 21428 13234 21440
rect 15304 21400 15332 21440
rect 16574 21428 16580 21440
rect 16632 21428 16638 21480
rect 16850 21428 16856 21480
rect 16908 21468 16914 21480
rect 16945 21471 17003 21477
rect 16945 21468 16957 21471
rect 16908 21440 16957 21468
rect 16908 21428 16914 21440
rect 16945 21437 16957 21440
rect 16991 21437 17003 21471
rect 16945 21431 17003 21437
rect 22465 21471 22523 21477
rect 22465 21437 22477 21471
rect 22511 21437 22523 21471
rect 22465 21431 22523 21437
rect 22649 21471 22707 21477
rect 22649 21437 22661 21471
rect 22695 21468 22707 21471
rect 25038 21468 25044 21480
rect 22695 21440 25044 21468
rect 22695 21437 22707 21440
rect 22649 21431 22707 21437
rect 18325 21403 18383 21409
rect 15304 21372 16252 21400
rect 1762 21332 1768 21344
rect 1723 21304 1768 21332
rect 1762 21292 1768 21304
rect 1820 21292 1826 21344
rect 12802 21332 12808 21344
rect 12763 21304 12808 21332
rect 12802 21292 12808 21304
rect 12860 21292 12866 21344
rect 15197 21335 15255 21341
rect 15197 21301 15209 21335
rect 15243 21332 15255 21335
rect 15286 21332 15292 21344
rect 15243 21304 15292 21332
rect 15243 21301 15255 21304
rect 15197 21295 15255 21301
rect 15286 21292 15292 21304
rect 15344 21292 15350 21344
rect 16114 21332 16120 21344
rect 16075 21304 16120 21332
rect 16114 21292 16120 21304
rect 16172 21292 16178 21344
rect 16224 21332 16252 21372
rect 18325 21369 18337 21403
rect 18371 21400 18383 21403
rect 22278 21400 22284 21412
rect 18371 21372 22284 21400
rect 18371 21369 18383 21372
rect 18325 21363 18383 21369
rect 22278 21360 22284 21372
rect 22336 21360 22342 21412
rect 22370 21360 22376 21412
rect 22428 21400 22434 21412
rect 22480 21400 22508 21431
rect 25038 21428 25044 21440
rect 25096 21468 25102 21480
rect 26142 21468 26148 21480
rect 25096 21440 26148 21468
rect 25096 21428 25102 21440
rect 26142 21428 26148 21440
rect 26200 21428 26206 21480
rect 27890 21468 27896 21480
rect 27851 21440 27896 21468
rect 27890 21428 27896 21440
rect 27948 21428 27954 21480
rect 27982 21428 27988 21480
rect 28040 21468 28046 21480
rect 28460 21468 28488 21508
rect 28626 21496 28632 21508
rect 28684 21496 28690 21548
rect 35894 21496 35900 21548
rect 35952 21536 35958 21548
rect 35989 21539 36047 21545
rect 35989 21536 36001 21539
rect 35952 21508 36001 21536
rect 35952 21496 35958 21508
rect 35989 21505 36001 21508
rect 36035 21505 36047 21539
rect 35989 21499 36047 21505
rect 38194 21496 38200 21548
rect 38252 21536 38258 21548
rect 38657 21539 38715 21545
rect 38657 21536 38669 21539
rect 38252 21508 38669 21536
rect 38252 21496 38258 21508
rect 38657 21505 38669 21508
rect 38703 21505 38715 21539
rect 38657 21499 38715 21505
rect 28810 21468 28816 21480
rect 28040 21440 28085 21468
rect 28460 21440 28816 21468
rect 28040 21428 28046 21440
rect 28810 21428 28816 21440
rect 28868 21428 28874 21480
rect 35802 21468 35808 21480
rect 35268 21440 35808 21468
rect 22428 21372 22508 21400
rect 22428 21360 22434 21372
rect 23014 21360 23020 21412
rect 23072 21400 23078 21412
rect 25590 21400 25596 21412
rect 23072 21372 25596 21400
rect 23072 21360 23078 21372
rect 25590 21360 25596 21372
rect 25648 21360 25654 21412
rect 28258 21400 28264 21412
rect 26344 21372 28264 21400
rect 17310 21332 17316 21344
rect 16224 21304 17316 21332
rect 17310 21292 17316 21304
rect 17368 21292 17374 21344
rect 19978 21332 19984 21344
rect 19939 21304 19984 21332
rect 19978 21292 19984 21304
rect 20036 21292 20042 21344
rect 20070 21292 20076 21344
rect 20128 21332 20134 21344
rect 26344 21332 26372 21372
rect 28258 21360 28264 21372
rect 28316 21360 28322 21412
rect 20128 21304 26372 21332
rect 27433 21335 27491 21341
rect 20128 21292 20134 21304
rect 27433 21301 27445 21335
rect 27479 21332 27491 21335
rect 28350 21332 28356 21344
rect 27479 21304 28356 21332
rect 27479 21301 27491 21304
rect 27433 21295 27491 21301
rect 28350 21292 28356 21304
rect 28408 21292 28414 21344
rect 28537 21335 28595 21341
rect 28537 21301 28549 21335
rect 28583 21332 28595 21335
rect 28718 21332 28724 21344
rect 28583 21304 28724 21332
rect 28583 21301 28595 21304
rect 28537 21295 28595 21301
rect 28718 21292 28724 21304
rect 28776 21292 28782 21344
rect 34698 21292 34704 21344
rect 34756 21332 34762 21344
rect 35268 21341 35296 21440
rect 35802 21428 35808 21440
rect 35860 21468 35866 21480
rect 36081 21471 36139 21477
rect 36081 21468 36093 21471
rect 35860 21440 36093 21468
rect 35860 21428 35866 21440
rect 36081 21437 36093 21440
rect 36127 21437 36139 21471
rect 36081 21431 36139 21437
rect 36265 21471 36323 21477
rect 36265 21437 36277 21471
rect 36311 21468 36323 21471
rect 36630 21468 36636 21480
rect 36311 21440 36636 21468
rect 36311 21437 36323 21440
rect 36265 21431 36323 21437
rect 36630 21428 36636 21440
rect 36688 21428 36694 21480
rect 38764 21477 38792 21576
rect 58250 21564 58256 21576
rect 58308 21564 58314 21616
rect 58066 21536 58072 21548
rect 58027 21508 58072 21536
rect 58066 21496 58072 21508
rect 58124 21496 58130 21548
rect 38749 21471 38807 21477
rect 38749 21468 38761 21471
rect 37936 21440 38761 21468
rect 35253 21335 35311 21341
rect 35253 21332 35265 21335
rect 34756 21304 35265 21332
rect 34756 21292 34762 21304
rect 35253 21301 35265 21304
rect 35299 21301 35311 21335
rect 35618 21332 35624 21344
rect 35579 21304 35624 21332
rect 35253 21295 35311 21301
rect 35618 21292 35624 21304
rect 35676 21292 35682 21344
rect 35710 21292 35716 21344
rect 35768 21332 35774 21344
rect 37936 21341 37964 21440
rect 38749 21437 38761 21440
rect 38795 21437 38807 21471
rect 38749 21431 38807 21437
rect 38838 21428 38844 21480
rect 38896 21468 38902 21480
rect 41690 21468 41696 21480
rect 38896 21440 41696 21468
rect 38896 21428 38902 21440
rect 41690 21428 41696 21440
rect 41748 21428 41754 21480
rect 38378 21360 38384 21412
rect 38436 21400 38442 21412
rect 52730 21400 52736 21412
rect 38436 21372 52736 21400
rect 38436 21360 38442 21372
rect 52730 21360 52736 21372
rect 52788 21360 52794 21412
rect 53190 21360 53196 21412
rect 53248 21400 53254 21412
rect 58158 21400 58164 21412
rect 53248 21372 58164 21400
rect 53248 21360 53254 21372
rect 58158 21360 58164 21372
rect 58216 21360 58222 21412
rect 37921 21335 37979 21341
rect 37921 21332 37933 21335
rect 35768 21304 37933 21332
rect 35768 21292 35774 21304
rect 37921 21301 37933 21304
rect 37967 21301 37979 21335
rect 37921 21295 37979 21301
rect 38289 21335 38347 21341
rect 38289 21301 38301 21335
rect 38335 21332 38347 21335
rect 38470 21332 38476 21344
rect 38335 21304 38476 21332
rect 38335 21301 38347 21304
rect 38289 21295 38347 21301
rect 38470 21292 38476 21304
rect 38528 21292 38534 21344
rect 50982 21292 50988 21344
rect 51040 21332 51046 21344
rect 52086 21332 52092 21344
rect 51040 21304 52092 21332
rect 51040 21292 51046 21304
rect 52086 21292 52092 21304
rect 52144 21292 52150 21344
rect 58250 21332 58256 21344
rect 58211 21304 58256 21332
rect 58250 21292 58256 21304
rect 58308 21292 58314 21344
rect 1104 21242 58880 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 58880 21242
rect 1104 21168 58880 21190
rect 15930 21128 15936 21140
rect 15891 21100 15936 21128
rect 15930 21088 15936 21100
rect 15988 21088 15994 21140
rect 16022 21088 16028 21140
rect 16080 21128 16086 21140
rect 19981 21131 20039 21137
rect 19981 21128 19993 21131
rect 16080 21100 19993 21128
rect 16080 21088 16086 21100
rect 19981 21097 19993 21100
rect 20027 21097 20039 21131
rect 27614 21128 27620 21140
rect 19981 21091 20039 21097
rect 22066 21100 27620 21128
rect 12710 21060 12716 21072
rect 11716 21032 12716 21060
rect 11716 21004 11744 21032
rect 12710 21020 12716 21032
rect 12768 21060 12774 21072
rect 16040 21060 16068 21088
rect 12768 21032 16068 21060
rect 12768 21020 12774 21032
rect 11698 20992 11704 21004
rect 11659 20964 11704 20992
rect 11698 20952 11704 20964
rect 11756 20952 11762 21004
rect 12161 20995 12219 21001
rect 12161 20961 12173 20995
rect 12207 20992 12219 20995
rect 12250 20992 12256 21004
rect 12207 20964 12256 20992
rect 12207 20961 12219 20964
rect 12161 20955 12219 20961
rect 12250 20952 12256 20964
rect 12308 20952 12314 21004
rect 13170 20992 13176 21004
rect 12820 20964 13176 20992
rect 11793 20927 11851 20933
rect 11793 20893 11805 20927
rect 11839 20893 11851 20927
rect 11793 20887 11851 20893
rect 11146 20748 11152 20800
rect 11204 20788 11210 20800
rect 11808 20788 11836 20887
rect 12710 20884 12716 20936
rect 12768 20924 12774 20936
rect 12820 20933 12848 20964
rect 13170 20952 13176 20964
rect 13228 20992 13234 21004
rect 13630 20992 13636 21004
rect 13228 20964 13636 20992
rect 13228 20952 13234 20964
rect 13630 20952 13636 20964
rect 13688 20952 13694 21004
rect 12805 20927 12863 20933
rect 12805 20924 12817 20927
rect 12768 20896 12817 20924
rect 12768 20884 12774 20896
rect 12805 20893 12817 20896
rect 12851 20893 12863 20927
rect 12805 20887 12863 20893
rect 12989 20927 13047 20933
rect 12989 20893 13001 20927
rect 13035 20924 13047 20927
rect 13740 20924 13768 21032
rect 16298 21020 16304 21072
rect 16356 21060 16362 21072
rect 19429 21063 19487 21069
rect 19429 21060 19441 21063
rect 16356 21032 19441 21060
rect 16356 21020 16362 21032
rect 19429 21029 19441 21032
rect 19475 21060 19487 21063
rect 22066 21060 22094 21100
rect 27614 21088 27620 21100
rect 27672 21088 27678 21140
rect 27890 21088 27896 21140
rect 27948 21128 27954 21140
rect 28718 21128 28724 21140
rect 27948 21100 28724 21128
rect 27948 21088 27954 21100
rect 28718 21088 28724 21100
rect 28776 21128 28782 21140
rect 28776 21100 31754 21128
rect 28776 21088 28782 21100
rect 19475 21032 22094 21060
rect 27341 21063 27399 21069
rect 19475 21029 19487 21032
rect 19429 21023 19487 21029
rect 27341 21029 27353 21063
rect 27387 21029 27399 21063
rect 27341 21023 27399 21029
rect 30653 21063 30711 21069
rect 30653 21029 30665 21063
rect 30699 21029 30711 21063
rect 31726 21060 31754 21100
rect 32490 21088 32496 21140
rect 32548 21128 32554 21140
rect 58250 21128 58256 21140
rect 32548 21100 58256 21128
rect 32548 21088 32554 21100
rect 58250 21088 58256 21100
rect 58308 21088 58314 21140
rect 53190 21060 53196 21072
rect 31726 21032 53196 21060
rect 30653 21023 30711 21029
rect 16666 20992 16672 21004
rect 15488 20964 16672 20992
rect 13035 20896 13768 20924
rect 15289 20927 15347 20933
rect 13035 20893 13047 20896
rect 12989 20887 13047 20893
rect 15289 20893 15301 20927
rect 15335 20924 15347 20927
rect 15378 20924 15384 20936
rect 15335 20896 15384 20924
rect 15335 20893 15347 20896
rect 15289 20887 15347 20893
rect 15378 20884 15384 20896
rect 15436 20884 15442 20936
rect 15488 20933 15516 20964
rect 16666 20952 16672 20964
rect 16724 20952 16730 21004
rect 17954 20992 17960 21004
rect 17915 20964 17960 20992
rect 17954 20952 17960 20964
rect 18012 20952 18018 21004
rect 19518 20952 19524 21004
rect 19576 20992 19582 21004
rect 22005 20995 22063 21001
rect 22005 20992 22017 20995
rect 19576 20964 22017 20992
rect 19576 20952 19582 20964
rect 22005 20961 22017 20964
rect 22051 20961 22063 20995
rect 22005 20955 22063 20961
rect 15473 20927 15531 20933
rect 15473 20893 15485 20927
rect 15519 20893 15531 20927
rect 15473 20887 15531 20893
rect 15562 20884 15568 20936
rect 15620 20924 15626 20936
rect 15838 20924 15844 20936
rect 15620 20896 15844 20924
rect 15620 20884 15626 20896
rect 15838 20884 15844 20896
rect 15896 20924 15902 20936
rect 15933 20927 15991 20933
rect 15933 20924 15945 20927
rect 15896 20896 15945 20924
rect 15896 20884 15902 20896
rect 15933 20893 15945 20896
rect 15979 20893 15991 20927
rect 15933 20887 15991 20893
rect 16022 20884 16028 20936
rect 16080 20924 16086 20936
rect 16117 20927 16175 20933
rect 16117 20924 16129 20927
rect 16080 20896 16129 20924
rect 16080 20884 16086 20896
rect 16117 20893 16129 20896
rect 16163 20924 16175 20927
rect 16390 20924 16396 20936
rect 16163 20896 16396 20924
rect 16163 20893 16175 20896
rect 16117 20887 16175 20893
rect 16390 20884 16396 20896
rect 16448 20884 16454 20936
rect 16577 20927 16635 20933
rect 16577 20893 16589 20927
rect 16623 20924 16635 20927
rect 16758 20924 16764 20936
rect 16623 20896 16764 20924
rect 16623 20893 16635 20896
rect 16577 20887 16635 20893
rect 16758 20884 16764 20896
rect 16816 20884 16822 20936
rect 17218 20884 17224 20936
rect 17276 20924 17282 20936
rect 19797 20927 19855 20933
rect 19797 20924 19809 20927
rect 17276 20896 19809 20924
rect 17276 20884 17282 20896
rect 19797 20893 19809 20896
rect 19843 20924 19855 20927
rect 20162 20924 20168 20936
rect 19843 20896 20168 20924
rect 19843 20893 19855 20896
rect 19797 20887 19855 20893
rect 20162 20884 20168 20896
rect 20220 20884 20226 20936
rect 20901 20927 20959 20933
rect 20901 20893 20913 20927
rect 20947 20924 20959 20927
rect 22738 20924 22744 20936
rect 20947 20896 22744 20924
rect 20947 20893 20959 20896
rect 20901 20887 20959 20893
rect 22738 20884 22744 20896
rect 22796 20884 22802 20936
rect 23014 20884 23020 20936
rect 23072 20924 23078 20936
rect 23661 20927 23719 20933
rect 23661 20924 23673 20927
rect 23072 20896 23673 20924
rect 23072 20884 23078 20896
rect 23661 20893 23673 20896
rect 23707 20893 23719 20927
rect 23842 20924 23848 20936
rect 23803 20896 23848 20924
rect 23661 20887 23719 20893
rect 23842 20884 23848 20896
rect 23900 20884 23906 20936
rect 24581 20927 24639 20933
rect 24581 20893 24593 20927
rect 24627 20924 24639 20927
rect 26234 20924 26240 20936
rect 24627 20896 26240 20924
rect 24627 20893 24639 20896
rect 24581 20887 24639 20893
rect 26234 20884 26240 20896
rect 26292 20884 26298 20936
rect 26421 20927 26479 20933
rect 26421 20893 26433 20927
rect 26467 20893 26479 20927
rect 26421 20887 26479 20893
rect 26513 20927 26571 20933
rect 26513 20893 26525 20927
rect 26559 20924 26571 20927
rect 27356 20924 27384 21023
rect 27522 20952 27528 21004
rect 27580 20992 27586 21004
rect 27801 20995 27859 21001
rect 27801 20992 27813 20995
rect 27580 20964 27813 20992
rect 27580 20952 27586 20964
rect 27801 20961 27813 20964
rect 27847 20961 27859 20995
rect 27982 20992 27988 21004
rect 27943 20964 27988 20992
rect 27801 20955 27859 20961
rect 27982 20952 27988 20964
rect 28040 20952 28046 21004
rect 28350 20952 28356 21004
rect 28408 20992 28414 21004
rect 28408 20964 28764 20992
rect 28408 20952 28414 20964
rect 26559 20896 27384 20924
rect 26559 20893 26571 20896
rect 26513 20887 26571 20893
rect 12621 20859 12679 20865
rect 12621 20825 12633 20859
rect 12667 20856 12679 20859
rect 13262 20856 13268 20868
rect 12667 20828 13268 20856
rect 12667 20825 12679 20828
rect 12621 20819 12679 20825
rect 13262 20816 13268 20828
rect 13320 20856 13326 20868
rect 19334 20856 19340 20868
rect 13320 20828 15516 20856
rect 13320 20816 13326 20828
rect 12894 20788 12900 20800
rect 11204 20760 12900 20788
rect 11204 20748 11210 20760
rect 12894 20748 12900 20760
rect 12952 20748 12958 20800
rect 13078 20748 13084 20800
rect 13136 20788 13142 20800
rect 13173 20791 13231 20797
rect 13173 20788 13185 20791
rect 13136 20760 13185 20788
rect 13136 20748 13142 20760
rect 13173 20757 13185 20760
rect 13219 20757 13231 20791
rect 15378 20788 15384 20800
rect 15339 20760 15384 20788
rect 13173 20751 13231 20757
rect 15378 20748 15384 20760
rect 15436 20748 15442 20800
rect 15488 20788 15516 20828
rect 17880 20828 19340 20856
rect 17880 20788 17908 20828
rect 19334 20816 19340 20828
rect 19392 20816 19398 20868
rect 20070 20856 20076 20868
rect 19628 20828 20076 20856
rect 15488 20760 17908 20788
rect 18138 20748 18144 20800
rect 18196 20788 18202 20800
rect 19628 20797 19656 20828
rect 20070 20816 20076 20828
rect 20128 20816 20134 20868
rect 24029 20859 24087 20865
rect 24029 20825 24041 20859
rect 24075 20856 24087 20859
rect 24826 20859 24884 20865
rect 24826 20856 24838 20859
rect 24075 20828 24838 20856
rect 24075 20825 24087 20828
rect 24029 20819 24087 20825
rect 24826 20825 24838 20828
rect 24872 20825 24884 20859
rect 26436 20856 26464 20887
rect 26436 20828 26924 20856
rect 24826 20819 24884 20825
rect 19613 20791 19671 20797
rect 19613 20788 19625 20791
rect 18196 20760 19625 20788
rect 18196 20748 18202 20760
rect 19613 20757 19625 20760
rect 19659 20757 19671 20791
rect 19613 20751 19671 20757
rect 19702 20748 19708 20800
rect 19760 20788 19766 20800
rect 20254 20788 20260 20800
rect 19760 20760 20260 20788
rect 19760 20748 19766 20760
rect 20254 20748 20260 20760
rect 20312 20748 20318 20800
rect 23474 20748 23480 20800
rect 23532 20788 23538 20800
rect 25222 20788 25228 20800
rect 23532 20760 25228 20788
rect 23532 20748 23538 20760
rect 25222 20748 25228 20760
rect 25280 20748 25286 20800
rect 25958 20788 25964 20800
rect 25919 20760 25964 20788
rect 25958 20748 25964 20760
rect 26016 20748 26022 20800
rect 26694 20788 26700 20800
rect 26655 20760 26700 20788
rect 26694 20748 26700 20760
rect 26752 20748 26758 20800
rect 26896 20788 26924 20828
rect 26970 20816 26976 20868
rect 27028 20856 27034 20868
rect 27065 20859 27123 20865
rect 27065 20856 27077 20859
rect 27028 20828 27077 20856
rect 27028 20816 27034 20828
rect 27065 20825 27077 20828
rect 27111 20856 27123 20859
rect 27540 20856 27568 20952
rect 27706 20924 27712 20936
rect 27667 20896 27712 20924
rect 27706 20884 27712 20896
rect 27764 20884 27770 20936
rect 28736 20933 28764 20964
rect 28629 20927 28687 20933
rect 28629 20893 28641 20927
rect 28675 20893 28687 20927
rect 28629 20887 28687 20893
rect 28721 20927 28779 20933
rect 28721 20893 28733 20927
rect 28767 20893 28779 20927
rect 28721 20887 28779 20893
rect 27111 20828 27568 20856
rect 28644 20856 28672 20887
rect 29730 20884 29736 20936
rect 29788 20924 29794 20936
rect 29825 20927 29883 20933
rect 29825 20924 29837 20927
rect 29788 20896 29837 20924
rect 29788 20884 29794 20896
rect 29825 20893 29837 20896
rect 29871 20893 29883 20927
rect 29825 20887 29883 20893
rect 30009 20927 30067 20933
rect 30009 20893 30021 20927
rect 30055 20924 30067 20927
rect 30668 20924 30696 21023
rect 53190 21020 53196 21032
rect 53248 21020 53254 21072
rect 53285 21063 53343 21069
rect 53285 21029 53297 21063
rect 53331 21060 53343 21063
rect 53331 21032 53972 21060
rect 53331 21029 53343 21032
rect 53285 21023 53343 21029
rect 30742 20952 30748 21004
rect 30800 20992 30806 21004
rect 31202 20992 31208 21004
rect 30800 20964 31208 20992
rect 30800 20952 30806 20964
rect 31202 20952 31208 20964
rect 31260 20952 31266 21004
rect 35986 20992 35992 21004
rect 35947 20964 35992 20992
rect 35986 20952 35992 20964
rect 36044 20952 36050 21004
rect 37274 20952 37280 21004
rect 37332 20992 37338 21004
rect 38289 20995 38347 21001
rect 38289 20992 38301 20995
rect 37332 20964 38301 20992
rect 37332 20952 37338 20964
rect 38289 20961 38301 20964
rect 38335 20961 38347 20995
rect 38289 20955 38347 20961
rect 41690 20952 41696 21004
rect 41748 20992 41754 21004
rect 42061 20995 42119 21001
rect 42061 20992 42073 20995
rect 41748 20964 42073 20992
rect 41748 20952 41754 20964
rect 42061 20961 42073 20964
rect 42107 20961 42119 20995
rect 42061 20955 42119 20961
rect 52086 20952 52092 21004
rect 52144 20992 52150 21004
rect 52144 20964 53788 20992
rect 52144 20952 52150 20964
rect 34882 20924 34888 20936
rect 30055 20896 30696 20924
rect 34843 20896 34888 20924
rect 30055 20893 30067 20896
rect 30009 20887 30067 20893
rect 34882 20884 34888 20896
rect 34940 20924 34946 20936
rect 38194 20924 38200 20936
rect 34940 20896 38200 20924
rect 34940 20884 34946 20896
rect 38194 20884 38200 20896
rect 38252 20884 38258 20936
rect 38470 20924 38476 20936
rect 38431 20896 38476 20924
rect 38470 20884 38476 20896
rect 38528 20884 38534 20936
rect 41138 20884 41144 20936
rect 41196 20924 41202 20936
rect 42705 20927 42763 20933
rect 42705 20924 42717 20927
rect 41196 20896 42717 20924
rect 41196 20884 41202 20896
rect 42705 20893 42717 20896
rect 42751 20893 42763 20927
rect 42886 20924 42892 20936
rect 42847 20896 42892 20924
rect 42705 20887 42763 20893
rect 42886 20884 42892 20896
rect 42944 20884 42950 20936
rect 42978 20884 42984 20936
rect 43036 20924 43042 20936
rect 43901 20927 43959 20933
rect 43901 20924 43913 20927
rect 43036 20896 43913 20924
rect 43036 20884 43042 20896
rect 43901 20893 43913 20896
rect 43947 20893 43959 20927
rect 43901 20887 43959 20893
rect 44358 20884 44364 20936
rect 44416 20924 44422 20936
rect 47489 20927 47547 20933
rect 47489 20924 47501 20927
rect 44416 20896 47501 20924
rect 44416 20884 44422 20896
rect 47489 20893 47501 20896
rect 47535 20893 47547 20927
rect 47854 20924 47860 20936
rect 47815 20896 47860 20924
rect 47489 20887 47547 20893
rect 47854 20884 47860 20896
rect 47912 20884 47918 20936
rect 52730 20924 52736 20936
rect 52691 20896 52736 20924
rect 52730 20884 52736 20896
rect 52788 20884 52794 20936
rect 53098 20924 53104 20936
rect 52840 20896 53104 20924
rect 29748 20856 29776 20884
rect 28644 20828 29776 20856
rect 27111 20825 27123 20828
rect 27065 20819 27123 20825
rect 36630 20816 36636 20868
rect 36688 20856 36694 20868
rect 38838 20856 38844 20868
rect 36688 20828 38844 20856
rect 36688 20816 36694 20828
rect 38838 20816 38844 20828
rect 38896 20816 38902 20868
rect 41877 20859 41935 20865
rect 41877 20825 41889 20859
rect 41923 20856 41935 20859
rect 42518 20856 42524 20868
rect 41923 20828 42524 20856
rect 41923 20825 41935 20828
rect 41877 20819 41935 20825
rect 42518 20816 42524 20828
rect 42576 20856 42582 20868
rect 42576 20828 43208 20856
rect 42576 20816 42582 20828
rect 28442 20788 28448 20800
rect 26896 20760 28448 20788
rect 28442 20748 28448 20760
rect 28500 20748 28506 20800
rect 28902 20788 28908 20800
rect 28863 20760 28908 20788
rect 28902 20748 28908 20760
rect 28960 20748 28966 20800
rect 30193 20791 30251 20797
rect 30193 20757 30205 20791
rect 30239 20788 30251 20791
rect 30374 20788 30380 20800
rect 30239 20760 30380 20788
rect 30239 20757 30251 20760
rect 30193 20751 30251 20757
rect 30374 20748 30380 20760
rect 30432 20748 30438 20800
rect 31018 20788 31024 20800
rect 30979 20760 31024 20788
rect 31018 20748 31024 20760
rect 31076 20748 31082 20800
rect 31110 20748 31116 20800
rect 31168 20788 31174 20800
rect 31168 20760 31213 20788
rect 31168 20748 31174 20760
rect 31294 20748 31300 20800
rect 31352 20788 31358 20800
rect 32490 20788 32496 20800
rect 31352 20760 32496 20788
rect 31352 20748 31358 20760
rect 32490 20748 32496 20760
rect 32548 20748 32554 20800
rect 38654 20788 38660 20800
rect 38615 20760 38660 20788
rect 38654 20748 38660 20760
rect 38712 20748 38718 20800
rect 41414 20748 41420 20800
rect 41472 20788 41478 20800
rect 41509 20791 41567 20797
rect 41509 20788 41521 20791
rect 41472 20760 41521 20788
rect 41472 20748 41478 20760
rect 41509 20757 41521 20760
rect 41555 20757 41567 20791
rect 41509 20751 41567 20757
rect 41966 20748 41972 20800
rect 42024 20788 42030 20800
rect 43070 20788 43076 20800
rect 42024 20760 42069 20788
rect 43031 20760 43076 20788
rect 42024 20748 42030 20760
rect 43070 20748 43076 20760
rect 43128 20748 43134 20800
rect 43180 20788 43208 20828
rect 43438 20816 43444 20868
rect 43496 20856 43502 20868
rect 43533 20859 43591 20865
rect 43533 20856 43545 20859
rect 43496 20828 43545 20856
rect 43496 20816 43502 20828
rect 43533 20825 43545 20828
rect 43579 20825 43591 20859
rect 43533 20819 43591 20825
rect 43717 20859 43775 20865
rect 43717 20825 43729 20859
rect 43763 20825 43775 20859
rect 47670 20856 47676 20868
rect 47631 20828 47676 20856
rect 43717 20819 43775 20825
rect 43732 20788 43760 20819
rect 47670 20816 47676 20828
rect 47728 20816 47734 20868
rect 47765 20859 47823 20865
rect 47765 20825 47777 20859
rect 47811 20856 47823 20859
rect 49142 20856 49148 20868
rect 47811 20828 49148 20856
rect 47811 20825 47823 20828
rect 47765 20819 47823 20825
rect 49142 20816 49148 20828
rect 49200 20816 49206 20868
rect 50706 20816 50712 20868
rect 50764 20856 50770 20868
rect 52840 20856 52868 20896
rect 53098 20884 53104 20896
rect 53156 20884 53162 20936
rect 53760 20933 53788 20964
rect 53944 20933 53972 21032
rect 54110 20992 54116 21004
rect 54071 20964 54116 20992
rect 54110 20952 54116 20964
rect 54168 20952 54174 21004
rect 54573 20995 54631 21001
rect 54573 20961 54585 20995
rect 54619 20992 54631 20995
rect 55306 20992 55312 21004
rect 54619 20964 55312 20992
rect 54619 20961 54631 20964
rect 54573 20955 54631 20961
rect 55306 20952 55312 20964
rect 55364 20992 55370 21004
rect 55585 20995 55643 21001
rect 55585 20992 55597 20995
rect 55364 20964 55597 20992
rect 55364 20952 55370 20964
rect 55585 20961 55597 20964
rect 55631 20961 55643 20995
rect 55585 20955 55643 20961
rect 55692 20964 57928 20992
rect 53745 20927 53803 20933
rect 53745 20893 53757 20927
rect 53791 20893 53803 20927
rect 53745 20887 53803 20893
rect 53929 20927 53987 20933
rect 53929 20893 53941 20927
rect 53975 20893 53987 20927
rect 54478 20924 54484 20936
rect 53929 20887 53987 20893
rect 54036 20896 54484 20924
rect 50764 20828 52868 20856
rect 52917 20859 52975 20865
rect 50764 20816 50770 20828
rect 52917 20825 52929 20859
rect 52963 20825 52975 20859
rect 52917 20819 52975 20825
rect 53009 20859 53067 20865
rect 53009 20825 53021 20859
rect 53055 20856 53067 20859
rect 54036 20856 54064 20896
rect 54478 20884 54484 20896
rect 54536 20884 54542 20936
rect 54754 20924 54760 20936
rect 54715 20896 54760 20924
rect 54754 20884 54760 20896
rect 54812 20884 54818 20936
rect 54846 20884 54852 20936
rect 54904 20924 54910 20936
rect 55692 20924 55720 20964
rect 54904 20896 55720 20924
rect 55769 20927 55827 20933
rect 54904 20884 54910 20896
rect 55769 20893 55781 20927
rect 55815 20924 55827 20927
rect 56042 20924 56048 20936
rect 55815 20896 56048 20924
rect 55815 20893 55827 20896
rect 55769 20887 55827 20893
rect 56042 20884 56048 20896
rect 56100 20884 56106 20936
rect 57900 20933 57928 20964
rect 57885 20927 57943 20933
rect 57885 20893 57897 20927
rect 57931 20893 57943 20927
rect 57885 20887 57943 20893
rect 55674 20856 55680 20868
rect 53055 20828 54064 20856
rect 54588 20828 55680 20856
rect 53055 20825 53067 20828
rect 53009 20819 53067 20825
rect 43180 20760 43760 20788
rect 48041 20791 48099 20797
rect 48041 20757 48053 20791
rect 48087 20788 48099 20791
rect 48222 20788 48228 20800
rect 48087 20760 48228 20788
rect 48087 20757 48099 20760
rect 48041 20751 48099 20757
rect 48222 20748 48228 20760
rect 48280 20748 48286 20800
rect 52932 20788 52960 20819
rect 54588 20788 54616 20828
rect 55674 20816 55680 20828
rect 55732 20816 55738 20868
rect 58158 20856 58164 20868
rect 58119 20828 58164 20856
rect 58158 20816 58164 20828
rect 58216 20816 58222 20868
rect 52932 20760 54616 20788
rect 54941 20791 54999 20797
rect 54941 20757 54953 20791
rect 54987 20788 54999 20791
rect 55214 20788 55220 20800
rect 54987 20760 55220 20788
rect 54987 20757 54999 20760
rect 54941 20751 54999 20757
rect 55214 20748 55220 20760
rect 55272 20748 55278 20800
rect 55953 20791 56011 20797
rect 55953 20757 55965 20791
rect 55999 20788 56011 20791
rect 56686 20788 56692 20800
rect 55999 20760 56692 20788
rect 55999 20757 56011 20760
rect 55953 20751 56011 20757
rect 56686 20748 56692 20760
rect 56744 20748 56750 20800
rect 1104 20698 58880 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 58880 20698
rect 1104 20624 58880 20646
rect 12894 20544 12900 20596
rect 12952 20584 12958 20596
rect 18874 20584 18880 20596
rect 12952 20556 18880 20584
rect 12952 20544 12958 20556
rect 18874 20544 18880 20556
rect 18932 20544 18938 20596
rect 19334 20544 19340 20596
rect 19392 20584 19398 20596
rect 19705 20587 19763 20593
rect 19705 20584 19717 20587
rect 19392 20556 19717 20584
rect 19392 20544 19398 20556
rect 19705 20553 19717 20556
rect 19751 20553 19763 20587
rect 19705 20547 19763 20553
rect 19794 20544 19800 20596
rect 19852 20584 19858 20596
rect 25501 20587 25559 20593
rect 25501 20584 25513 20587
rect 19852 20556 25513 20584
rect 19852 20544 19858 20556
rect 25501 20553 25513 20556
rect 25547 20553 25559 20587
rect 25501 20547 25559 20553
rect 27706 20544 27712 20596
rect 27764 20584 27770 20596
rect 28166 20584 28172 20596
rect 27764 20556 28172 20584
rect 27764 20544 27770 20556
rect 28166 20544 28172 20556
rect 28224 20584 28230 20596
rect 28537 20587 28595 20593
rect 28537 20584 28549 20587
rect 28224 20556 28549 20584
rect 28224 20544 28230 20556
rect 28537 20553 28549 20556
rect 28583 20553 28595 20587
rect 28537 20547 28595 20553
rect 29472 20556 39344 20584
rect 11698 20516 11704 20528
rect 10980 20488 11704 20516
rect 1581 20451 1639 20457
rect 1581 20417 1593 20451
rect 1627 20448 1639 20451
rect 7374 20448 7380 20460
rect 1627 20420 7380 20448
rect 1627 20417 1639 20420
rect 1581 20411 1639 20417
rect 7374 20408 7380 20420
rect 7432 20408 7438 20460
rect 8018 20448 8024 20460
rect 7979 20420 8024 20448
rect 8018 20408 8024 20420
rect 8076 20408 8082 20460
rect 10980 20457 11008 20488
rect 11698 20476 11704 20488
rect 11756 20476 11762 20528
rect 13464 20488 18460 20516
rect 10965 20451 11023 20457
rect 10965 20417 10977 20451
rect 11011 20417 11023 20451
rect 11146 20448 11152 20460
rect 11107 20420 11152 20448
rect 10965 20411 11023 20417
rect 11146 20408 11152 20420
rect 11204 20408 11210 20460
rect 12428 20451 12486 20457
rect 12428 20417 12440 20451
rect 12474 20448 12486 20451
rect 13354 20448 13360 20460
rect 12474 20420 13360 20448
rect 12474 20417 12486 20420
rect 12428 20411 12486 20417
rect 13354 20408 13360 20420
rect 13412 20408 13418 20460
rect 1762 20380 1768 20392
rect 1723 20352 1768 20380
rect 1762 20340 1768 20352
rect 1820 20340 1826 20392
rect 11882 20340 11888 20392
rect 11940 20380 11946 20392
rect 12161 20383 12219 20389
rect 12161 20380 12173 20383
rect 11940 20352 12173 20380
rect 11940 20340 11946 20352
rect 12161 20349 12173 20352
rect 12207 20349 12219 20383
rect 12161 20343 12219 20349
rect 13464 20312 13492 20488
rect 14001 20451 14059 20457
rect 14001 20417 14013 20451
rect 14047 20448 14059 20451
rect 15378 20448 15384 20460
rect 14047 20420 15384 20448
rect 14047 20417 14059 20420
rect 14001 20411 14059 20417
rect 15378 20408 15384 20420
rect 15436 20408 15442 20460
rect 16666 20408 16672 20460
rect 16724 20448 16730 20460
rect 17589 20451 17647 20457
rect 17589 20448 17601 20451
rect 16724 20420 17601 20448
rect 16724 20408 16730 20420
rect 17589 20417 17601 20420
rect 17635 20417 17647 20451
rect 17862 20448 17868 20460
rect 17823 20420 17868 20448
rect 17589 20411 17647 20417
rect 17862 20408 17868 20420
rect 17920 20408 17926 20460
rect 18049 20451 18107 20457
rect 18049 20417 18061 20451
rect 18095 20417 18107 20451
rect 18432 20451 18460 20488
rect 22094 20476 22100 20528
rect 22152 20516 22158 20528
rect 22250 20519 22308 20525
rect 22250 20516 22262 20519
rect 22152 20488 22262 20516
rect 22152 20476 22158 20488
rect 22250 20485 22262 20488
rect 22296 20485 22308 20519
rect 22250 20479 22308 20485
rect 26694 20476 26700 20528
rect 26752 20516 26758 20528
rect 27402 20519 27460 20525
rect 27402 20516 27414 20519
rect 26752 20488 27414 20516
rect 26752 20476 26758 20488
rect 27402 20485 27414 20488
rect 27448 20485 27460 20519
rect 27402 20479 27460 20485
rect 18506 20451 18512 20460
rect 18432 20423 18512 20451
rect 18049 20411 18107 20417
rect 15838 20340 15844 20392
rect 15896 20380 15902 20392
rect 17218 20380 17224 20392
rect 15896 20352 17224 20380
rect 15896 20340 15902 20352
rect 17218 20340 17224 20352
rect 17276 20340 17282 20392
rect 18064 20380 18092 20411
rect 18506 20408 18512 20423
rect 18564 20448 18570 20460
rect 18564 20420 18657 20448
rect 18564 20408 18570 20420
rect 19334 20408 19340 20460
rect 19392 20448 19398 20460
rect 21269 20451 21327 20457
rect 21269 20448 21281 20451
rect 19392 20420 21281 20448
rect 19392 20408 19398 20420
rect 21269 20417 21281 20420
rect 21315 20417 21327 20451
rect 21450 20448 21456 20460
rect 21411 20420 21456 20448
rect 21269 20411 21327 20417
rect 21450 20408 21456 20420
rect 21508 20408 21514 20460
rect 24302 20448 24308 20460
rect 21560 20420 24164 20448
rect 24263 20420 24308 20448
rect 19426 20380 19432 20392
rect 18064 20352 19432 20380
rect 19426 20340 19432 20352
rect 19484 20340 19490 20392
rect 13541 20315 13599 20321
rect 13541 20312 13553 20315
rect 13464 20284 13553 20312
rect 13541 20281 13553 20284
rect 13587 20281 13599 20315
rect 13541 20275 13599 20281
rect 13630 20272 13636 20324
rect 13688 20312 13694 20324
rect 13688 20284 17540 20312
rect 13688 20272 13694 20284
rect 9398 20244 9404 20256
rect 9359 20216 9404 20244
rect 9398 20204 9404 20216
rect 9456 20204 9462 20256
rect 11054 20244 11060 20256
rect 11015 20216 11060 20244
rect 11054 20204 11060 20216
rect 11112 20204 11118 20256
rect 15194 20244 15200 20256
rect 15155 20216 15200 20244
rect 15194 20204 15200 20216
rect 15252 20204 15258 20256
rect 16574 20204 16580 20256
rect 16632 20244 16638 20256
rect 17405 20247 17463 20253
rect 17405 20244 17417 20247
rect 16632 20216 17417 20244
rect 16632 20204 16638 20216
rect 17405 20213 17417 20216
rect 17451 20213 17463 20247
rect 17512 20244 17540 20284
rect 17586 20272 17592 20324
rect 17644 20312 17650 20324
rect 21560 20312 21588 20420
rect 22002 20380 22008 20392
rect 21963 20352 22008 20380
rect 22002 20340 22008 20352
rect 22060 20340 22066 20392
rect 24136 20380 24164 20420
rect 24302 20408 24308 20420
rect 24360 20408 24366 20460
rect 26234 20408 26240 20460
rect 26292 20448 26298 20460
rect 27154 20448 27160 20460
rect 26292 20420 27160 20448
rect 26292 20408 26298 20420
rect 27154 20408 27160 20420
rect 27212 20408 27218 20460
rect 29472 20457 29500 20556
rect 34882 20516 34888 20528
rect 31726 20488 34888 20516
rect 29457 20451 29515 20457
rect 29457 20448 29469 20451
rect 27264 20420 29469 20448
rect 25314 20380 25320 20392
rect 24136 20352 25320 20380
rect 25314 20340 25320 20352
rect 25372 20340 25378 20392
rect 25498 20340 25504 20392
rect 25556 20380 25562 20392
rect 27264 20380 27292 20420
rect 29457 20417 29469 20420
rect 29503 20417 29515 20451
rect 29457 20411 29515 20417
rect 31726 20380 31754 20488
rect 34882 20476 34888 20488
rect 34940 20476 34946 20528
rect 39316 20516 39344 20556
rect 39942 20544 39948 20596
rect 40000 20584 40006 20596
rect 43898 20584 43904 20596
rect 40000 20556 43904 20584
rect 40000 20544 40006 20556
rect 43898 20544 43904 20556
rect 43956 20544 43962 20596
rect 44082 20584 44088 20596
rect 44043 20556 44088 20584
rect 44082 20544 44088 20556
rect 44140 20544 44146 20596
rect 49142 20544 49148 20596
rect 49200 20584 49206 20596
rect 49513 20587 49571 20593
rect 49513 20584 49525 20587
rect 49200 20556 49525 20584
rect 49200 20544 49206 20556
rect 49513 20553 49525 20556
rect 49559 20553 49571 20587
rect 54478 20584 54484 20596
rect 54439 20556 54484 20584
rect 49513 20547 49571 20553
rect 54478 20544 54484 20556
rect 54536 20544 54542 20596
rect 56321 20587 56379 20593
rect 56321 20553 56333 20587
rect 56367 20584 56379 20587
rect 56594 20584 56600 20596
rect 56367 20556 56600 20584
rect 56367 20553 56379 20556
rect 56321 20547 56379 20553
rect 56594 20544 56600 20556
rect 56652 20584 56658 20596
rect 57882 20584 57888 20596
rect 56652 20556 57888 20584
rect 56652 20544 56658 20556
rect 57882 20544 57888 20556
rect 57940 20544 57946 20596
rect 42518 20516 42524 20528
rect 39316 20488 42524 20516
rect 42518 20476 42524 20488
rect 42576 20476 42582 20528
rect 42972 20519 43030 20525
rect 42972 20485 42984 20519
rect 43018 20516 43030 20519
rect 43070 20516 43076 20528
rect 43018 20488 43076 20516
rect 43018 20485 43030 20488
rect 42972 20479 43030 20485
rect 43070 20476 43076 20488
rect 43128 20476 43134 20528
rect 43530 20476 43536 20528
rect 43588 20516 43594 20528
rect 46017 20519 46075 20525
rect 46017 20516 46029 20519
rect 43588 20488 46029 20516
rect 43588 20476 43594 20488
rect 46017 20485 46029 20488
rect 46063 20485 46075 20519
rect 51442 20516 51448 20528
rect 46017 20479 46075 20485
rect 48148 20488 51448 20516
rect 33505 20451 33563 20457
rect 33505 20417 33517 20451
rect 33551 20448 33563 20451
rect 34606 20448 34612 20460
rect 33551 20420 34612 20448
rect 33551 20417 33563 20420
rect 33505 20411 33563 20417
rect 34606 20408 34612 20420
rect 34664 20408 34670 20460
rect 36078 20408 36084 20460
rect 36136 20448 36142 20460
rect 37645 20451 37703 20457
rect 37645 20448 37657 20451
rect 36136 20420 37657 20448
rect 36136 20408 36142 20420
rect 37645 20417 37657 20420
rect 37691 20417 37703 20451
rect 37645 20411 37703 20417
rect 38381 20451 38439 20457
rect 38381 20417 38393 20451
rect 38427 20448 38439 20451
rect 38746 20448 38752 20460
rect 38427 20420 38752 20448
rect 38427 20417 38439 20420
rect 38381 20411 38439 20417
rect 38746 20408 38752 20420
rect 38804 20408 38810 20460
rect 41414 20408 41420 20460
rect 41472 20448 41478 20460
rect 44358 20448 44364 20460
rect 41472 20420 41517 20448
rect 42536 20420 44364 20448
rect 41472 20408 41478 20420
rect 33321 20383 33379 20389
rect 33321 20380 33333 20383
rect 25556 20352 27292 20380
rect 28184 20352 31754 20380
rect 32416 20352 33333 20380
rect 25556 20340 25562 20352
rect 17644 20284 21588 20312
rect 17644 20272 17650 20284
rect 19794 20244 19800 20256
rect 17512 20216 19800 20244
rect 17405 20207 17463 20213
rect 19794 20204 19800 20216
rect 19852 20204 19858 20256
rect 20070 20204 20076 20256
rect 20128 20244 20134 20256
rect 21269 20247 21327 20253
rect 21269 20244 21281 20247
rect 20128 20216 21281 20244
rect 20128 20204 20134 20216
rect 21269 20213 21281 20216
rect 21315 20213 21327 20247
rect 21269 20207 21327 20213
rect 23198 20204 23204 20256
rect 23256 20244 23262 20256
rect 23385 20247 23443 20253
rect 23385 20244 23397 20247
rect 23256 20216 23397 20244
rect 23256 20204 23262 20216
rect 23385 20213 23397 20216
rect 23431 20213 23443 20247
rect 23385 20207 23443 20213
rect 24210 20204 24216 20256
rect 24268 20244 24274 20256
rect 28184 20244 28212 20352
rect 28258 20272 28264 20324
rect 28316 20312 28322 20324
rect 30653 20315 30711 20321
rect 30653 20312 30665 20315
rect 28316 20284 30665 20312
rect 28316 20272 28322 20284
rect 30653 20281 30665 20284
rect 30699 20281 30711 20315
rect 32416 20312 32444 20352
rect 33321 20349 33333 20352
rect 33367 20349 33379 20383
rect 33321 20343 33379 20349
rect 35161 20383 35219 20389
rect 35161 20349 35173 20383
rect 35207 20349 35219 20383
rect 35161 20343 35219 20349
rect 30653 20275 30711 20281
rect 31726 20284 32444 20312
rect 24268 20216 28212 20244
rect 24268 20204 24274 20216
rect 29730 20204 29736 20256
rect 29788 20244 29794 20256
rect 31726 20244 31754 20284
rect 32490 20272 32496 20324
rect 32548 20312 32554 20324
rect 35176 20312 35204 20343
rect 35342 20340 35348 20392
rect 35400 20380 35406 20392
rect 35437 20383 35495 20389
rect 35437 20380 35449 20383
rect 35400 20352 35449 20380
rect 35400 20340 35406 20352
rect 35437 20349 35449 20352
rect 35483 20349 35495 20383
rect 35437 20343 35495 20349
rect 35802 20340 35808 20392
rect 35860 20380 35866 20392
rect 37274 20380 37280 20392
rect 35860 20352 37280 20380
rect 35860 20340 35866 20352
rect 37274 20340 37280 20352
rect 37332 20380 37338 20392
rect 37461 20383 37519 20389
rect 37461 20380 37473 20383
rect 37332 20352 37473 20380
rect 37332 20340 37338 20352
rect 37461 20349 37473 20352
rect 37507 20349 37519 20383
rect 38654 20380 38660 20392
rect 38615 20352 38660 20380
rect 37461 20343 37519 20349
rect 38654 20340 38660 20352
rect 38712 20340 38718 20392
rect 41138 20340 41144 20392
rect 41196 20380 41202 20392
rect 41233 20383 41291 20389
rect 41233 20380 41245 20383
rect 41196 20352 41245 20380
rect 41196 20340 41202 20352
rect 41233 20349 41245 20352
rect 41279 20349 41291 20383
rect 42536 20380 42564 20420
rect 44358 20408 44364 20420
rect 44416 20408 44422 20460
rect 47026 20448 47032 20460
rect 46987 20420 47032 20448
rect 47026 20408 47032 20420
rect 47084 20408 47090 20460
rect 48148 20392 48176 20488
rect 48406 20457 48412 20460
rect 48400 20411 48412 20457
rect 48464 20448 48470 20460
rect 50264 20457 50292 20488
rect 51442 20476 51448 20488
rect 51500 20516 51506 20528
rect 56502 20516 56508 20528
rect 51500 20488 56508 20516
rect 51500 20476 51506 20488
rect 50522 20457 50528 20460
rect 50249 20451 50307 20457
rect 48464 20420 48500 20448
rect 48406 20408 48412 20411
rect 48464 20408 48470 20420
rect 50249 20417 50261 20451
rect 50295 20417 50307 20451
rect 50249 20411 50307 20417
rect 50516 20411 50528 20457
rect 50580 20448 50586 20460
rect 53116 20457 53144 20488
rect 53101 20451 53159 20457
rect 50580 20420 50616 20448
rect 50522 20408 50528 20411
rect 50580 20408 50586 20420
rect 53101 20417 53113 20451
rect 53147 20417 53159 20451
rect 53101 20411 53159 20417
rect 53368 20451 53426 20457
rect 53368 20417 53380 20451
rect 53414 20448 53426 20451
rect 54110 20448 54116 20460
rect 53414 20420 54116 20448
rect 53414 20417 53426 20420
rect 53368 20411 53426 20417
rect 54110 20408 54116 20420
rect 54168 20408 54174 20460
rect 54956 20457 54984 20488
rect 56502 20476 56508 20488
rect 56560 20476 56566 20528
rect 55214 20457 55220 20460
rect 54941 20451 54999 20457
rect 54941 20417 54953 20451
rect 54987 20417 54999 20451
rect 55208 20448 55220 20457
rect 55175 20420 55220 20448
rect 54941 20411 54999 20417
rect 55208 20411 55220 20420
rect 55214 20408 55220 20411
rect 55272 20408 55278 20460
rect 42702 20380 42708 20392
rect 41233 20343 41291 20349
rect 41340 20352 42564 20380
rect 42663 20352 42708 20380
rect 32548 20284 35204 20312
rect 32548 20272 32554 20284
rect 39666 20272 39672 20324
rect 39724 20312 39730 20324
rect 41340 20312 41368 20352
rect 42702 20340 42708 20352
rect 42760 20340 42766 20392
rect 46842 20380 46848 20392
rect 46803 20352 46848 20380
rect 46842 20340 46848 20352
rect 46900 20340 46906 20392
rect 48130 20380 48136 20392
rect 48091 20352 48136 20380
rect 48130 20340 48136 20352
rect 48188 20340 48194 20392
rect 39724 20284 41368 20312
rect 41432 20284 41736 20312
rect 39724 20272 39730 20284
rect 33686 20244 33692 20256
rect 29788 20216 31754 20244
rect 33647 20216 33692 20244
rect 29788 20204 29794 20216
rect 33686 20204 33692 20216
rect 33744 20204 33750 20256
rect 35894 20204 35900 20256
rect 35952 20244 35958 20256
rect 36541 20247 36599 20253
rect 36541 20244 36553 20247
rect 35952 20216 36553 20244
rect 35952 20204 35958 20216
rect 36541 20213 36553 20216
rect 36587 20213 36599 20247
rect 37826 20244 37832 20256
rect 37787 20216 37832 20244
rect 36541 20207 36599 20213
rect 37826 20204 37832 20216
rect 37884 20204 37890 20256
rect 38194 20204 38200 20256
rect 38252 20244 38258 20256
rect 39758 20244 39764 20256
rect 38252 20216 39764 20244
rect 38252 20204 38258 20216
rect 39758 20204 39764 20216
rect 39816 20204 39822 20256
rect 40218 20204 40224 20256
rect 40276 20244 40282 20256
rect 41432 20244 41460 20284
rect 41598 20244 41604 20256
rect 40276 20216 41460 20244
rect 41559 20216 41604 20244
rect 40276 20204 40282 20216
rect 41598 20204 41604 20216
rect 41656 20204 41662 20256
rect 41708 20244 41736 20284
rect 45278 20272 45284 20324
rect 45336 20312 45342 20324
rect 46293 20315 46351 20321
rect 46293 20312 46305 20315
rect 45336 20284 46305 20312
rect 45336 20272 45342 20284
rect 46293 20281 46305 20284
rect 46339 20312 46351 20315
rect 51626 20312 51632 20324
rect 46339 20284 47532 20312
rect 51587 20284 51632 20312
rect 46339 20281 46351 20284
rect 46293 20275 46351 20281
rect 43438 20244 43444 20256
rect 41708 20216 43444 20244
rect 43438 20204 43444 20216
rect 43496 20244 43502 20256
rect 43806 20244 43812 20256
rect 43496 20216 43812 20244
rect 43496 20204 43502 20216
rect 43806 20204 43812 20216
rect 43864 20204 43870 20256
rect 47210 20244 47216 20256
rect 47171 20216 47216 20244
rect 47210 20204 47216 20216
rect 47268 20204 47274 20256
rect 47504 20244 47532 20284
rect 51626 20272 51632 20284
rect 51684 20272 51690 20324
rect 50982 20244 50988 20256
rect 47504 20216 50988 20244
rect 50982 20204 50988 20216
rect 51040 20204 51046 20256
rect 53098 20204 53104 20256
rect 53156 20244 53162 20256
rect 54386 20244 54392 20256
rect 53156 20216 54392 20244
rect 53156 20204 53162 20216
rect 54386 20204 54392 20216
rect 54444 20244 54450 20256
rect 55858 20244 55864 20256
rect 54444 20216 55864 20244
rect 54444 20204 54450 20216
rect 55858 20204 55864 20216
rect 55916 20204 55922 20256
rect 1104 20154 58880 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 58880 20154
rect 1104 20080 58880 20102
rect 13630 20040 13636 20052
rect 1596 20012 13636 20040
rect 1596 19845 1624 20012
rect 13630 20000 13636 20012
rect 13688 20000 13694 20052
rect 14918 20000 14924 20052
rect 14976 20040 14982 20052
rect 16025 20043 16083 20049
rect 14976 20012 15976 20040
rect 14976 20000 14982 20012
rect 9398 19972 9404 19984
rect 9359 19944 9404 19972
rect 9398 19932 9404 19944
rect 9456 19932 9462 19984
rect 15948 19972 15976 20012
rect 16025 20009 16037 20043
rect 16071 20040 16083 20043
rect 20806 20040 20812 20052
rect 16071 20012 20484 20040
rect 20767 20012 20812 20040
rect 16071 20009 16083 20012
rect 16025 20003 16083 20009
rect 19150 19972 19156 19984
rect 15948 19944 19156 19972
rect 19150 19932 19156 19944
rect 19208 19932 19214 19984
rect 9585 19907 9643 19913
rect 9585 19904 9597 19907
rect 6288 19876 9597 19904
rect 6288 19845 6316 19876
rect 9585 19873 9597 19876
rect 9631 19873 9643 19907
rect 9585 19867 9643 19873
rect 10229 19907 10287 19913
rect 10229 19873 10241 19907
rect 10275 19873 10287 19907
rect 13170 19904 13176 19916
rect 13131 19876 13176 19904
rect 10229 19867 10287 19873
rect 1581 19839 1639 19845
rect 1581 19805 1593 19839
rect 1627 19805 1639 19839
rect 1581 19799 1639 19805
rect 6273 19839 6331 19845
rect 6273 19805 6285 19839
rect 6319 19805 6331 19839
rect 6273 19799 6331 19805
rect 9306 19796 9312 19848
rect 9364 19836 9370 19848
rect 10244 19836 10272 19867
rect 13170 19864 13176 19876
rect 13228 19864 13234 19916
rect 20456 19904 20484 20012
rect 20806 20000 20812 20012
rect 20864 20000 20870 20052
rect 22738 20040 22744 20052
rect 22699 20012 22744 20040
rect 22738 20000 22744 20012
rect 22796 20000 22802 20052
rect 24302 20000 24308 20052
rect 24360 20040 24366 20052
rect 31849 20043 31907 20049
rect 31849 20040 31861 20043
rect 24360 20012 31861 20040
rect 24360 20000 24366 20012
rect 31849 20009 31861 20012
rect 31895 20009 31907 20043
rect 35342 20040 35348 20052
rect 35303 20012 35348 20040
rect 31849 20003 31907 20009
rect 35342 20000 35348 20012
rect 35400 20000 35406 20052
rect 54389 20043 54447 20049
rect 35544 20012 52684 20040
rect 21450 19932 21456 19984
rect 21508 19972 21514 19984
rect 25406 19972 25412 19984
rect 21508 19944 25412 19972
rect 21508 19932 21514 19944
rect 25406 19932 25412 19944
rect 25464 19932 25470 19984
rect 35544 19972 35572 20012
rect 25608 19944 35572 19972
rect 25498 19904 25504 19916
rect 16500 19876 19564 19904
rect 20456 19876 25504 19904
rect 9364 19808 10272 19836
rect 10321 19839 10379 19845
rect 9364 19796 9370 19808
rect 10321 19805 10333 19839
rect 10367 19805 10379 19839
rect 10321 19799 10379 19805
rect 11425 19839 11483 19845
rect 11425 19805 11437 19839
rect 11471 19836 11483 19839
rect 12802 19836 12808 19848
rect 11471 19808 12808 19836
rect 11471 19805 11483 19808
rect 11425 19799 11483 19805
rect 1854 19768 1860 19780
rect 1815 19740 1860 19768
rect 1854 19728 1860 19740
rect 1912 19728 1918 19780
rect 9125 19771 9183 19777
rect 9125 19737 9137 19771
rect 9171 19768 9183 19771
rect 9582 19768 9588 19780
rect 9171 19740 9588 19768
rect 9171 19737 9183 19740
rect 9125 19731 9183 19737
rect 9582 19728 9588 19740
rect 9640 19728 9646 19780
rect 10336 19768 10364 19799
rect 12802 19796 12808 19808
rect 12860 19796 12866 19848
rect 14642 19836 14648 19848
rect 14603 19808 14648 19836
rect 14642 19796 14648 19808
rect 14700 19796 14706 19848
rect 14912 19839 14970 19845
rect 14912 19805 14924 19839
rect 14958 19836 14970 19839
rect 15194 19836 15200 19848
rect 14958 19808 15200 19836
rect 14958 19805 14970 19808
rect 14912 19799 14970 19805
rect 15194 19796 15200 19808
rect 15252 19796 15258 19848
rect 10336 19740 12434 19768
rect 7466 19700 7472 19712
rect 7427 19672 7472 19700
rect 7466 19660 7472 19672
rect 7524 19660 7530 19712
rect 9214 19660 9220 19712
rect 9272 19700 9278 19712
rect 10336 19700 10364 19740
rect 10686 19700 10692 19712
rect 9272 19672 10364 19700
rect 10647 19672 10692 19700
rect 9272 19660 9278 19672
rect 10686 19660 10692 19672
rect 10744 19660 10750 19712
rect 12406 19700 12434 19740
rect 16500 19700 16528 19876
rect 16577 19839 16635 19845
rect 16577 19805 16589 19839
rect 16623 19805 16635 19839
rect 16577 19799 16635 19805
rect 12406 19672 16528 19700
rect 16592 19700 16620 19799
rect 16850 19796 16856 19848
rect 16908 19836 16914 19848
rect 19429 19839 19487 19845
rect 19429 19836 19441 19839
rect 16908 19808 19441 19836
rect 16908 19796 16914 19808
rect 19429 19805 19441 19808
rect 19475 19805 19487 19839
rect 19536 19836 19564 19876
rect 25498 19864 25504 19876
rect 25556 19864 25562 19916
rect 25608 19913 25636 19944
rect 35802 19932 35808 19984
rect 35860 19932 35866 19984
rect 37737 19975 37795 19981
rect 37737 19941 37749 19975
rect 37783 19972 37795 19975
rect 39666 19972 39672 19984
rect 37783 19944 39672 19972
rect 37783 19941 37795 19944
rect 37737 19935 37795 19941
rect 39666 19932 39672 19944
rect 39724 19932 39730 19984
rect 42518 19972 42524 19984
rect 42479 19944 42524 19972
rect 42518 19932 42524 19944
rect 42576 19932 42582 19984
rect 44450 19972 44456 19984
rect 44411 19944 44456 19972
rect 44450 19932 44456 19944
rect 44508 19932 44514 19984
rect 48406 19972 48412 19984
rect 48367 19944 48412 19972
rect 48406 19932 48412 19944
rect 48464 19932 48470 19984
rect 52656 19972 52684 20012
rect 54389 20009 54401 20043
rect 54435 20040 54447 20043
rect 54754 20040 54760 20052
rect 54435 20012 54760 20040
rect 54435 20009 54447 20012
rect 54389 20003 54447 20009
rect 54754 20000 54760 20012
rect 54812 20000 54818 20052
rect 56042 20040 56048 20052
rect 56003 20012 56048 20040
rect 56042 20000 56048 20012
rect 56100 20000 56106 20052
rect 52656 19944 55352 19972
rect 25593 19907 25651 19913
rect 25593 19873 25605 19907
rect 25639 19873 25651 19907
rect 27614 19904 27620 19916
rect 27575 19876 27620 19904
rect 25593 19867 25651 19873
rect 27614 19864 27620 19876
rect 27672 19864 27678 19916
rect 34977 19907 35035 19913
rect 34977 19873 34989 19907
rect 35023 19904 35035 19907
rect 35820 19904 35848 19932
rect 38286 19904 38292 19916
rect 35023 19876 35848 19904
rect 38247 19876 38292 19904
rect 35023 19873 35035 19876
rect 34977 19867 35035 19873
rect 38286 19864 38292 19876
rect 38344 19864 38350 19916
rect 47670 19864 47676 19916
rect 47728 19904 47734 19916
rect 51074 19904 51080 19916
rect 47728 19876 48452 19904
rect 47728 19864 47734 19876
rect 20806 19836 20812 19848
rect 19536 19808 20812 19836
rect 19429 19799 19487 19805
rect 20806 19796 20812 19808
rect 20864 19796 20870 19848
rect 21545 19839 21603 19845
rect 21545 19805 21557 19839
rect 21591 19836 21603 19839
rect 22278 19836 22284 19848
rect 21591 19808 22284 19836
rect 21591 19805 21603 19808
rect 21545 19799 21603 19805
rect 22278 19796 22284 19808
rect 22336 19836 22342 19848
rect 23198 19836 23204 19848
rect 22336 19808 23204 19836
rect 22336 19796 22342 19808
rect 23198 19796 23204 19808
rect 23256 19796 23262 19848
rect 24857 19839 24915 19845
rect 24857 19836 24869 19839
rect 23768 19808 24869 19836
rect 18877 19771 18935 19777
rect 18877 19737 18889 19771
rect 18923 19768 18935 19771
rect 19674 19771 19732 19777
rect 19674 19768 19686 19771
rect 18923 19740 19686 19768
rect 18923 19737 18935 19740
rect 18877 19731 18935 19737
rect 19674 19737 19686 19740
rect 19720 19737 19732 19771
rect 19674 19731 19732 19737
rect 22186 19728 22192 19780
rect 22244 19768 22250 19780
rect 23106 19768 23112 19780
rect 22244 19740 23112 19768
rect 22244 19728 22250 19740
rect 23106 19728 23112 19740
rect 23164 19728 23170 19780
rect 23768 19712 23796 19808
rect 24857 19805 24869 19808
rect 24903 19805 24915 19839
rect 24857 19799 24915 19805
rect 19334 19700 19340 19712
rect 16592 19672 19340 19700
rect 19334 19660 19340 19672
rect 19392 19660 19398 19712
rect 20162 19660 20168 19712
rect 20220 19700 20226 19712
rect 23750 19700 23756 19712
rect 20220 19672 23756 19700
rect 20220 19660 20226 19672
rect 23750 19660 23756 19672
rect 23808 19660 23814 19712
rect 24872 19700 24900 19799
rect 24946 19796 24952 19848
rect 25004 19836 25010 19848
rect 25133 19839 25191 19845
rect 25004 19808 25049 19836
rect 25004 19796 25010 19808
rect 25133 19805 25145 19839
rect 25179 19805 25191 19839
rect 25133 19799 25191 19805
rect 25148 19768 25176 19799
rect 25314 19796 25320 19848
rect 25372 19836 25378 19848
rect 26329 19839 26387 19845
rect 26329 19836 26341 19839
rect 25372 19808 26341 19836
rect 25372 19796 25378 19808
rect 26329 19805 26341 19808
rect 26375 19805 26387 19839
rect 29730 19836 29736 19848
rect 29691 19808 29736 19836
rect 26329 19799 26387 19805
rect 25866 19768 25872 19780
rect 25148 19740 25872 19768
rect 25866 19728 25872 19740
rect 25924 19728 25930 19780
rect 26344 19768 26372 19799
rect 29730 19796 29736 19808
rect 29788 19796 29794 19848
rect 29917 19839 29975 19845
rect 29917 19805 29929 19839
rect 29963 19836 29975 19839
rect 30466 19836 30472 19848
rect 29963 19808 30472 19836
rect 29963 19805 29975 19808
rect 29917 19799 29975 19805
rect 30466 19796 30472 19808
rect 30524 19796 30530 19848
rect 30650 19836 30656 19848
rect 30611 19808 30656 19836
rect 30650 19796 30656 19808
rect 30708 19836 30714 19848
rect 35161 19839 35219 19845
rect 30708 19808 31754 19836
rect 30708 19796 30714 19808
rect 31726 19768 31754 19808
rect 35161 19805 35173 19839
rect 35207 19836 35219 19839
rect 35618 19836 35624 19848
rect 35207 19808 35624 19836
rect 35207 19805 35219 19808
rect 35161 19799 35219 19805
rect 35618 19796 35624 19808
rect 35676 19796 35682 19848
rect 35805 19839 35863 19845
rect 35805 19805 35817 19839
rect 35851 19836 35863 19839
rect 38746 19836 38752 19848
rect 35851 19808 38752 19836
rect 35851 19805 35863 19808
rect 35805 19799 35863 19805
rect 38746 19796 38752 19808
rect 38804 19836 38810 19848
rect 41141 19839 41199 19845
rect 41141 19836 41153 19839
rect 38804 19808 41153 19836
rect 38804 19796 38810 19808
rect 41141 19805 41153 19808
rect 41187 19836 41199 19839
rect 42702 19836 42708 19848
rect 41187 19808 42708 19836
rect 41187 19805 41199 19808
rect 41141 19799 41199 19805
rect 42702 19796 42708 19808
rect 42760 19836 42766 19848
rect 43073 19839 43131 19845
rect 43073 19836 43085 19839
rect 42760 19808 43085 19836
rect 42760 19796 42766 19808
rect 43073 19805 43085 19808
rect 43119 19836 43131 19839
rect 45370 19836 45376 19848
rect 43119 19808 45376 19836
rect 43119 19805 43131 19808
rect 43073 19799 43131 19805
rect 45370 19796 45376 19808
rect 45428 19836 45434 19848
rect 46109 19839 46167 19845
rect 46109 19836 46121 19839
rect 45428 19808 46121 19836
rect 45428 19796 45434 19808
rect 46109 19805 46121 19808
rect 46155 19805 46167 19839
rect 46109 19799 46167 19805
rect 46376 19839 46434 19845
rect 46376 19805 46388 19839
rect 46422 19836 46434 19839
rect 47210 19836 47216 19848
rect 46422 19808 47216 19836
rect 46422 19805 46434 19808
rect 46376 19799 46434 19805
rect 47210 19796 47216 19808
rect 47268 19796 47274 19848
rect 48041 19839 48099 19845
rect 48041 19805 48053 19839
rect 48087 19805 48099 19839
rect 48222 19836 48228 19848
rect 48183 19808 48228 19836
rect 48041 19799 48099 19805
rect 35894 19768 35900 19780
rect 26344 19740 30696 19768
rect 31726 19740 35900 19768
rect 24946 19700 24952 19712
rect 24872 19672 24952 19700
rect 24946 19660 24952 19672
rect 25004 19660 25010 19712
rect 30101 19703 30159 19709
rect 30101 19669 30113 19703
rect 30147 19700 30159 19703
rect 30558 19700 30564 19712
rect 30147 19672 30564 19700
rect 30147 19669 30159 19672
rect 30101 19663 30159 19669
rect 30558 19660 30564 19672
rect 30616 19660 30622 19712
rect 30668 19700 30696 19740
rect 35894 19728 35900 19740
rect 35952 19728 35958 19780
rect 36072 19771 36130 19777
rect 36072 19737 36084 19771
rect 36118 19768 36130 19771
rect 37826 19768 37832 19780
rect 36118 19740 37832 19768
rect 36118 19737 36130 19740
rect 36072 19731 36130 19737
rect 37826 19728 37832 19740
rect 37884 19728 37890 19780
rect 38286 19728 38292 19780
rect 38344 19768 38350 19780
rect 40218 19768 40224 19780
rect 38344 19740 40224 19768
rect 38344 19728 38350 19740
rect 40218 19728 40224 19740
rect 40276 19768 40282 19780
rect 40313 19771 40371 19777
rect 40313 19768 40325 19771
rect 40276 19740 40325 19768
rect 40276 19728 40282 19740
rect 40313 19737 40325 19740
rect 40359 19737 40371 19771
rect 40313 19731 40371 19737
rect 40497 19771 40555 19777
rect 40497 19737 40509 19771
rect 40543 19737 40555 19771
rect 40497 19731 40555 19737
rect 41408 19771 41466 19777
rect 41408 19737 41420 19771
rect 41454 19768 41466 19771
rect 41598 19768 41604 19780
rect 41454 19740 41604 19768
rect 41454 19737 41466 19740
rect 41408 19731 41466 19737
rect 36354 19700 36360 19712
rect 30668 19672 36360 19700
rect 36354 19660 36360 19672
rect 36412 19700 36418 19712
rect 37185 19703 37243 19709
rect 37185 19700 37197 19703
rect 36412 19672 37197 19700
rect 36412 19660 36418 19672
rect 37185 19669 37197 19672
rect 37231 19700 37243 19703
rect 38105 19703 38163 19709
rect 38105 19700 38117 19703
rect 37231 19672 38117 19700
rect 37231 19669 37243 19672
rect 37185 19663 37243 19669
rect 38105 19669 38117 19672
rect 38151 19669 38163 19703
rect 38105 19663 38163 19669
rect 38197 19703 38255 19709
rect 38197 19669 38209 19703
rect 38243 19700 38255 19703
rect 38654 19700 38660 19712
rect 38243 19672 38660 19700
rect 38243 19669 38255 19672
rect 38197 19663 38255 19669
rect 38654 19660 38660 19672
rect 38712 19660 38718 19712
rect 39758 19660 39764 19712
rect 39816 19700 39822 19712
rect 40512 19700 40540 19731
rect 41598 19728 41604 19740
rect 41656 19728 41662 19780
rect 42150 19728 42156 19780
rect 42208 19768 42214 19780
rect 43318 19771 43376 19777
rect 43318 19768 43330 19771
rect 42208 19740 43330 19768
rect 42208 19728 42214 19740
rect 43318 19737 43330 19740
rect 43364 19737 43376 19771
rect 45278 19768 45284 19780
rect 45239 19740 45284 19768
rect 43318 19731 43376 19737
rect 45278 19728 45284 19740
rect 45336 19728 45342 19780
rect 45554 19728 45560 19780
rect 45612 19768 45618 19780
rect 45649 19771 45707 19777
rect 45649 19768 45661 19771
rect 45612 19740 45661 19768
rect 45612 19728 45618 19740
rect 45649 19737 45661 19740
rect 45695 19768 45707 19771
rect 46842 19768 46848 19780
rect 45695 19740 46848 19768
rect 45695 19737 45707 19740
rect 45649 19731 45707 19737
rect 46842 19728 46848 19740
rect 46900 19768 46906 19780
rect 48056 19768 48084 19799
rect 48222 19796 48228 19808
rect 48280 19796 48286 19848
rect 48314 19768 48320 19780
rect 46900 19740 48320 19768
rect 46900 19728 46906 19740
rect 48314 19728 48320 19740
rect 48372 19728 48378 19780
rect 48424 19768 48452 19876
rect 50540 19876 51080 19904
rect 49694 19796 49700 19848
rect 49752 19836 49758 19848
rect 50341 19839 50399 19845
rect 50341 19836 50353 19839
rect 49752 19808 50353 19836
rect 49752 19796 49758 19808
rect 50341 19805 50353 19808
rect 50387 19805 50399 19839
rect 50341 19799 50399 19805
rect 50540 19777 50568 19876
rect 51074 19864 51080 19876
rect 51132 19864 51138 19916
rect 51442 19904 51448 19916
rect 51403 19876 51448 19904
rect 51442 19864 51448 19876
rect 51500 19864 51506 19916
rect 54570 19904 54576 19916
rect 54036 19876 54576 19904
rect 50706 19836 50712 19848
rect 50667 19808 50712 19836
rect 50706 19796 50712 19808
rect 50764 19796 50770 19848
rect 51092 19836 51120 19864
rect 53834 19836 53840 19848
rect 51092 19808 52408 19836
rect 53795 19808 53840 19836
rect 50525 19771 50583 19777
rect 50525 19768 50537 19771
rect 48424 19740 50537 19768
rect 50525 19737 50537 19740
rect 50571 19737 50583 19771
rect 50525 19731 50583 19737
rect 50617 19771 50675 19777
rect 50617 19737 50629 19771
rect 50663 19737 50675 19771
rect 50617 19731 50675 19737
rect 51712 19771 51770 19777
rect 51712 19737 51724 19771
rect 51758 19768 51770 19771
rect 52270 19768 52276 19780
rect 51758 19740 52276 19768
rect 51758 19737 51770 19740
rect 51712 19731 51770 19737
rect 39816 19672 40540 19700
rect 40681 19703 40739 19709
rect 39816 19660 39822 19672
rect 40681 19669 40693 19703
rect 40727 19700 40739 19703
rect 42794 19700 42800 19712
rect 40727 19672 42800 19700
rect 40727 19669 40739 19672
rect 40681 19663 40739 19669
rect 42794 19660 42800 19672
rect 42852 19660 42858 19712
rect 43070 19660 43076 19712
rect 43128 19700 43134 19712
rect 43714 19700 43720 19712
rect 43128 19672 43720 19700
rect 43128 19660 43134 19672
rect 43714 19660 43720 19672
rect 43772 19660 43778 19712
rect 46290 19660 46296 19712
rect 46348 19700 46354 19712
rect 47489 19703 47547 19709
rect 47489 19700 47501 19703
rect 46348 19672 47501 19700
rect 46348 19660 46354 19672
rect 47489 19669 47501 19672
rect 47535 19700 47547 19703
rect 49510 19700 49516 19712
rect 47535 19672 49516 19700
rect 47535 19669 47547 19672
rect 47489 19663 47547 19669
rect 49510 19660 49516 19672
rect 49568 19660 49574 19712
rect 49970 19660 49976 19712
rect 50028 19700 50034 19712
rect 50632 19700 50660 19731
rect 52270 19728 52276 19740
rect 52328 19728 52334 19780
rect 52380 19768 52408 19808
rect 53834 19796 53840 19808
rect 53892 19796 53898 19848
rect 54036 19777 54064 19876
rect 54570 19864 54576 19876
rect 54628 19864 54634 19916
rect 54205 19839 54263 19845
rect 54205 19805 54217 19839
rect 54251 19836 54263 19839
rect 54294 19836 54300 19848
rect 54251 19808 54300 19836
rect 54251 19805 54263 19808
rect 54205 19799 54263 19805
rect 54294 19796 54300 19808
rect 54352 19796 54358 19848
rect 55324 19836 55352 19944
rect 56502 19864 56508 19916
rect 56560 19904 56566 19916
rect 56597 19907 56655 19913
rect 56597 19904 56609 19907
rect 56560 19876 56609 19904
rect 56560 19864 56566 19876
rect 56597 19873 56609 19876
rect 56643 19873 56655 19907
rect 56597 19867 56655 19873
rect 55493 19839 55551 19845
rect 55493 19836 55505 19839
rect 55324 19808 55505 19836
rect 55493 19805 55505 19808
rect 55539 19805 55551 19839
rect 55674 19836 55680 19848
rect 55635 19808 55680 19836
rect 55493 19799 55551 19805
rect 55674 19796 55680 19808
rect 55732 19796 55738 19848
rect 55858 19836 55864 19848
rect 55819 19808 55864 19836
rect 55858 19796 55864 19808
rect 55916 19796 55922 19848
rect 56686 19796 56692 19848
rect 56744 19836 56750 19848
rect 56853 19839 56911 19845
rect 56853 19836 56865 19839
rect 56744 19808 56865 19836
rect 56744 19796 56750 19808
rect 56853 19805 56865 19808
rect 56899 19805 56911 19839
rect 56853 19799 56911 19805
rect 54021 19771 54079 19777
rect 54021 19768 54033 19771
rect 52380 19740 54033 19768
rect 54021 19737 54033 19740
rect 54067 19737 54079 19771
rect 54021 19731 54079 19737
rect 54113 19771 54171 19777
rect 54113 19737 54125 19771
rect 54159 19768 54171 19771
rect 55769 19771 55827 19777
rect 54159 19740 55628 19768
rect 54159 19737 54171 19740
rect 54113 19731 54171 19737
rect 50028 19672 50660 19700
rect 50028 19660 50034 19672
rect 50706 19660 50712 19712
rect 50764 19700 50770 19712
rect 50893 19703 50951 19709
rect 50893 19700 50905 19703
rect 50764 19672 50905 19700
rect 50764 19660 50770 19672
rect 50893 19669 50905 19672
rect 50939 19669 50951 19703
rect 50893 19663 50951 19669
rect 51258 19660 51264 19712
rect 51316 19700 51322 19712
rect 52825 19703 52883 19709
rect 52825 19700 52837 19703
rect 51316 19672 52837 19700
rect 51316 19660 51322 19672
rect 52825 19669 52837 19672
rect 52871 19700 52883 19703
rect 54662 19700 54668 19712
rect 52871 19672 54668 19700
rect 52871 19669 52883 19672
rect 52825 19663 52883 19669
rect 54662 19660 54668 19672
rect 54720 19660 54726 19712
rect 55600 19700 55628 19740
rect 55769 19737 55781 19771
rect 55815 19768 55827 19771
rect 56134 19768 56140 19780
rect 55815 19740 56140 19768
rect 55815 19737 55827 19740
rect 55769 19731 55827 19737
rect 56134 19728 56140 19740
rect 56192 19768 56198 19780
rect 56192 19740 58020 19768
rect 56192 19728 56198 19740
rect 56594 19700 56600 19712
rect 55600 19672 56600 19700
rect 56594 19660 56600 19672
rect 56652 19660 56658 19712
rect 57992 19709 58020 19740
rect 57977 19703 58035 19709
rect 57977 19669 57989 19703
rect 58023 19669 58035 19703
rect 57977 19663 58035 19669
rect 1104 19610 58880 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 58880 19610
rect 1104 19536 58880 19558
rect 8205 19499 8263 19505
rect 8205 19465 8217 19499
rect 8251 19496 8263 19499
rect 13449 19499 13507 19505
rect 8251 19468 13400 19496
rect 8251 19465 8263 19468
rect 8205 19459 8263 19465
rect 7092 19431 7150 19437
rect 7092 19397 7104 19431
rect 7138 19428 7150 19431
rect 7466 19428 7472 19440
rect 7138 19400 7472 19428
rect 7138 19397 7150 19400
rect 7092 19391 7150 19397
rect 7466 19388 7472 19400
rect 7524 19388 7530 19440
rect 13372 19428 13400 19468
rect 13449 19465 13461 19499
rect 13495 19496 13507 19499
rect 30650 19496 30656 19508
rect 13495 19468 30656 19496
rect 13495 19465 13507 19468
rect 13449 19459 13507 19465
rect 30650 19456 30656 19468
rect 30708 19456 30714 19508
rect 33778 19456 33784 19508
rect 33836 19496 33842 19508
rect 33873 19499 33931 19505
rect 33873 19496 33885 19499
rect 33836 19468 33885 19496
rect 33836 19456 33842 19468
rect 33873 19465 33885 19468
rect 33919 19465 33931 19499
rect 34606 19496 34612 19508
rect 34567 19468 34612 19496
rect 33873 19459 33931 19465
rect 18509 19431 18567 19437
rect 13372 19400 16988 19428
rect 1581 19363 1639 19369
rect 1581 19329 1593 19363
rect 1627 19329 1639 19363
rect 1854 19360 1860 19372
rect 1815 19332 1860 19360
rect 1581 19323 1639 19329
rect 1596 19292 1624 19323
rect 1854 19320 1860 19332
rect 1912 19320 1918 19372
rect 6822 19360 6828 19372
rect 6783 19332 6828 19360
rect 6822 19320 6828 19332
rect 6880 19320 6886 19372
rect 8849 19363 8907 19369
rect 8849 19329 8861 19363
rect 8895 19360 8907 19363
rect 10686 19360 10692 19372
rect 8895 19332 10692 19360
rect 8895 19329 8907 19332
rect 8849 19323 8907 19329
rect 10686 19320 10692 19332
rect 10744 19320 10750 19372
rect 11882 19360 11888 19372
rect 11843 19332 11888 19360
rect 11882 19320 11888 19332
rect 11940 19360 11946 19372
rect 14001 19363 14059 19369
rect 11940 19332 13952 19360
rect 11940 19320 11946 19332
rect 12158 19292 12164 19304
rect 1596 19264 2452 19292
rect 12119 19264 12164 19292
rect 2424 19168 2452 19264
rect 12158 19252 12164 19264
rect 12216 19252 12222 19304
rect 13924 19292 13952 19332
rect 14001 19329 14013 19363
rect 14047 19360 14059 19363
rect 15286 19360 15292 19372
rect 14047 19332 15292 19360
rect 14047 19329 14059 19332
rect 14001 19323 14059 19329
rect 15286 19320 15292 19332
rect 15344 19320 15350 19372
rect 16850 19360 16856 19372
rect 16811 19332 16856 19360
rect 16850 19320 16856 19332
rect 16908 19320 16914 19372
rect 16960 19360 16988 19400
rect 18509 19397 18521 19431
rect 18555 19428 18567 19431
rect 22640 19431 22698 19437
rect 18555 19400 22600 19428
rect 18555 19397 18567 19400
rect 18509 19391 18567 19397
rect 17770 19360 17776 19372
rect 16960 19332 17776 19360
rect 17770 19320 17776 19332
rect 17828 19320 17834 19372
rect 19150 19360 19156 19372
rect 19111 19332 19156 19360
rect 19150 19320 19156 19332
rect 19208 19360 19214 19372
rect 20162 19360 20168 19372
rect 19208 19332 20168 19360
rect 19208 19320 19214 19332
rect 20162 19320 20168 19332
rect 20220 19320 20226 19372
rect 22002 19320 22008 19372
rect 22060 19360 22066 19372
rect 22373 19363 22431 19369
rect 22373 19360 22385 19363
rect 22060 19332 22385 19360
rect 22060 19320 22066 19332
rect 22373 19329 22385 19332
rect 22419 19329 22431 19363
rect 22572 19360 22600 19400
rect 22640 19397 22652 19431
rect 22686 19428 22698 19431
rect 24854 19428 24860 19440
rect 22686 19400 24860 19428
rect 22686 19397 22698 19400
rect 22640 19391 22698 19397
rect 24854 19388 24860 19400
rect 24912 19388 24918 19440
rect 25590 19388 25596 19440
rect 25648 19428 25654 19440
rect 30006 19428 30012 19440
rect 25648 19400 30012 19428
rect 25648 19388 25654 19400
rect 30006 19388 30012 19400
rect 30064 19388 30070 19440
rect 32760 19431 32818 19437
rect 30300 19400 31754 19428
rect 30300 19372 30328 19400
rect 24210 19360 24216 19372
rect 22572 19332 24216 19360
rect 22373 19323 22431 19329
rect 24210 19320 24216 19332
rect 24268 19320 24274 19372
rect 24302 19320 24308 19372
rect 24360 19360 24366 19372
rect 24360 19332 24405 19360
rect 24360 19320 24366 19332
rect 26970 19320 26976 19372
rect 27028 19360 27034 19372
rect 27157 19363 27215 19369
rect 27157 19360 27169 19363
rect 27028 19332 27169 19360
rect 27028 19320 27034 19332
rect 27157 19329 27169 19332
rect 27203 19329 27215 19363
rect 30282 19360 30288 19372
rect 30195 19332 30288 19360
rect 27157 19323 27215 19329
rect 14642 19292 14648 19304
rect 13924 19264 14648 19292
rect 14642 19252 14648 19264
rect 14700 19292 14706 19304
rect 16868 19292 16896 19320
rect 14700 19264 16896 19292
rect 17129 19295 17187 19301
rect 14700 19252 14706 19264
rect 17129 19261 17141 19295
rect 17175 19292 17187 19295
rect 17954 19292 17960 19304
rect 17175 19264 17960 19292
rect 17175 19261 17187 19264
rect 17129 19255 17187 19261
rect 17954 19252 17960 19264
rect 18012 19252 18018 19304
rect 20714 19292 20720 19304
rect 20675 19264 20720 19292
rect 20714 19252 20720 19264
rect 20772 19252 20778 19304
rect 25406 19292 25412 19304
rect 25367 19264 25412 19292
rect 25406 19252 25412 19264
rect 25464 19252 25470 19304
rect 21450 19224 21456 19236
rect 17788 19196 21456 19224
rect 2406 19156 2412 19168
rect 2367 19128 2412 19156
rect 2406 19116 2412 19128
rect 2464 19116 2470 19168
rect 10042 19156 10048 19168
rect 10003 19128 10048 19156
rect 10042 19116 10048 19128
rect 10100 19116 10106 19168
rect 15194 19156 15200 19168
rect 15155 19128 15200 19156
rect 15194 19116 15200 19128
rect 15252 19116 15258 19168
rect 16022 19116 16028 19168
rect 16080 19156 16086 19168
rect 17788 19156 17816 19196
rect 21450 19184 21456 19196
rect 21508 19184 21514 19236
rect 23474 19224 23480 19236
rect 23308 19196 23480 19224
rect 16080 19128 17816 19156
rect 16080 19116 16086 19128
rect 17862 19116 17868 19168
rect 17920 19156 17926 19168
rect 23308 19156 23336 19196
rect 23474 19184 23480 19196
rect 23532 19184 23538 19236
rect 23750 19224 23756 19236
rect 23711 19196 23756 19224
rect 23750 19184 23756 19196
rect 23808 19184 23814 19236
rect 27172 19224 27200 19323
rect 30282 19320 30288 19332
rect 30340 19320 30346 19372
rect 30374 19320 30380 19372
rect 30432 19360 30438 19372
rect 30541 19363 30599 19369
rect 30541 19360 30553 19363
rect 30432 19332 30553 19360
rect 30432 19320 30438 19332
rect 30541 19329 30553 19332
rect 30587 19329 30599 19363
rect 31726 19360 31754 19400
rect 32760 19397 32772 19431
rect 32806 19428 32818 19431
rect 33686 19428 33692 19440
rect 32806 19400 33692 19428
rect 32806 19397 32818 19400
rect 32760 19391 32818 19397
rect 33686 19388 33692 19400
rect 33744 19388 33750 19440
rect 33888 19428 33916 19459
rect 34606 19456 34612 19468
rect 34664 19456 34670 19508
rect 35066 19496 35072 19508
rect 35027 19468 35072 19496
rect 35066 19456 35072 19468
rect 35124 19456 35130 19508
rect 35989 19499 36047 19505
rect 35989 19465 36001 19499
rect 36035 19496 36047 19499
rect 36078 19496 36084 19508
rect 36035 19468 36084 19496
rect 36035 19465 36047 19468
rect 35989 19459 36047 19465
rect 36078 19456 36084 19468
rect 36136 19456 36142 19508
rect 36354 19496 36360 19508
rect 36315 19468 36360 19496
rect 36354 19456 36360 19468
rect 36412 19456 36418 19508
rect 36446 19456 36452 19508
rect 36504 19496 36510 19508
rect 59170 19496 59176 19508
rect 36504 19468 37274 19496
rect 36504 19456 36510 19468
rect 34977 19431 35035 19437
rect 34977 19428 34989 19431
rect 33888 19400 34989 19428
rect 34977 19397 34989 19400
rect 35023 19397 35035 19431
rect 37246 19428 37274 19468
rect 41432 19468 59176 19496
rect 41432 19428 41460 19468
rect 59170 19456 59176 19468
rect 59228 19456 59234 19508
rect 42889 19431 42947 19437
rect 42889 19428 42901 19431
rect 37246 19400 41460 19428
rect 41616 19400 42901 19428
rect 34977 19391 35035 19397
rect 32490 19360 32496 19372
rect 31726 19332 32496 19360
rect 30541 19323 30599 19329
rect 32490 19320 32496 19332
rect 32548 19320 32554 19372
rect 33134 19320 33140 19372
rect 33192 19360 33198 19372
rect 39942 19360 39948 19372
rect 33192 19332 39948 19360
rect 33192 19320 33198 19332
rect 39942 19320 39948 19332
rect 40000 19320 40006 19372
rect 40770 19320 40776 19372
rect 40828 19360 40834 19372
rect 41616 19360 41644 19400
rect 42889 19397 42901 19400
rect 42935 19397 42947 19431
rect 42889 19391 42947 19397
rect 43714 19388 43720 19440
rect 43772 19428 43778 19440
rect 43809 19431 43867 19437
rect 43809 19428 43821 19431
rect 43772 19400 43821 19428
rect 43772 19388 43778 19400
rect 43809 19397 43821 19400
rect 43855 19397 43867 19431
rect 43809 19391 43867 19397
rect 43898 19388 43904 19440
rect 43956 19428 43962 19440
rect 51166 19428 51172 19440
rect 43956 19400 50936 19428
rect 51127 19400 51172 19428
rect 43956 19388 43962 19400
rect 40828 19332 41644 19360
rect 41877 19363 41935 19369
rect 40828 19320 40834 19332
rect 41877 19329 41889 19363
rect 41923 19360 41935 19363
rect 42613 19363 42671 19369
rect 42613 19360 42625 19363
rect 41923 19332 42625 19360
rect 41923 19329 41935 19332
rect 41877 19323 41935 19329
rect 42613 19329 42625 19332
rect 42659 19329 42671 19363
rect 42794 19360 42800 19372
rect 42755 19332 42800 19360
rect 42613 19323 42671 19329
rect 42794 19320 42800 19332
rect 42852 19320 42858 19372
rect 43162 19369 43168 19372
rect 42981 19363 43039 19369
rect 42981 19329 42993 19363
rect 43027 19329 43039 19363
rect 42981 19323 43039 19329
rect 43119 19363 43168 19369
rect 43119 19329 43131 19363
rect 43165 19329 43168 19363
rect 43119 19323 43168 19329
rect 34333 19295 34391 19301
rect 34333 19261 34345 19295
rect 34379 19292 34391 19295
rect 34698 19292 34704 19304
rect 34379 19264 34704 19292
rect 34379 19261 34391 19264
rect 34333 19255 34391 19261
rect 34698 19252 34704 19264
rect 34756 19292 34762 19304
rect 35066 19292 35072 19304
rect 34756 19264 35072 19292
rect 34756 19252 34762 19264
rect 35066 19252 35072 19264
rect 35124 19252 35130 19304
rect 35253 19295 35311 19301
rect 35253 19261 35265 19295
rect 35299 19292 35311 19295
rect 36630 19292 36636 19304
rect 35299 19264 36636 19292
rect 35299 19261 35311 19264
rect 35253 19255 35311 19261
rect 36630 19252 36636 19264
rect 36688 19252 36694 19304
rect 37274 19252 37280 19304
rect 37332 19292 37338 19304
rect 41693 19295 41751 19301
rect 41693 19292 41705 19295
rect 37332 19264 41705 19292
rect 37332 19252 37338 19264
rect 41693 19261 41705 19264
rect 41739 19261 41751 19295
rect 41693 19255 41751 19261
rect 31662 19224 31668 19236
rect 27172 19196 28764 19224
rect 17920 19128 23336 19156
rect 17920 19116 17926 19128
rect 23382 19116 23388 19168
rect 23440 19156 23446 19168
rect 26050 19156 26056 19168
rect 23440 19128 26056 19156
rect 23440 19116 23446 19128
rect 26050 19116 26056 19128
rect 26108 19116 26114 19168
rect 28350 19156 28356 19168
rect 28311 19128 28356 19156
rect 28350 19116 28356 19128
rect 28408 19116 28414 19168
rect 28736 19156 28764 19196
rect 31220 19196 31668 19224
rect 31018 19156 31024 19168
rect 28736 19128 31024 19156
rect 31018 19116 31024 19128
rect 31076 19156 31082 19168
rect 31220 19156 31248 19196
rect 31662 19184 31668 19196
rect 31720 19184 31726 19236
rect 33686 19184 33692 19236
rect 33744 19224 33750 19236
rect 42242 19224 42248 19236
rect 33744 19196 42248 19224
rect 33744 19184 33750 19196
rect 42242 19184 42248 19196
rect 42300 19184 42306 19236
rect 35710 19156 35716 19168
rect 31076 19128 31248 19156
rect 35671 19128 35716 19156
rect 31076 19116 31082 19128
rect 35710 19116 35716 19128
rect 35768 19116 35774 19168
rect 36446 19116 36452 19168
rect 36504 19156 36510 19168
rect 41874 19156 41880 19168
rect 36504 19128 41880 19156
rect 36504 19116 36510 19128
rect 41874 19116 41880 19128
rect 41932 19116 41938 19168
rect 42061 19159 42119 19165
rect 42061 19125 42073 19159
rect 42107 19156 42119 19159
rect 42150 19156 42156 19168
rect 42107 19128 42156 19156
rect 42107 19125 42119 19128
rect 42061 19119 42119 19125
rect 42150 19116 42156 19128
rect 42208 19116 42214 19168
rect 42996 19156 43024 19323
rect 43162 19320 43168 19323
rect 43220 19320 43226 19372
rect 45370 19360 45376 19372
rect 45331 19332 45376 19360
rect 45370 19320 45376 19332
rect 45428 19320 45434 19372
rect 45646 19369 45652 19372
rect 45640 19323 45652 19369
rect 45704 19360 45710 19372
rect 45704 19332 45740 19360
rect 45646 19320 45652 19323
rect 45704 19320 45710 19332
rect 47578 19320 47584 19372
rect 47636 19360 47642 19372
rect 47765 19363 47823 19369
rect 47765 19360 47777 19363
rect 47636 19332 47777 19360
rect 47636 19320 47642 19332
rect 47765 19329 47777 19332
rect 47811 19329 47823 19363
rect 47765 19323 47823 19329
rect 47854 19320 47860 19372
rect 47912 19360 47918 19372
rect 48041 19363 48099 19369
rect 48041 19360 48053 19363
rect 47912 19332 48053 19360
rect 47912 19320 47918 19332
rect 48041 19329 48053 19332
rect 48087 19360 48099 19363
rect 48222 19360 48228 19372
rect 48087 19332 48228 19360
rect 48087 19329 48099 19332
rect 48041 19323 48099 19329
rect 48222 19320 48228 19332
rect 48280 19360 48286 19372
rect 50154 19360 50160 19372
rect 48280 19332 50160 19360
rect 48280 19320 48286 19332
rect 50154 19320 50160 19332
rect 50212 19320 50218 19372
rect 50249 19363 50307 19369
rect 50249 19329 50261 19363
rect 50295 19360 50307 19363
rect 50706 19360 50712 19372
rect 50295 19332 50712 19360
rect 50295 19329 50307 19332
rect 50249 19323 50307 19329
rect 50706 19320 50712 19332
rect 50764 19320 50770 19372
rect 50908 19369 50936 19400
rect 51166 19388 51172 19400
rect 51224 19388 51230 19440
rect 52454 19428 52460 19440
rect 51276 19400 52460 19428
rect 50893 19363 50951 19369
rect 50893 19329 50905 19363
rect 50939 19329 50951 19363
rect 51074 19360 51080 19372
rect 51035 19332 51080 19360
rect 50893 19323 50951 19329
rect 51074 19320 51080 19332
rect 51132 19320 51138 19372
rect 51276 19369 51304 19400
rect 52454 19388 52460 19400
rect 52512 19428 52518 19440
rect 54294 19428 54300 19440
rect 52512 19400 54300 19428
rect 52512 19388 52518 19400
rect 54294 19388 54300 19400
rect 54352 19388 54358 19440
rect 51261 19363 51319 19369
rect 51261 19329 51273 19363
rect 51307 19329 51319 19363
rect 52089 19363 52147 19369
rect 52089 19360 52101 19363
rect 51261 19323 51319 19329
rect 51460 19332 52101 19360
rect 43257 19295 43315 19301
rect 43257 19261 43269 19295
rect 43303 19292 43315 19295
rect 44450 19292 44456 19304
rect 43303 19264 44456 19292
rect 43303 19261 43315 19264
rect 43257 19255 43315 19261
rect 44450 19252 44456 19264
rect 44508 19252 44514 19304
rect 48314 19252 48320 19304
rect 48372 19292 48378 19304
rect 50065 19295 50123 19301
rect 50065 19292 50077 19295
rect 48372 19264 50077 19292
rect 48372 19252 48378 19264
rect 50065 19261 50077 19264
rect 50111 19292 50123 19295
rect 51350 19292 51356 19304
rect 50111 19264 51356 19292
rect 50111 19261 50123 19264
rect 50065 19255 50123 19261
rect 51350 19252 51356 19264
rect 51408 19252 51414 19304
rect 46382 19184 46388 19236
rect 46440 19224 46446 19236
rect 51460 19233 51488 19332
rect 52089 19329 52101 19332
rect 52135 19329 52147 19363
rect 52270 19360 52276 19372
rect 52231 19332 52276 19360
rect 52089 19323 52147 19329
rect 52270 19320 52276 19332
rect 52328 19320 52334 19372
rect 51534 19252 51540 19304
rect 51592 19292 51598 19304
rect 51905 19295 51963 19301
rect 51905 19292 51917 19295
rect 51592 19264 51917 19292
rect 51592 19252 51598 19264
rect 51905 19261 51917 19264
rect 51951 19261 51963 19295
rect 51905 19255 51963 19261
rect 51445 19227 51503 19233
rect 46440 19196 51074 19224
rect 46440 19184 46446 19196
rect 43254 19156 43260 19168
rect 42996 19128 43260 19156
rect 43254 19116 43260 19128
rect 43312 19116 43318 19168
rect 43898 19156 43904 19168
rect 43859 19128 43904 19156
rect 43898 19116 43904 19128
rect 43956 19116 43962 19168
rect 46658 19116 46664 19168
rect 46716 19156 46722 19168
rect 46753 19159 46811 19165
rect 46753 19156 46765 19159
rect 46716 19128 46765 19156
rect 46716 19116 46722 19128
rect 46753 19125 46765 19128
rect 46799 19125 46811 19159
rect 46753 19119 46811 19125
rect 46934 19116 46940 19168
rect 46992 19156 46998 19168
rect 47670 19156 47676 19168
rect 46992 19128 47676 19156
rect 46992 19116 46998 19128
rect 47670 19116 47676 19128
rect 47728 19116 47734 19168
rect 50433 19159 50491 19165
rect 50433 19125 50445 19159
rect 50479 19156 50491 19159
rect 50614 19156 50620 19168
rect 50479 19128 50620 19156
rect 50479 19125 50491 19128
rect 50433 19119 50491 19125
rect 50614 19116 50620 19128
rect 50672 19116 50678 19168
rect 51046 19156 51074 19196
rect 51445 19193 51457 19227
rect 51491 19193 51503 19227
rect 51445 19187 51503 19193
rect 58066 19156 58072 19168
rect 51046 19128 58072 19156
rect 58066 19116 58072 19128
rect 58124 19116 58130 19168
rect 1104 19066 58880 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 58880 19066
rect 1104 18992 58880 19014
rect 12158 18912 12164 18964
rect 12216 18952 12222 18964
rect 12621 18955 12679 18961
rect 12621 18952 12633 18955
rect 12216 18924 12633 18952
rect 12216 18912 12222 18924
rect 12621 18921 12633 18924
rect 12667 18921 12679 18955
rect 22094 18952 22100 18964
rect 12621 18915 12679 18921
rect 14476 18924 22100 18952
rect 10505 18887 10563 18893
rect 10505 18853 10517 18887
rect 10551 18884 10563 18887
rect 14476 18884 14504 18924
rect 22094 18912 22100 18924
rect 22152 18912 22158 18964
rect 22649 18955 22707 18961
rect 22649 18952 22661 18955
rect 22204 18924 22661 18952
rect 10551 18856 14504 18884
rect 15841 18887 15899 18893
rect 10551 18853 10563 18856
rect 10505 18847 10563 18853
rect 15841 18853 15853 18887
rect 15887 18884 15899 18887
rect 17586 18884 17592 18896
rect 15887 18856 17592 18884
rect 15887 18853 15899 18856
rect 15841 18847 15899 18853
rect 17586 18844 17592 18856
rect 17644 18844 17650 18896
rect 19426 18884 19432 18896
rect 17880 18856 19432 18884
rect 16390 18776 16396 18828
rect 16448 18816 16454 18828
rect 17880 18816 17908 18856
rect 19426 18844 19432 18856
rect 19484 18844 19490 18896
rect 20806 18844 20812 18896
rect 20864 18884 20870 18896
rect 22204 18884 22232 18924
rect 22649 18921 22661 18924
rect 22695 18921 22707 18955
rect 28350 18952 28356 18964
rect 22649 18915 22707 18921
rect 23400 18924 28356 18952
rect 20864 18856 22232 18884
rect 20864 18844 20870 18856
rect 18046 18816 18052 18828
rect 16448 18788 17908 18816
rect 18007 18788 18052 18816
rect 16448 18776 16454 18788
rect 18046 18776 18052 18788
rect 18104 18776 18110 18828
rect 1581 18751 1639 18757
rect 1581 18717 1593 18751
rect 1627 18748 1639 18751
rect 6273 18751 6331 18757
rect 1627 18720 2452 18748
rect 1627 18717 1639 18720
rect 1581 18711 1639 18717
rect 2424 18692 2452 18720
rect 6273 18717 6285 18751
rect 6319 18717 6331 18751
rect 6273 18711 6331 18717
rect 1854 18680 1860 18692
rect 1815 18652 1860 18680
rect 1854 18640 1860 18652
rect 1912 18640 1918 18692
rect 2406 18680 2412 18692
rect 2367 18652 2412 18680
rect 2406 18640 2412 18652
rect 2464 18640 2470 18692
rect 6288 18680 6316 18711
rect 6822 18708 6828 18760
rect 6880 18748 6886 18760
rect 8202 18748 8208 18760
rect 6880 18720 8208 18748
rect 6880 18708 6886 18720
rect 8202 18708 8208 18720
rect 8260 18748 8266 18760
rect 9125 18751 9183 18757
rect 9125 18748 9137 18751
rect 8260 18720 9137 18748
rect 8260 18708 8266 18720
rect 9125 18717 9137 18720
rect 9171 18717 9183 18751
rect 9125 18711 9183 18717
rect 11425 18751 11483 18757
rect 11425 18717 11437 18751
rect 11471 18748 11483 18751
rect 13722 18748 13728 18760
rect 11471 18720 13728 18748
rect 11471 18717 11483 18720
rect 11425 18711 11483 18717
rect 13722 18708 13728 18720
rect 13780 18708 13786 18760
rect 14461 18751 14519 18757
rect 14461 18717 14473 18751
rect 14507 18748 14519 18751
rect 14550 18748 14556 18760
rect 14507 18720 14556 18748
rect 14507 18717 14519 18720
rect 14461 18711 14519 18717
rect 14550 18708 14556 18720
rect 14608 18708 14614 18760
rect 14728 18751 14786 18757
rect 14728 18717 14740 18751
rect 14774 18748 14786 18751
rect 15194 18748 15200 18760
rect 14774 18720 15200 18748
rect 14774 18717 14786 18720
rect 14728 18711 14786 18717
rect 15194 18708 15200 18720
rect 15252 18708 15258 18760
rect 16574 18748 16580 18760
rect 16535 18720 16580 18748
rect 16574 18708 16580 18720
rect 16632 18708 16638 18760
rect 19429 18751 19487 18757
rect 19429 18717 19441 18751
rect 19475 18748 19487 18751
rect 21269 18751 21327 18757
rect 19475 18720 21128 18748
rect 19475 18717 19487 18720
rect 19429 18711 19487 18717
rect 7006 18680 7012 18692
rect 6288 18652 7012 18680
rect 7006 18640 7012 18652
rect 7064 18640 7070 18692
rect 9392 18683 9450 18689
rect 9392 18649 9404 18683
rect 9438 18680 9450 18683
rect 9674 18680 9680 18692
rect 9438 18652 9680 18680
rect 9438 18649 9450 18652
rect 9392 18643 9450 18649
rect 9674 18640 9680 18652
rect 9732 18640 9738 18692
rect 12342 18640 12348 18692
rect 12400 18680 12406 18692
rect 19696 18683 19754 18689
rect 12400 18652 18460 18680
rect 12400 18640 12406 18652
rect 7098 18572 7104 18624
rect 7156 18612 7162 18624
rect 7469 18615 7527 18621
rect 7469 18612 7481 18615
rect 7156 18584 7481 18612
rect 7156 18572 7162 18584
rect 7469 18581 7481 18584
rect 7515 18581 7527 18615
rect 18432 18612 18460 18652
rect 19696 18649 19708 18683
rect 19742 18680 19754 18683
rect 20990 18680 20996 18692
rect 19742 18652 20996 18680
rect 19742 18649 19754 18652
rect 19696 18643 19754 18649
rect 20990 18640 20996 18652
rect 21048 18640 21054 18692
rect 21100 18680 21128 18720
rect 21269 18717 21281 18751
rect 21315 18748 21327 18751
rect 23400 18748 23428 18924
rect 28350 18912 28356 18924
rect 28408 18912 28414 18964
rect 36446 18952 36452 18964
rect 28460 18924 36452 18952
rect 25317 18887 25375 18893
rect 25317 18853 25329 18887
rect 25363 18884 25375 18887
rect 26694 18884 26700 18896
rect 25363 18856 26700 18884
rect 25363 18853 25375 18856
rect 25317 18847 25375 18853
rect 26694 18844 26700 18856
rect 26752 18844 26758 18896
rect 27062 18844 27068 18896
rect 27120 18884 27126 18896
rect 28460 18884 28488 18924
rect 36446 18912 36452 18924
rect 36504 18912 36510 18964
rect 36998 18912 37004 18964
rect 37056 18952 37062 18964
rect 45557 18955 45615 18961
rect 37056 18924 45508 18952
rect 37056 18912 37062 18924
rect 33686 18884 33692 18896
rect 27120 18856 28488 18884
rect 31312 18856 33692 18884
rect 27120 18844 27126 18856
rect 25961 18819 26019 18825
rect 25961 18785 25973 18819
rect 26007 18816 26019 18819
rect 26050 18816 26056 18828
rect 26007 18788 26056 18816
rect 26007 18785 26019 18788
rect 25961 18779 26019 18785
rect 26050 18776 26056 18788
rect 26108 18816 26114 18828
rect 28258 18816 28264 18828
rect 26108 18788 28264 18816
rect 26108 18776 26114 18788
rect 28258 18776 28264 18788
rect 28316 18776 28322 18828
rect 28350 18776 28356 18828
rect 28408 18816 28414 18828
rect 28408 18788 28453 18816
rect 28408 18776 28414 18788
rect 29454 18776 29460 18828
rect 29512 18816 29518 18828
rect 30282 18816 30288 18828
rect 29512 18788 30288 18816
rect 29512 18776 29518 18788
rect 30282 18776 30288 18788
rect 30340 18776 30346 18828
rect 21315 18720 23428 18748
rect 21315 18717 21327 18720
rect 21269 18711 21327 18717
rect 23474 18708 23480 18760
rect 23532 18748 23538 18760
rect 24581 18751 24639 18757
rect 24581 18748 24593 18751
rect 23532 18720 24593 18748
rect 23532 18708 23538 18720
rect 24581 18717 24593 18720
rect 24627 18717 24639 18751
rect 24762 18748 24768 18760
rect 24723 18720 24768 18748
rect 24581 18711 24639 18717
rect 24762 18708 24768 18720
rect 24820 18708 24826 18760
rect 25774 18748 25780 18760
rect 25735 18720 25780 18748
rect 25774 18708 25780 18720
rect 25832 18708 25838 18760
rect 26510 18748 26516 18760
rect 26471 18720 26516 18748
rect 26510 18708 26516 18720
rect 26568 18748 26574 18760
rect 30006 18748 30012 18760
rect 26568 18720 30012 18748
rect 26568 18708 26574 18720
rect 30006 18708 30012 18720
rect 30064 18708 30070 18760
rect 30558 18757 30564 18760
rect 30552 18748 30564 18757
rect 30519 18720 30564 18748
rect 30552 18711 30564 18720
rect 30558 18708 30564 18711
rect 30616 18708 30622 18760
rect 22002 18680 22008 18692
rect 21100 18652 22008 18680
rect 22002 18640 22008 18652
rect 22060 18640 22066 18692
rect 22186 18640 22192 18692
rect 22244 18680 22250 18692
rect 28350 18680 28356 18692
rect 22244 18652 28356 18680
rect 22244 18640 22250 18652
rect 28350 18640 28356 18652
rect 28408 18640 28414 18692
rect 28626 18640 28632 18692
rect 28684 18680 28690 18692
rect 30650 18680 30656 18692
rect 28684 18652 30656 18680
rect 28684 18640 28690 18652
rect 30650 18640 30656 18652
rect 30708 18640 30714 18692
rect 31312 18680 31340 18856
rect 33686 18844 33692 18856
rect 33744 18844 33750 18896
rect 35710 18884 35716 18896
rect 35623 18856 35716 18884
rect 35710 18844 35716 18856
rect 35768 18884 35774 18896
rect 36081 18887 36139 18893
rect 36081 18884 36093 18887
rect 35768 18856 36093 18884
rect 35768 18844 35774 18856
rect 36081 18853 36093 18856
rect 36127 18884 36139 18887
rect 36354 18884 36360 18896
rect 36127 18856 36360 18884
rect 36127 18853 36139 18856
rect 36081 18847 36139 18853
rect 36354 18844 36360 18856
rect 36412 18844 36418 18896
rect 36817 18887 36875 18893
rect 36817 18853 36829 18887
rect 36863 18884 36875 18887
rect 42610 18884 42616 18896
rect 36863 18856 42616 18884
rect 36863 18853 36875 18856
rect 36817 18847 36875 18853
rect 42610 18844 42616 18856
rect 42668 18844 42674 18896
rect 42705 18887 42763 18893
rect 42705 18853 42717 18887
rect 42751 18884 42763 18887
rect 42886 18884 42892 18896
rect 42751 18856 42892 18884
rect 42751 18853 42763 18856
rect 42705 18847 42763 18853
rect 42886 18844 42892 18856
rect 42944 18844 42950 18896
rect 43254 18884 43260 18896
rect 43088 18856 43260 18884
rect 31478 18776 31484 18828
rect 31536 18816 31542 18828
rect 31754 18816 31760 18828
rect 31536 18788 31760 18816
rect 31536 18776 31542 18788
rect 31754 18776 31760 18788
rect 31812 18776 31818 18828
rect 37461 18819 37519 18825
rect 37461 18785 37473 18819
rect 37507 18816 37519 18819
rect 38286 18816 38292 18828
rect 37507 18788 38292 18816
rect 37507 18785 37519 18788
rect 37461 18779 37519 18785
rect 38286 18776 38292 18788
rect 38344 18776 38350 18828
rect 38657 18819 38715 18825
rect 38657 18785 38669 18819
rect 38703 18816 38715 18819
rect 40034 18816 40040 18828
rect 38703 18788 40040 18816
rect 38703 18785 38715 18788
rect 38657 18779 38715 18785
rect 40034 18776 40040 18788
rect 40092 18776 40098 18828
rect 41233 18819 41291 18825
rect 41233 18785 41245 18819
rect 41279 18816 41291 18819
rect 42242 18816 42248 18828
rect 41279 18788 42248 18816
rect 41279 18785 41291 18788
rect 41233 18779 41291 18785
rect 31662 18708 31668 18760
rect 31720 18748 31726 18760
rect 32217 18751 32275 18757
rect 32217 18748 32229 18751
rect 31720 18720 32229 18748
rect 31720 18708 31726 18720
rect 32217 18717 32229 18720
rect 32263 18717 32275 18751
rect 32217 18711 32275 18717
rect 32401 18751 32459 18757
rect 32401 18717 32413 18751
rect 32447 18717 32459 18751
rect 32401 18711 32459 18717
rect 33781 18751 33839 18757
rect 33781 18717 33793 18751
rect 33827 18748 33839 18751
rect 33827 18720 35848 18748
rect 33827 18717 33839 18720
rect 33781 18711 33839 18717
rect 31128 18652 31340 18680
rect 20809 18615 20867 18621
rect 20809 18612 20821 18615
rect 18432 18584 20821 18612
rect 7469 18575 7527 18581
rect 20809 18581 20821 18584
rect 20855 18612 20867 18615
rect 22278 18612 22284 18624
rect 20855 18584 22284 18612
rect 20855 18581 20867 18584
rect 20809 18575 20867 18581
rect 22278 18572 22284 18584
rect 22336 18572 22342 18624
rect 23382 18572 23388 18624
rect 23440 18612 23446 18624
rect 24673 18615 24731 18621
rect 24673 18612 24685 18615
rect 23440 18584 24685 18612
rect 23440 18572 23446 18584
rect 24673 18581 24685 18584
rect 24719 18581 24731 18615
rect 24673 18575 24731 18581
rect 25685 18615 25743 18621
rect 25685 18581 25697 18615
rect 25731 18612 25743 18615
rect 26786 18612 26792 18624
rect 25731 18584 26792 18612
rect 25731 18581 25743 18584
rect 25685 18575 25743 18581
rect 26786 18572 26792 18584
rect 26844 18572 26850 18624
rect 26878 18572 26884 18624
rect 26936 18612 26942 18624
rect 31128 18612 31156 18652
rect 31386 18640 31392 18692
rect 31444 18680 31450 18692
rect 32416 18680 32444 18711
rect 31444 18652 32444 18680
rect 31444 18640 31450 18652
rect 33686 18640 33692 18692
rect 33744 18680 33750 18692
rect 34057 18683 34115 18689
rect 34057 18680 34069 18683
rect 33744 18652 34069 18680
rect 33744 18640 33750 18652
rect 34057 18649 34069 18652
rect 34103 18649 34115 18683
rect 35820 18680 35848 18720
rect 35894 18708 35900 18760
rect 35952 18748 35958 18760
rect 37185 18751 37243 18757
rect 37185 18748 37197 18751
rect 35952 18720 37197 18748
rect 35952 18708 35958 18720
rect 37185 18717 37197 18720
rect 37231 18717 37243 18751
rect 38838 18748 38844 18760
rect 38799 18720 38844 18748
rect 37185 18711 37243 18717
rect 38838 18708 38844 18720
rect 38896 18708 38902 18760
rect 41248 18748 41276 18779
rect 42242 18776 42248 18788
rect 42300 18776 42306 18828
rect 38948 18720 41276 18748
rect 42890 18745 42948 18751
rect 42890 18738 42902 18745
rect 42936 18738 42948 18745
rect 36722 18680 36728 18692
rect 35820 18652 36728 18680
rect 34057 18643 34115 18649
rect 36722 18640 36728 18652
rect 36780 18640 36786 18692
rect 38378 18640 38384 18692
rect 38436 18680 38442 18692
rect 38948 18680 38976 18720
rect 38436 18652 38976 18680
rect 38436 18640 38442 18652
rect 39206 18640 39212 18692
rect 39264 18680 39270 18692
rect 42886 18686 42892 18738
rect 42944 18686 42950 18738
rect 43088 18689 43116 18856
rect 43254 18844 43260 18856
rect 43312 18884 43318 18896
rect 45278 18884 45284 18896
rect 43312 18856 45284 18884
rect 43312 18844 43318 18856
rect 45278 18844 45284 18856
rect 45336 18844 45342 18896
rect 45480 18884 45508 18924
rect 45557 18921 45569 18955
rect 45603 18952 45615 18955
rect 45646 18952 45652 18964
rect 45603 18924 45652 18952
rect 45603 18921 45615 18924
rect 45557 18915 45615 18921
rect 45646 18912 45652 18924
rect 45704 18912 45710 18964
rect 46569 18955 46627 18961
rect 46569 18921 46581 18955
rect 46615 18952 46627 18955
rect 47026 18952 47032 18964
rect 46615 18924 47032 18952
rect 46615 18921 46627 18924
rect 46569 18915 46627 18921
rect 47026 18912 47032 18924
rect 47084 18912 47090 18964
rect 58066 18952 58072 18964
rect 58027 18924 58072 18952
rect 58066 18912 58072 18924
rect 58124 18912 58130 18964
rect 53834 18884 53840 18896
rect 45480 18856 53840 18884
rect 53834 18844 53840 18856
rect 53892 18844 53898 18896
rect 43349 18819 43407 18825
rect 43349 18785 43361 18819
rect 43395 18816 43407 18819
rect 44082 18816 44088 18828
rect 43395 18788 44088 18816
rect 43395 18785 43407 18788
rect 43349 18779 43407 18785
rect 44082 18776 44088 18788
rect 44140 18776 44146 18828
rect 53926 18816 53932 18828
rect 44192 18788 53932 18816
rect 43622 18708 43628 18760
rect 43680 18748 43686 18760
rect 44192 18748 44220 18788
rect 53926 18776 53932 18788
rect 53984 18776 53990 18828
rect 55030 18776 55036 18828
rect 55088 18816 55094 18828
rect 58434 18816 58440 18828
rect 55088 18788 55720 18816
rect 55088 18776 55094 18788
rect 43680 18720 44220 18748
rect 45281 18751 45339 18757
rect 43680 18708 43686 18720
rect 45281 18717 45293 18751
rect 45327 18717 45339 18751
rect 45281 18711 45339 18717
rect 45373 18751 45431 18757
rect 45373 18717 45385 18751
rect 45419 18748 45431 18751
rect 45922 18748 45928 18760
rect 45419 18720 45928 18748
rect 45419 18717 45431 18720
rect 45373 18711 45431 18717
rect 42982 18683 43040 18689
rect 39264 18652 42012 18680
rect 39264 18640 39270 18652
rect 26936 18584 31156 18612
rect 26936 18572 26942 18584
rect 31202 18572 31208 18624
rect 31260 18612 31266 18624
rect 31665 18615 31723 18621
rect 31665 18612 31677 18615
rect 31260 18584 31677 18612
rect 31260 18572 31266 18584
rect 31665 18581 31677 18584
rect 31711 18581 31723 18615
rect 31665 18575 31723 18581
rect 32585 18615 32643 18621
rect 32585 18581 32597 18615
rect 32631 18612 32643 18615
rect 33042 18612 33048 18624
rect 32631 18584 33048 18612
rect 32631 18581 32643 18584
rect 32585 18575 32643 18581
rect 33042 18572 33048 18584
rect 33100 18572 33106 18624
rect 34514 18572 34520 18624
rect 34572 18612 34578 18624
rect 35434 18612 35440 18624
rect 34572 18584 35440 18612
rect 34572 18572 34578 18584
rect 35434 18572 35440 18584
rect 35492 18572 35498 18624
rect 37182 18572 37188 18624
rect 37240 18612 37246 18624
rect 37277 18615 37335 18621
rect 37277 18612 37289 18615
rect 37240 18584 37289 18612
rect 37240 18572 37246 18584
rect 37277 18581 37289 18584
rect 37323 18581 37335 18615
rect 39022 18612 39028 18624
rect 38983 18584 39028 18612
rect 37277 18575 37335 18581
rect 39022 18572 39028 18584
rect 39080 18572 39086 18624
rect 40586 18612 40592 18624
rect 40547 18584 40592 18612
rect 40586 18572 40592 18584
rect 40644 18572 40650 18624
rect 40954 18612 40960 18624
rect 40915 18584 40960 18612
rect 40954 18572 40960 18584
rect 41012 18572 41018 18624
rect 41049 18615 41107 18621
rect 41049 18581 41061 18615
rect 41095 18612 41107 18615
rect 41874 18612 41880 18624
rect 41095 18584 41880 18612
rect 41095 18581 41107 18584
rect 41049 18575 41107 18581
rect 41874 18572 41880 18584
rect 41932 18572 41938 18624
rect 41984 18612 42012 18652
rect 42982 18649 42994 18683
rect 43028 18649 43040 18683
rect 42982 18643 43040 18649
rect 43073 18683 43131 18689
rect 43073 18649 43085 18683
rect 43119 18649 43131 18683
rect 43073 18643 43131 18649
rect 42996 18612 43024 18643
rect 43162 18640 43168 18692
rect 43220 18689 43226 18692
rect 43220 18683 43269 18689
rect 43220 18649 43223 18683
rect 43257 18680 43269 18683
rect 43714 18680 43720 18692
rect 43257 18652 43720 18680
rect 43257 18649 43269 18652
rect 43220 18643 43269 18649
rect 43220 18640 43226 18643
rect 43714 18640 43720 18652
rect 43772 18640 43778 18692
rect 45296 18680 45324 18711
rect 45922 18708 45928 18720
rect 45980 18708 45986 18760
rect 46014 18708 46020 18760
rect 46072 18748 46078 18760
rect 46290 18748 46296 18760
rect 46072 18720 46117 18748
rect 46251 18720 46296 18748
rect 46072 18708 46078 18720
rect 46290 18708 46296 18720
rect 46348 18708 46354 18760
rect 46382 18708 46388 18760
rect 46440 18748 46446 18760
rect 47854 18748 47860 18760
rect 46440 18720 47860 18748
rect 46440 18708 46446 18720
rect 47854 18708 47860 18720
rect 47912 18708 47918 18760
rect 48314 18748 48320 18760
rect 48275 18720 48320 18748
rect 48314 18708 48320 18720
rect 48372 18708 48378 18760
rect 48498 18748 48504 18760
rect 48459 18720 48504 18748
rect 48498 18708 48504 18720
rect 48556 18708 48562 18760
rect 51350 18708 51356 18760
rect 51408 18748 51414 18760
rect 55306 18748 55312 18760
rect 51408 18720 55312 18748
rect 51408 18708 51414 18720
rect 55306 18708 55312 18720
rect 55364 18748 55370 18760
rect 55692 18757 55720 18788
rect 55784 18788 58440 18816
rect 55493 18751 55551 18757
rect 55493 18748 55505 18751
rect 55364 18720 55505 18748
rect 55364 18708 55370 18720
rect 55493 18717 55505 18720
rect 55539 18717 55551 18751
rect 55493 18711 55551 18717
rect 55677 18751 55735 18757
rect 55677 18717 55689 18751
rect 55723 18717 55735 18751
rect 55677 18711 55735 18717
rect 45554 18680 45560 18692
rect 45296 18652 45560 18680
rect 45554 18640 45560 18652
rect 45612 18640 45618 18692
rect 46201 18683 46259 18689
rect 46201 18680 46213 18683
rect 45655 18652 46213 18680
rect 41984 18584 43024 18612
rect 45278 18572 45284 18624
rect 45336 18612 45342 18624
rect 45655 18612 45683 18652
rect 46201 18649 46213 18652
rect 46247 18680 46259 18683
rect 46750 18680 46756 18692
rect 46247 18652 46756 18680
rect 46247 18649 46259 18652
rect 46201 18643 46259 18649
rect 46750 18640 46756 18652
rect 46808 18640 46814 18692
rect 46842 18640 46848 18692
rect 46900 18680 46906 18692
rect 47121 18683 47179 18689
rect 47121 18680 47133 18683
rect 46900 18652 47133 18680
rect 46900 18640 46906 18652
rect 47121 18649 47133 18652
rect 47167 18649 47179 18683
rect 47121 18643 47179 18649
rect 47489 18683 47547 18689
rect 47489 18649 47501 18683
rect 47535 18680 47547 18683
rect 47578 18680 47584 18692
rect 47535 18652 47584 18680
rect 47535 18649 47547 18652
rect 47489 18643 47547 18649
rect 47578 18640 47584 18652
rect 47636 18640 47642 18692
rect 49694 18680 49700 18692
rect 47688 18652 49700 18680
rect 45336 18584 45683 18612
rect 45336 18572 45342 18584
rect 45830 18572 45836 18624
rect 45888 18612 45894 18624
rect 47688 18612 47716 18652
rect 49694 18640 49700 18652
rect 49752 18640 49758 18692
rect 53834 18640 53840 18692
rect 53892 18680 53898 18692
rect 55784 18680 55812 18788
rect 58434 18776 58440 18788
rect 58492 18776 58498 18828
rect 56594 18708 56600 18760
rect 56652 18748 56658 18760
rect 56965 18751 57023 18757
rect 56965 18748 56977 18751
rect 56652 18720 56977 18748
rect 56652 18708 56658 18720
rect 56965 18717 56977 18720
rect 57011 18717 57023 18751
rect 57974 18748 57980 18760
rect 57935 18720 57980 18748
rect 56965 18711 57023 18717
rect 57974 18708 57980 18720
rect 58032 18708 58038 18760
rect 57238 18680 57244 18692
rect 53892 18652 55812 18680
rect 57199 18652 57244 18680
rect 53892 18640 53898 18652
rect 57238 18640 57244 18652
rect 57296 18640 57302 18692
rect 45888 18584 47716 18612
rect 48685 18615 48743 18621
rect 45888 18572 45894 18584
rect 48685 18581 48697 18615
rect 48731 18612 48743 18615
rect 48774 18612 48780 18624
rect 48731 18584 48780 18612
rect 48731 18581 48743 18584
rect 48685 18575 48743 18581
rect 48774 18572 48780 18584
rect 48832 18572 48838 18624
rect 55858 18612 55864 18624
rect 55819 18584 55864 18612
rect 55858 18572 55864 18584
rect 55916 18572 55922 18624
rect 1104 18522 58880 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 58880 18522
rect 1104 18448 58880 18470
rect 6822 18368 6828 18420
rect 6880 18368 6886 18420
rect 7929 18411 7987 18417
rect 7929 18377 7941 18411
rect 7975 18408 7987 18411
rect 20898 18408 20904 18420
rect 7975 18380 20904 18408
rect 7975 18377 7987 18380
rect 7929 18371 7987 18377
rect 20898 18368 20904 18380
rect 20956 18368 20962 18420
rect 20990 18368 20996 18420
rect 21048 18408 21054 18420
rect 22005 18411 22063 18417
rect 22005 18408 22017 18411
rect 21048 18380 22017 18408
rect 21048 18368 21054 18380
rect 22005 18377 22017 18380
rect 22051 18377 22063 18411
rect 22005 18371 22063 18377
rect 22094 18368 22100 18420
rect 22152 18408 22158 18420
rect 22152 18380 22508 18408
rect 22152 18368 22158 18380
rect 6840 18340 6868 18368
rect 12710 18340 12716 18352
rect 6564 18312 6868 18340
rect 11992 18312 12716 18340
rect 6564 18281 6592 18312
rect 6549 18275 6607 18281
rect 6549 18241 6561 18275
rect 6595 18241 6607 18275
rect 6549 18235 6607 18241
rect 6816 18275 6874 18281
rect 6816 18241 6828 18275
rect 6862 18272 6874 18275
rect 7098 18272 7104 18284
rect 6862 18244 7104 18272
rect 6862 18241 6874 18244
rect 6816 18235 6874 18241
rect 7098 18232 7104 18244
rect 7156 18232 7162 18284
rect 8110 18232 8116 18284
rect 8168 18272 8174 18284
rect 11992 18281 12020 18312
rect 12710 18300 12716 18312
rect 12768 18300 12774 18352
rect 16301 18343 16359 18349
rect 16301 18309 16313 18343
rect 16347 18340 16359 18343
rect 17862 18340 17868 18352
rect 16347 18312 17868 18340
rect 16347 18309 16359 18312
rect 16301 18303 16359 18309
rect 17862 18300 17868 18312
rect 17920 18300 17926 18352
rect 22186 18340 22192 18352
rect 19168 18312 22192 18340
rect 8573 18275 8631 18281
rect 8573 18272 8585 18275
rect 8168 18244 8585 18272
rect 8168 18232 8174 18244
rect 8573 18241 8585 18244
rect 8619 18241 8631 18275
rect 8573 18235 8631 18241
rect 11977 18275 12035 18281
rect 11977 18241 11989 18275
rect 12023 18241 12035 18275
rect 11977 18235 12035 18241
rect 12250 18232 12256 18284
rect 12308 18272 12314 18284
rect 12805 18275 12863 18281
rect 12805 18272 12817 18275
rect 12308 18244 12817 18272
rect 12308 18232 12314 18244
rect 12805 18241 12817 18244
rect 12851 18241 12863 18275
rect 16022 18272 16028 18284
rect 15983 18244 16028 18272
rect 12805 18235 12863 18241
rect 16022 18232 16028 18244
rect 16080 18232 16086 18284
rect 16117 18275 16175 18281
rect 16117 18241 16129 18275
rect 16163 18272 16175 18275
rect 16390 18272 16396 18284
rect 16163 18244 16396 18272
rect 16163 18241 16175 18244
rect 16117 18235 16175 18241
rect 16390 18232 16396 18244
rect 16448 18232 16454 18284
rect 16850 18232 16856 18284
rect 16908 18272 16914 18284
rect 19168 18281 19196 18312
rect 22186 18300 22192 18312
rect 22244 18300 22250 18352
rect 22370 18340 22376 18352
rect 22331 18312 22376 18340
rect 22370 18300 22376 18312
rect 22428 18300 22434 18352
rect 22480 18340 22508 18380
rect 23566 18368 23572 18420
rect 23624 18408 23630 18420
rect 24302 18408 24308 18420
rect 23624 18380 24308 18408
rect 23624 18368 23630 18380
rect 24302 18368 24308 18380
rect 24360 18408 24366 18420
rect 28810 18408 28816 18420
rect 24360 18380 28816 18408
rect 24360 18368 24366 18380
rect 28810 18368 28816 18380
rect 28868 18368 28874 18420
rect 30466 18368 30472 18420
rect 30524 18408 30530 18420
rect 30837 18411 30895 18417
rect 30837 18408 30849 18411
rect 30524 18380 30849 18408
rect 30524 18368 30530 18380
rect 30837 18377 30849 18380
rect 30883 18377 30895 18411
rect 30837 18371 30895 18377
rect 31297 18411 31355 18417
rect 31297 18377 31309 18411
rect 31343 18408 31355 18411
rect 40954 18408 40960 18420
rect 31343 18380 40960 18408
rect 31343 18377 31355 18380
rect 31297 18371 31355 18377
rect 40954 18368 40960 18380
rect 41012 18368 41018 18420
rect 42061 18411 42119 18417
rect 42061 18377 42073 18411
rect 42107 18408 42119 18411
rect 42107 18380 42564 18408
rect 42107 18377 42119 18380
rect 42061 18371 42119 18377
rect 26970 18340 26976 18352
rect 22480 18312 26976 18340
rect 26970 18300 26976 18312
rect 27028 18300 27034 18352
rect 27792 18343 27850 18349
rect 27792 18309 27804 18343
rect 27838 18340 27850 18343
rect 28902 18340 28908 18352
rect 27838 18312 28908 18340
rect 27838 18309 27850 18312
rect 27792 18303 27850 18309
rect 28902 18300 28908 18312
rect 28960 18300 28966 18352
rect 41782 18340 41788 18352
rect 31036 18312 38884 18340
rect 17129 18275 17187 18281
rect 17129 18272 17141 18275
rect 16908 18244 17141 18272
rect 16908 18232 16914 18244
rect 17129 18241 17141 18244
rect 17175 18241 17187 18275
rect 17129 18235 17187 18241
rect 17396 18275 17454 18281
rect 17396 18241 17408 18275
rect 17442 18272 17454 18275
rect 19153 18275 19211 18281
rect 17442 18244 18552 18272
rect 17442 18241 17454 18244
rect 17396 18235 17454 18241
rect 11054 18164 11060 18216
rect 11112 18204 11118 18216
rect 11885 18207 11943 18213
rect 11885 18204 11897 18207
rect 11112 18176 11897 18204
rect 11112 18164 11118 18176
rect 11885 18173 11897 18176
rect 11931 18173 11943 18207
rect 18524 18204 18552 18244
rect 19153 18241 19165 18275
rect 19199 18241 19211 18275
rect 19153 18235 19211 18241
rect 19242 18232 19248 18284
rect 19300 18272 19306 18284
rect 21634 18272 21640 18284
rect 19300 18244 21640 18272
rect 19300 18232 19306 18244
rect 21634 18232 21640 18244
rect 21692 18232 21698 18284
rect 22278 18232 22284 18284
rect 22336 18272 22342 18284
rect 22465 18275 22523 18281
rect 22465 18272 22477 18275
rect 22336 18244 22477 18272
rect 22336 18232 22342 18244
rect 22465 18241 22477 18244
rect 22511 18241 22523 18275
rect 23566 18272 23572 18284
rect 23527 18244 23572 18272
rect 22465 18235 22523 18241
rect 23566 18232 23572 18244
rect 23624 18232 23630 18284
rect 23661 18275 23719 18281
rect 23661 18241 23673 18275
rect 23707 18241 23719 18275
rect 23661 18235 23719 18241
rect 24305 18275 24363 18281
rect 24305 18241 24317 18275
rect 24351 18241 24363 18275
rect 24305 18235 24363 18241
rect 19426 18204 19432 18216
rect 18524 18176 19432 18204
rect 11885 18167 11943 18173
rect 19426 18164 19432 18176
rect 19484 18164 19490 18216
rect 22649 18207 22707 18213
rect 22649 18173 22661 18207
rect 22695 18204 22707 18207
rect 23290 18204 23296 18216
rect 22695 18176 23296 18204
rect 22695 18173 22707 18176
rect 22649 18167 22707 18173
rect 23290 18164 23296 18176
rect 23348 18164 23354 18216
rect 23474 18164 23480 18216
rect 23532 18204 23538 18216
rect 23676 18204 23704 18235
rect 23532 18176 23704 18204
rect 24320 18204 24348 18235
rect 24762 18232 24768 18284
rect 24820 18272 24826 18284
rect 27062 18272 27068 18284
rect 24820 18244 27068 18272
rect 24820 18232 24826 18244
rect 27062 18232 27068 18244
rect 27120 18232 27126 18284
rect 27154 18232 27160 18284
rect 27212 18272 27218 18284
rect 27525 18275 27583 18281
rect 27525 18272 27537 18275
rect 27212 18244 27537 18272
rect 27212 18232 27218 18244
rect 27525 18241 27537 18244
rect 27571 18241 27583 18275
rect 27525 18235 27583 18241
rect 28258 18232 28264 18284
rect 28316 18272 28322 18284
rect 29546 18272 29552 18284
rect 28316 18244 29552 18272
rect 28316 18232 28322 18244
rect 29546 18232 29552 18244
rect 29604 18232 29610 18284
rect 29733 18275 29791 18281
rect 29733 18241 29745 18275
rect 29779 18241 29791 18275
rect 29733 18235 29791 18241
rect 29748 18204 29776 18235
rect 29822 18232 29828 18284
rect 29880 18272 29886 18284
rect 30009 18275 30067 18281
rect 29880 18244 29925 18272
rect 29880 18232 29886 18244
rect 30009 18241 30021 18275
rect 30055 18241 30067 18275
rect 30009 18235 30067 18241
rect 30101 18275 30159 18281
rect 30101 18241 30113 18275
rect 30147 18272 30236 18275
rect 31036 18272 31064 18312
rect 31202 18272 31208 18284
rect 30147 18247 31064 18272
rect 30147 18241 30159 18247
rect 30208 18244 31064 18247
rect 31163 18244 31208 18272
rect 30101 18235 30159 18241
rect 29914 18204 29920 18216
rect 24320 18176 27568 18204
rect 29748 18176 29920 18204
rect 23532 18164 23538 18176
rect 12345 18139 12403 18145
rect 12345 18105 12357 18139
rect 12391 18136 12403 18139
rect 12526 18136 12532 18148
rect 12391 18108 12532 18136
rect 12391 18105 12403 18108
rect 12345 18099 12403 18105
rect 12526 18096 12532 18108
rect 12584 18096 12590 18148
rect 18509 18139 18567 18145
rect 18509 18105 18521 18139
rect 18555 18136 18567 18139
rect 18555 18108 20484 18136
rect 18555 18105 18567 18108
rect 18509 18099 18567 18105
rect 9766 18068 9772 18080
rect 9727 18040 9772 18068
rect 9766 18028 9772 18040
rect 9824 18028 9830 18080
rect 13446 18028 13452 18080
rect 13504 18068 13510 18080
rect 14001 18071 14059 18077
rect 14001 18068 14013 18071
rect 13504 18040 14013 18068
rect 13504 18028 13510 18040
rect 14001 18037 14013 18040
rect 14047 18037 14059 18071
rect 14001 18031 14059 18037
rect 16022 18028 16028 18080
rect 16080 18068 16086 18080
rect 16206 18068 16212 18080
rect 16080 18040 16212 18068
rect 16080 18028 16086 18040
rect 16206 18028 16212 18040
rect 16264 18028 16270 18080
rect 16390 18028 16396 18080
rect 16448 18068 16454 18080
rect 20349 18071 20407 18077
rect 20349 18068 20361 18071
rect 16448 18040 20361 18068
rect 16448 18028 16454 18040
rect 20349 18037 20361 18040
rect 20395 18037 20407 18071
rect 20456 18068 20484 18108
rect 23382 18096 23388 18148
rect 23440 18136 23446 18148
rect 25501 18139 25559 18145
rect 25501 18136 25513 18139
rect 23440 18108 25513 18136
rect 23440 18096 23446 18108
rect 25501 18105 25513 18108
rect 25547 18105 25559 18139
rect 25501 18099 25559 18105
rect 26234 18096 26240 18148
rect 26292 18136 26298 18148
rect 27154 18136 27160 18148
rect 26292 18108 27160 18136
rect 26292 18096 26298 18108
rect 27154 18096 27160 18108
rect 27212 18096 27218 18148
rect 23566 18068 23572 18080
rect 20456 18040 23572 18068
rect 20349 18031 20407 18037
rect 23566 18028 23572 18040
rect 23624 18028 23630 18080
rect 23845 18071 23903 18077
rect 23845 18037 23857 18071
rect 23891 18068 23903 18071
rect 26510 18068 26516 18080
rect 23891 18040 26516 18068
rect 23891 18037 23903 18040
rect 23845 18031 23903 18037
rect 26510 18028 26516 18040
rect 26568 18028 26574 18080
rect 27540 18068 27568 18176
rect 29914 18164 29920 18176
rect 29972 18164 29978 18216
rect 30024 18204 30052 18235
rect 31202 18232 31208 18244
rect 31260 18232 31266 18284
rect 32122 18232 32128 18284
rect 32180 18272 32186 18284
rect 33870 18272 33876 18284
rect 32180 18244 33876 18272
rect 32180 18232 32186 18244
rect 33870 18232 33876 18244
rect 33928 18232 33934 18284
rect 34698 18272 34704 18284
rect 34659 18244 34704 18272
rect 34698 18232 34704 18244
rect 34756 18272 34762 18284
rect 35437 18275 35495 18281
rect 35437 18272 35449 18275
rect 34756 18244 35449 18272
rect 34756 18232 34762 18244
rect 35437 18241 35449 18244
rect 35483 18241 35495 18275
rect 38746 18272 38752 18284
rect 38707 18244 38752 18272
rect 35437 18235 35495 18241
rect 38746 18232 38752 18244
rect 38804 18232 38810 18284
rect 30190 18204 30196 18216
rect 30024 18176 30196 18204
rect 30190 18164 30196 18176
rect 30248 18164 30254 18216
rect 31481 18207 31539 18213
rect 31481 18173 31493 18207
rect 31527 18204 31539 18207
rect 31662 18204 31668 18216
rect 31527 18176 31668 18204
rect 31527 18173 31539 18176
rect 31481 18167 31539 18173
rect 31662 18164 31668 18176
rect 31720 18164 31726 18216
rect 35342 18164 35348 18216
rect 35400 18204 35406 18216
rect 35529 18207 35587 18213
rect 35529 18204 35541 18207
rect 35400 18176 35541 18204
rect 35400 18164 35406 18176
rect 35529 18173 35541 18176
rect 35575 18173 35587 18207
rect 35529 18167 35587 18173
rect 35618 18164 35624 18216
rect 35676 18204 35682 18216
rect 35713 18207 35771 18213
rect 35713 18204 35725 18207
rect 35676 18176 35725 18204
rect 35676 18164 35682 18176
rect 35713 18173 35725 18176
rect 35759 18204 35771 18207
rect 38378 18204 38384 18216
rect 35759 18176 38384 18204
rect 35759 18173 35771 18176
rect 35713 18167 35771 18173
rect 38378 18164 38384 18176
rect 38436 18164 38442 18216
rect 38856 18204 38884 18312
rect 41386 18312 41644 18340
rect 41743 18312 41788 18340
rect 39022 18272 39028 18284
rect 38983 18244 39028 18272
rect 39022 18232 39028 18244
rect 39080 18232 39086 18284
rect 41386 18204 41414 18312
rect 41509 18275 41567 18281
rect 41509 18241 41521 18275
rect 41555 18241 41567 18275
rect 41509 18235 41567 18241
rect 38856 18176 41414 18204
rect 33321 18139 33379 18145
rect 33321 18136 33333 18139
rect 28460 18108 33333 18136
rect 28460 18068 28488 18108
rect 33321 18105 33333 18108
rect 33367 18105 33379 18139
rect 33321 18099 33379 18105
rect 33962 18096 33968 18148
rect 34020 18136 34026 18148
rect 35069 18139 35127 18145
rect 35069 18136 35081 18139
rect 34020 18108 35081 18136
rect 34020 18096 34026 18108
rect 35069 18105 35081 18108
rect 35115 18105 35127 18139
rect 35069 18099 35127 18105
rect 27540 18040 28488 18068
rect 28810 18028 28816 18080
rect 28868 18068 28874 18080
rect 28905 18071 28963 18077
rect 28905 18068 28917 18071
rect 28868 18040 28917 18068
rect 28868 18028 28874 18040
rect 28905 18037 28917 18040
rect 28951 18037 28963 18071
rect 28905 18031 28963 18037
rect 29549 18071 29607 18077
rect 29549 18037 29561 18071
rect 29595 18068 29607 18071
rect 29914 18068 29920 18080
rect 29595 18040 29920 18068
rect 29595 18037 29607 18040
rect 29549 18031 29607 18037
rect 29914 18028 29920 18040
rect 29972 18028 29978 18080
rect 30006 18028 30012 18080
rect 30064 18068 30070 18080
rect 33778 18068 33784 18080
rect 30064 18040 33784 18068
rect 30064 18028 30070 18040
rect 33778 18028 33784 18040
rect 33836 18068 33842 18080
rect 34422 18068 34428 18080
rect 33836 18040 34428 18068
rect 33836 18028 33842 18040
rect 34422 18028 34428 18040
rect 34480 18028 34486 18080
rect 36630 18028 36636 18080
rect 36688 18068 36694 18080
rect 39022 18068 39028 18080
rect 36688 18040 39028 18068
rect 36688 18028 36694 18040
rect 39022 18028 39028 18040
rect 39080 18028 39086 18080
rect 40034 18028 40040 18080
rect 40092 18068 40098 18080
rect 40129 18071 40187 18077
rect 40129 18068 40141 18071
rect 40092 18040 40141 18068
rect 40092 18028 40098 18040
rect 40129 18037 40141 18040
rect 40175 18068 40187 18071
rect 40954 18068 40960 18080
rect 40175 18040 40960 18068
rect 40175 18037 40187 18040
rect 40129 18031 40187 18037
rect 40954 18028 40960 18040
rect 41012 18028 41018 18080
rect 41524 18068 41552 18235
rect 41616 18136 41644 18312
rect 41782 18300 41788 18312
rect 41840 18300 41846 18352
rect 42426 18340 42432 18352
rect 41892 18312 42432 18340
rect 41892 18281 41920 18312
rect 42426 18300 42432 18312
rect 42484 18300 42490 18352
rect 41693 18275 41751 18281
rect 41693 18241 41705 18275
rect 41739 18241 41751 18275
rect 41693 18235 41751 18241
rect 41877 18275 41935 18281
rect 41877 18241 41889 18275
rect 41923 18241 41935 18275
rect 42536 18272 42564 18380
rect 42610 18368 42616 18420
rect 42668 18408 42674 18420
rect 45830 18408 45836 18420
rect 42668 18380 45836 18408
rect 42668 18368 42674 18380
rect 45830 18368 45836 18380
rect 45888 18368 45894 18420
rect 45922 18368 45928 18420
rect 45980 18408 45986 18420
rect 46385 18411 46443 18417
rect 46385 18408 46397 18411
rect 45980 18380 46397 18408
rect 45980 18368 45986 18380
rect 46385 18377 46397 18380
rect 46431 18377 46443 18411
rect 46385 18371 46443 18377
rect 46566 18368 46572 18420
rect 46624 18408 46630 18420
rect 53834 18408 53840 18420
rect 46624 18380 53840 18408
rect 46624 18368 46630 18380
rect 53834 18368 53840 18380
rect 53892 18368 53898 18420
rect 53926 18368 53932 18420
rect 53984 18408 53990 18420
rect 54021 18411 54079 18417
rect 54021 18408 54033 18411
rect 53984 18380 54033 18408
rect 53984 18368 53990 18380
rect 54021 18377 54033 18380
rect 54067 18377 54079 18411
rect 54021 18371 54079 18377
rect 54941 18411 54999 18417
rect 54941 18377 54953 18411
rect 54987 18408 54999 18411
rect 55030 18408 55036 18420
rect 54987 18380 55036 18408
rect 54987 18377 54999 18380
rect 54941 18371 54999 18377
rect 42794 18300 42800 18352
rect 42852 18340 42858 18352
rect 42981 18343 43039 18349
rect 42981 18340 42993 18343
rect 42852 18312 42993 18340
rect 42852 18300 42858 18312
rect 42981 18309 42993 18312
rect 43027 18309 43039 18343
rect 42981 18303 43039 18309
rect 45278 18300 45284 18352
rect 45336 18340 45342 18352
rect 46017 18343 46075 18349
rect 46017 18340 46029 18343
rect 45336 18312 46029 18340
rect 45336 18300 45342 18312
rect 46017 18309 46029 18312
rect 46063 18309 46075 18343
rect 46017 18303 46075 18309
rect 46109 18343 46167 18349
rect 46109 18309 46121 18343
rect 46155 18340 46167 18343
rect 46658 18340 46664 18352
rect 46155 18312 46664 18340
rect 46155 18309 46167 18312
rect 46109 18303 46167 18309
rect 46658 18300 46664 18312
rect 46716 18300 46722 18352
rect 46934 18300 46940 18352
rect 46992 18340 46998 18352
rect 50062 18340 50068 18352
rect 46992 18312 50068 18340
rect 46992 18300 46998 18312
rect 50062 18300 50068 18312
rect 50120 18300 50126 18352
rect 51046 18312 53972 18340
rect 42613 18275 42671 18281
rect 42613 18272 42625 18275
rect 42536 18244 42625 18272
rect 41877 18235 41935 18241
rect 42613 18241 42625 18244
rect 42659 18241 42671 18275
rect 42613 18235 42671 18241
rect 41708 18204 41736 18235
rect 42702 18232 42708 18284
rect 42760 18272 42766 18284
rect 42760 18244 42805 18272
rect 42760 18232 42766 18244
rect 42886 18232 42892 18284
rect 42944 18272 42950 18284
rect 42944 18244 42989 18272
rect 42944 18232 42950 18244
rect 43070 18232 43076 18284
rect 43128 18281 43134 18284
rect 43128 18272 43136 18281
rect 43346 18272 43352 18284
rect 43128 18244 43352 18272
rect 43128 18235 43136 18244
rect 43128 18232 43134 18235
rect 43346 18232 43352 18244
rect 43404 18232 43410 18284
rect 44174 18232 44180 18284
rect 44232 18272 44238 18284
rect 45833 18275 45891 18281
rect 45833 18272 45845 18275
rect 44232 18244 45845 18272
rect 44232 18232 44238 18244
rect 45833 18241 45845 18244
rect 45879 18241 45891 18275
rect 45833 18235 45891 18241
rect 46201 18275 46259 18281
rect 46201 18241 46213 18275
rect 46247 18272 46259 18275
rect 46382 18272 46388 18284
rect 46247 18244 46388 18272
rect 46247 18241 46259 18244
rect 46201 18235 46259 18241
rect 46382 18232 46388 18244
rect 46440 18232 46446 18284
rect 48774 18281 48780 18284
rect 48768 18272 48780 18281
rect 48735 18244 48780 18272
rect 48768 18235 48780 18244
rect 48774 18232 48780 18235
rect 48832 18232 48838 18284
rect 49602 18232 49608 18284
rect 49660 18272 49666 18284
rect 51046 18272 51074 18312
rect 49660 18244 51074 18272
rect 49660 18232 49666 18244
rect 42150 18204 42156 18216
rect 41708 18176 42156 18204
rect 42150 18164 42156 18176
rect 42208 18164 42214 18216
rect 42242 18164 42248 18216
rect 42300 18204 42306 18216
rect 43162 18204 43168 18216
rect 42300 18176 43168 18204
rect 42300 18164 42306 18176
rect 43162 18164 43168 18176
rect 43220 18164 43226 18216
rect 48130 18164 48136 18216
rect 48188 18204 48194 18216
rect 48501 18207 48559 18213
rect 48501 18204 48513 18207
rect 48188 18176 48513 18204
rect 48188 18164 48194 18176
rect 48501 18173 48513 18176
rect 48547 18173 48559 18207
rect 48501 18167 48559 18173
rect 43257 18139 43315 18145
rect 43257 18136 43269 18139
rect 41616 18108 43269 18136
rect 43257 18105 43269 18108
rect 43303 18105 43315 18139
rect 43257 18099 43315 18105
rect 49436 18108 50016 18136
rect 49436 18068 49464 18108
rect 41524 18040 49464 18068
rect 49602 18028 49608 18080
rect 49660 18068 49666 18080
rect 49881 18071 49939 18077
rect 49881 18068 49893 18071
rect 49660 18040 49893 18068
rect 49660 18028 49666 18040
rect 49881 18037 49893 18040
rect 49927 18037 49939 18071
rect 49988 18068 50016 18108
rect 52178 18068 52184 18080
rect 49988 18040 52184 18068
rect 49881 18031 49939 18037
rect 52178 18028 52184 18040
rect 52236 18028 52242 18080
rect 53944 18068 53972 18312
rect 54036 18272 54064 18371
rect 55030 18368 55036 18380
rect 55088 18368 55094 18420
rect 57146 18408 57152 18420
rect 55692 18380 57152 18408
rect 54665 18343 54723 18349
rect 54665 18309 54677 18343
rect 54711 18340 54723 18343
rect 55692 18340 55720 18380
rect 57146 18368 57152 18380
rect 57204 18368 57210 18420
rect 56502 18340 56508 18352
rect 54711 18312 55720 18340
rect 55784 18312 56508 18340
rect 54711 18309 54723 18312
rect 54665 18303 54723 18309
rect 54389 18275 54447 18281
rect 54389 18272 54401 18275
rect 54036 18244 54401 18272
rect 54389 18241 54401 18244
rect 54435 18241 54447 18275
rect 54570 18272 54576 18284
rect 54531 18244 54576 18272
rect 54389 18235 54447 18241
rect 54570 18232 54576 18244
rect 54628 18232 54634 18284
rect 55784 18281 55812 18312
rect 56502 18300 56508 18312
rect 56560 18300 56566 18352
rect 54757 18275 54815 18281
rect 54757 18241 54769 18275
rect 54803 18241 54815 18275
rect 54757 18235 54815 18241
rect 55769 18275 55827 18281
rect 55769 18241 55781 18275
rect 55815 18241 55827 18275
rect 55769 18235 55827 18241
rect 54772 18204 54800 18235
rect 55858 18232 55864 18284
rect 55916 18272 55922 18284
rect 56025 18275 56083 18281
rect 56025 18272 56037 18275
rect 55916 18244 56037 18272
rect 55916 18232 55922 18244
rect 56025 18241 56037 18244
rect 56071 18241 56083 18275
rect 56025 18235 56083 18241
rect 54404 18176 54800 18204
rect 54404 18148 54432 18176
rect 54386 18096 54392 18148
rect 54444 18096 54450 18148
rect 57606 18068 57612 18080
rect 53944 18040 57612 18068
rect 57606 18028 57612 18040
rect 57664 18028 57670 18080
rect 1104 17978 58880 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 58880 17978
rect 1104 17904 58880 17926
rect 8018 17864 8024 17876
rect 7979 17836 8024 17864
rect 8018 17824 8024 17836
rect 8076 17824 8082 17876
rect 9122 17864 9128 17876
rect 8220 17836 9128 17864
rect 7561 17799 7619 17805
rect 7561 17765 7573 17799
rect 7607 17796 7619 17799
rect 8110 17796 8116 17808
rect 7607 17768 8116 17796
rect 7607 17765 7619 17768
rect 7561 17759 7619 17765
rect 8110 17756 8116 17768
rect 8168 17756 8174 17808
rect 8220 17737 8248 17836
rect 9122 17824 9128 17836
rect 9180 17864 9186 17876
rect 9180 17836 9536 17864
rect 9180 17824 9186 17836
rect 9508 17808 9536 17836
rect 9674 17824 9680 17876
rect 9732 17864 9738 17876
rect 11333 17867 11391 17873
rect 11333 17864 11345 17867
rect 9732 17836 11345 17864
rect 9732 17824 9738 17836
rect 11333 17833 11345 17836
rect 11379 17833 11391 17867
rect 13354 17864 13360 17876
rect 13315 17836 13360 17864
rect 11333 17827 11391 17833
rect 13354 17824 13360 17836
rect 13412 17824 13418 17876
rect 14826 17824 14832 17876
rect 14884 17864 14890 17876
rect 15473 17867 15531 17873
rect 15473 17864 15485 17867
rect 14884 17836 15485 17864
rect 14884 17824 14890 17836
rect 15473 17833 15485 17836
rect 15519 17864 15531 17867
rect 15562 17864 15568 17876
rect 15519 17836 15568 17864
rect 15519 17833 15531 17836
rect 15473 17827 15531 17833
rect 15562 17824 15568 17836
rect 15620 17824 15626 17876
rect 15657 17867 15715 17873
rect 15657 17833 15669 17867
rect 15703 17864 15715 17867
rect 16666 17864 16672 17876
rect 15703 17836 16672 17864
rect 15703 17833 15715 17836
rect 15657 17827 15715 17833
rect 16666 17824 16672 17836
rect 16724 17824 16730 17876
rect 17310 17864 17316 17876
rect 17271 17836 17316 17864
rect 17310 17824 17316 17836
rect 17368 17824 17374 17876
rect 19334 17824 19340 17876
rect 19392 17864 19398 17876
rect 19429 17867 19487 17873
rect 19429 17864 19441 17867
rect 19392 17836 19441 17864
rect 19392 17824 19398 17836
rect 19429 17833 19441 17836
rect 19475 17833 19487 17867
rect 19429 17827 19487 17833
rect 19702 17824 19708 17876
rect 19760 17864 19766 17876
rect 23382 17864 23388 17876
rect 19760 17836 23388 17864
rect 19760 17824 19766 17836
rect 23382 17824 23388 17836
rect 23440 17824 23446 17876
rect 24578 17864 24584 17876
rect 24539 17836 24584 17864
rect 24578 17824 24584 17836
rect 24636 17824 24642 17876
rect 28626 17864 28632 17876
rect 26160 17836 27292 17864
rect 28587 17836 28632 17864
rect 9490 17756 9496 17808
rect 9548 17796 9554 17808
rect 12986 17796 12992 17808
rect 9548 17768 12992 17796
rect 9548 17756 9554 17768
rect 12986 17756 12992 17768
rect 13044 17756 13050 17808
rect 13170 17796 13176 17808
rect 13131 17768 13176 17796
rect 13170 17756 13176 17768
rect 13228 17756 13234 17808
rect 21269 17799 21327 17805
rect 21269 17796 21281 17799
rect 13280 17768 21281 17796
rect 7285 17731 7343 17737
rect 7285 17697 7297 17731
rect 7331 17728 7343 17731
rect 8205 17731 8263 17737
rect 8205 17728 8217 17731
rect 7331 17700 8217 17728
rect 7331 17697 7343 17700
rect 7285 17691 7343 17697
rect 8205 17697 8217 17700
rect 8251 17697 8263 17731
rect 8205 17691 8263 17697
rect 8481 17731 8539 17737
rect 8481 17697 8493 17731
rect 8527 17728 8539 17731
rect 9125 17731 9183 17737
rect 9125 17728 9137 17731
rect 8527 17700 9137 17728
rect 8527 17697 8539 17700
rect 8481 17691 8539 17697
rect 9125 17697 9137 17700
rect 9171 17728 9183 17731
rect 13280 17728 13308 17768
rect 21269 17765 21281 17768
rect 21315 17765 21327 17799
rect 26160 17796 26188 17836
rect 21269 17759 21327 17765
rect 23308 17768 26188 17796
rect 22646 17728 22652 17740
rect 9171 17700 13308 17728
rect 14660 17700 22652 17728
rect 9171 17697 9183 17700
rect 9125 17691 9183 17697
rect 1578 17660 1584 17672
rect 1539 17632 1584 17660
rect 1578 17620 1584 17632
rect 1636 17620 1642 17672
rect 7193 17663 7251 17669
rect 7193 17629 7205 17663
rect 7239 17629 7251 17663
rect 7193 17623 7251 17629
rect 8297 17663 8355 17669
rect 8297 17629 8309 17663
rect 8343 17629 8355 17663
rect 8297 17623 8355 17629
rect 8389 17663 8447 17669
rect 8389 17629 8401 17663
rect 8435 17660 8447 17663
rect 9214 17660 9220 17672
rect 8435 17657 8524 17660
rect 8588 17657 9220 17660
rect 8435 17632 9220 17657
rect 8435 17629 8447 17632
rect 8496 17629 8616 17632
rect 8389 17623 8447 17629
rect 1854 17592 1860 17604
rect 1815 17564 1860 17592
rect 1854 17552 1860 17564
rect 1912 17552 1918 17604
rect 7208 17592 7236 17623
rect 8312 17592 8340 17623
rect 9214 17620 9220 17632
rect 9272 17660 9278 17672
rect 9309 17663 9367 17669
rect 9309 17660 9321 17663
rect 9272 17632 9321 17660
rect 9272 17620 9278 17632
rect 9309 17629 9321 17632
rect 9355 17629 9367 17663
rect 9490 17660 9496 17672
rect 9451 17632 9496 17660
rect 9309 17623 9367 17629
rect 9490 17620 9496 17632
rect 9548 17620 9554 17672
rect 10042 17620 10048 17672
rect 10100 17660 10106 17672
rect 10137 17663 10195 17669
rect 10137 17660 10149 17663
rect 10100 17632 10149 17660
rect 10100 17620 10106 17632
rect 10137 17629 10149 17632
rect 10183 17629 10195 17663
rect 10137 17623 10195 17629
rect 12897 17663 12955 17669
rect 12897 17629 12909 17663
rect 12943 17660 12955 17663
rect 13078 17660 13084 17672
rect 12943 17632 13084 17660
rect 12943 17629 12955 17632
rect 12897 17623 12955 17629
rect 13078 17620 13084 17632
rect 13136 17620 13142 17672
rect 14660 17669 14688 17700
rect 22646 17688 22652 17700
rect 22704 17688 22710 17740
rect 23198 17728 23204 17740
rect 23159 17700 23204 17728
rect 23198 17688 23204 17700
rect 23256 17688 23262 17740
rect 14645 17663 14703 17669
rect 14645 17629 14657 17663
rect 14691 17629 14703 17663
rect 14826 17660 14832 17672
rect 14787 17632 14832 17660
rect 14645 17623 14703 17629
rect 14826 17620 14832 17632
rect 14884 17620 14890 17672
rect 16142 17663 16200 17669
rect 14936 17632 16068 17660
rect 9398 17592 9404 17604
rect 7208 17564 9404 17592
rect 9398 17552 9404 17564
rect 9456 17592 9462 17604
rect 14936 17592 14964 17632
rect 9456 17564 12434 17592
rect 9456 17552 9462 17564
rect 9582 17484 9588 17536
rect 9640 17524 9646 17536
rect 9677 17527 9735 17533
rect 9677 17524 9689 17527
rect 9640 17496 9689 17524
rect 9640 17484 9646 17496
rect 9677 17493 9689 17496
rect 9723 17493 9735 17527
rect 12406 17524 12434 17564
rect 14660 17564 14964 17592
rect 15289 17595 15347 17601
rect 14660 17524 14688 17564
rect 15289 17561 15301 17595
rect 15335 17592 15347 17595
rect 15930 17592 15936 17604
rect 15335 17564 15936 17592
rect 15335 17561 15347 17564
rect 15289 17555 15347 17561
rect 15930 17552 15936 17564
rect 15988 17552 15994 17604
rect 12406 17496 14688 17524
rect 14737 17527 14795 17533
rect 9677 17487 9735 17493
rect 14737 17493 14749 17527
rect 14783 17524 14795 17527
rect 15378 17524 15384 17536
rect 14783 17496 15384 17524
rect 14783 17493 14795 17496
rect 14737 17487 14795 17493
rect 15378 17484 15384 17496
rect 15436 17484 15442 17536
rect 15499 17527 15557 17533
rect 15499 17493 15511 17527
rect 15545 17524 15557 17527
rect 15838 17524 15844 17536
rect 15545 17496 15844 17524
rect 15545 17493 15557 17496
rect 15499 17487 15557 17493
rect 15838 17484 15844 17496
rect 15896 17484 15902 17536
rect 16040 17524 16068 17632
rect 16142 17629 16154 17663
rect 16188 17660 16200 17663
rect 19429 17663 19487 17669
rect 16188 17632 16344 17660
rect 16188 17629 16200 17632
rect 16142 17623 16200 17629
rect 16316 17604 16344 17632
rect 19429 17629 19441 17663
rect 19475 17660 19487 17663
rect 19518 17660 19524 17672
rect 19475 17632 19524 17660
rect 19475 17629 19487 17632
rect 19429 17623 19487 17629
rect 19518 17620 19524 17632
rect 19576 17620 19582 17672
rect 19613 17663 19671 17669
rect 19613 17629 19625 17663
rect 19659 17660 19671 17663
rect 19978 17660 19984 17672
rect 19659 17632 19984 17660
rect 19659 17629 19671 17632
rect 19613 17623 19671 17629
rect 19978 17620 19984 17632
rect 20036 17620 20042 17672
rect 20073 17663 20131 17669
rect 20073 17629 20085 17663
rect 20119 17660 20131 17663
rect 23308 17660 23336 17768
rect 24578 17688 24584 17740
rect 24636 17728 24642 17740
rect 25038 17728 25044 17740
rect 24636 17700 25044 17728
rect 24636 17688 24642 17700
rect 25038 17688 25044 17700
rect 25096 17728 25102 17740
rect 25133 17731 25191 17737
rect 25133 17728 25145 17731
rect 25096 17700 25145 17728
rect 25096 17688 25102 17700
rect 25133 17697 25145 17700
rect 25179 17728 25191 17731
rect 26050 17728 26056 17740
rect 25179 17700 26056 17728
rect 25179 17697 25191 17700
rect 25133 17691 25191 17697
rect 26050 17688 26056 17700
rect 26108 17688 26114 17740
rect 27264 17728 27292 17836
rect 28626 17824 28632 17836
rect 28684 17824 28690 17876
rect 30650 17864 30656 17876
rect 28966 17836 30656 17864
rect 27338 17756 27344 17808
rect 27396 17796 27402 17808
rect 28966 17796 28994 17836
rect 30650 17824 30656 17836
rect 30708 17824 30714 17876
rect 32125 17867 32183 17873
rect 32125 17833 32137 17867
rect 32171 17864 32183 17867
rect 38749 17867 38807 17873
rect 32171 17836 36768 17864
rect 32171 17833 32183 17836
rect 32125 17827 32183 17833
rect 27396 17768 28994 17796
rect 30285 17799 30343 17805
rect 27396 17756 27402 17768
rect 30285 17765 30297 17799
rect 30331 17796 30343 17799
rect 30374 17796 30380 17808
rect 30331 17768 30380 17796
rect 30331 17765 30343 17768
rect 30285 17759 30343 17765
rect 30374 17756 30380 17768
rect 30432 17756 30438 17808
rect 36740 17796 36768 17836
rect 38749 17833 38761 17867
rect 38795 17864 38807 17867
rect 38838 17864 38844 17876
rect 38795 17836 38844 17864
rect 38795 17833 38807 17836
rect 38749 17827 38807 17833
rect 38838 17824 38844 17836
rect 38896 17824 38902 17876
rect 46014 17864 46020 17876
rect 38948 17836 46020 17864
rect 38948 17796 38976 17836
rect 46014 17824 46020 17836
rect 46072 17824 46078 17876
rect 48409 17867 48467 17873
rect 48409 17833 48421 17867
rect 48455 17864 48467 17867
rect 48498 17864 48504 17876
rect 48455 17836 48504 17864
rect 48455 17833 48467 17836
rect 48409 17827 48467 17833
rect 48498 17824 48504 17836
rect 48556 17824 48562 17876
rect 52825 17867 52883 17873
rect 52825 17864 52837 17867
rect 50724 17836 52837 17864
rect 31680 17768 35112 17796
rect 36740 17768 38976 17796
rect 39040 17768 39436 17796
rect 27264 17700 28948 17728
rect 20119 17632 23336 17660
rect 23385 17663 23443 17669
rect 20119 17629 20131 17632
rect 20073 17623 20131 17629
rect 23385 17629 23397 17663
rect 23431 17660 23443 17663
rect 23474 17660 23480 17672
rect 23431 17632 23480 17660
rect 23431 17629 23443 17632
rect 23385 17623 23443 17629
rect 16298 17552 16304 17604
rect 16356 17552 16362 17604
rect 19702 17592 19708 17604
rect 17236 17564 19708 17592
rect 17236 17524 17264 17564
rect 19702 17552 19708 17564
rect 19760 17552 19766 17604
rect 16040 17496 17264 17524
rect 17770 17484 17776 17536
rect 17828 17524 17834 17536
rect 20088 17524 20116 17623
rect 23474 17620 23480 17632
rect 23532 17620 23538 17672
rect 24946 17660 24952 17672
rect 24907 17632 24952 17660
rect 24946 17620 24952 17632
rect 25004 17620 25010 17672
rect 26145 17663 26203 17669
rect 26145 17629 26157 17663
rect 26191 17660 26203 17663
rect 26234 17660 26240 17672
rect 26191 17632 26240 17660
rect 26191 17629 26203 17632
rect 26145 17623 26203 17629
rect 26234 17620 26240 17632
rect 26292 17620 26298 17672
rect 26412 17663 26470 17669
rect 26412 17629 26424 17663
rect 26458 17660 26470 17663
rect 26694 17660 26700 17672
rect 26458 17632 26700 17660
rect 26458 17629 26470 17632
rect 26412 17623 26470 17629
rect 26694 17620 26700 17632
rect 26752 17620 26758 17672
rect 27890 17660 27896 17672
rect 27172 17632 27896 17660
rect 23658 17552 23664 17604
rect 23716 17592 23722 17604
rect 27172 17592 27200 17632
rect 27890 17620 27896 17632
rect 27948 17620 27954 17672
rect 28074 17660 28080 17672
rect 28035 17632 28080 17660
rect 28074 17620 28080 17632
rect 28132 17620 28138 17672
rect 28166 17620 28172 17672
rect 28224 17660 28230 17672
rect 28353 17663 28411 17669
rect 28353 17660 28365 17663
rect 28224 17632 28365 17660
rect 28224 17620 28230 17632
rect 28353 17629 28365 17632
rect 28399 17629 28411 17663
rect 28353 17623 28411 17629
rect 28450 17663 28508 17669
rect 28450 17629 28462 17663
rect 28496 17629 28508 17663
rect 28920 17660 28948 17700
rect 30466 17688 30472 17740
rect 30524 17728 30530 17740
rect 31680 17737 31708 17768
rect 31665 17731 31723 17737
rect 31665 17728 31677 17731
rect 30524 17700 31677 17728
rect 30524 17688 30530 17700
rect 31665 17697 31677 17700
rect 31711 17697 31723 17731
rect 31665 17691 31723 17697
rect 32309 17731 32367 17737
rect 32309 17697 32321 17731
rect 32355 17697 32367 17731
rect 32309 17691 32367 17697
rect 30561 17663 30619 17669
rect 30561 17660 30573 17663
rect 28920 17632 30573 17660
rect 28450 17623 28508 17629
rect 30561 17629 30573 17632
rect 30607 17660 30619 17663
rect 31202 17660 31208 17672
rect 30607 17632 31208 17660
rect 30607 17629 30619 17632
rect 30561 17623 30619 17629
rect 23716 17564 27200 17592
rect 23716 17552 23722 17564
rect 27246 17552 27252 17604
rect 27304 17592 27310 17604
rect 28261 17595 28319 17601
rect 28261 17592 28273 17595
rect 27304 17564 28273 17592
rect 27304 17552 27310 17564
rect 28261 17561 28273 17564
rect 28307 17561 28319 17595
rect 28261 17555 28319 17561
rect 28460 17592 28488 17623
rect 31202 17620 31208 17632
rect 31260 17620 31266 17672
rect 31386 17660 31392 17672
rect 31347 17632 31392 17660
rect 31386 17620 31392 17632
rect 31444 17620 31450 17672
rect 32324 17660 32352 17691
rect 32398 17688 32404 17740
rect 32456 17728 32462 17740
rect 33042 17728 33048 17740
rect 32456 17700 32501 17728
rect 32692 17700 33048 17728
rect 32456 17688 32462 17700
rect 32140 17632 32352 17660
rect 32494 17663 32552 17669
rect 32140 17604 32168 17632
rect 32494 17629 32506 17663
rect 32540 17629 32552 17663
rect 32494 17623 32552 17629
rect 32585 17663 32643 17669
rect 32585 17629 32597 17663
rect 32631 17660 32643 17663
rect 32692 17660 32720 17700
rect 33042 17688 33048 17700
rect 33100 17688 33106 17740
rect 33778 17688 33784 17740
rect 33836 17728 33842 17740
rect 33873 17731 33931 17737
rect 33873 17728 33885 17731
rect 33836 17700 33885 17728
rect 33836 17688 33842 17700
rect 33873 17697 33885 17700
rect 33919 17697 33931 17731
rect 33873 17691 33931 17697
rect 32631 17632 32720 17660
rect 32631 17629 32643 17632
rect 32585 17623 32643 17629
rect 30466 17592 30472 17604
rect 28460 17564 30472 17592
rect 17828 17496 20116 17524
rect 23569 17527 23627 17533
rect 17828 17484 17834 17496
rect 23569 17493 23581 17527
rect 23615 17524 23627 17527
rect 24854 17524 24860 17536
rect 23615 17496 24860 17524
rect 23615 17493 23627 17496
rect 23569 17487 23627 17493
rect 24854 17484 24860 17496
rect 24912 17484 24918 17536
rect 25038 17484 25044 17536
rect 25096 17524 25102 17536
rect 25096 17496 25141 17524
rect 25096 17484 25102 17496
rect 25774 17484 25780 17536
rect 25832 17524 25838 17536
rect 27525 17527 27583 17533
rect 27525 17524 27537 17527
rect 25832 17496 27537 17524
rect 25832 17484 25838 17496
rect 27525 17493 27537 17496
rect 27571 17493 27583 17527
rect 27525 17487 27583 17493
rect 27614 17484 27620 17536
rect 27672 17524 27678 17536
rect 28460 17524 28488 17564
rect 30466 17552 30472 17564
rect 30524 17552 30530 17604
rect 30650 17552 30656 17604
rect 30708 17592 30714 17604
rect 30837 17595 30895 17601
rect 30837 17592 30849 17595
rect 30708 17564 30849 17592
rect 30708 17552 30714 17564
rect 30837 17561 30849 17564
rect 30883 17561 30895 17595
rect 30837 17555 30895 17561
rect 27672 17496 28488 17524
rect 27672 17484 27678 17496
rect 29914 17484 29920 17536
rect 29972 17524 29978 17536
rect 30745 17527 30803 17533
rect 30745 17524 30757 17527
rect 29972 17496 30757 17524
rect 29972 17484 29978 17496
rect 30745 17493 30757 17496
rect 30791 17493 30803 17527
rect 30852 17524 30880 17555
rect 32122 17552 32128 17604
rect 32180 17552 32186 17604
rect 32508 17592 32536 17623
rect 34422 17620 34428 17672
rect 34480 17660 34486 17672
rect 35084 17669 35112 17768
rect 35158 17688 35164 17740
rect 35216 17728 35222 17740
rect 39040 17728 39068 17768
rect 35216 17700 39068 17728
rect 35216 17688 35222 17700
rect 39114 17688 39120 17740
rect 39172 17728 39178 17740
rect 39301 17731 39359 17737
rect 39301 17728 39313 17731
rect 39172 17700 39313 17728
rect 39172 17688 39178 17700
rect 39301 17697 39313 17700
rect 39347 17697 39359 17731
rect 39408 17728 39436 17768
rect 39408 17700 40448 17728
rect 39301 17691 39359 17697
rect 34885 17663 34943 17669
rect 34885 17660 34897 17663
rect 34480 17632 34897 17660
rect 34480 17620 34486 17632
rect 34885 17629 34897 17632
rect 34931 17629 34943 17663
rect 34885 17623 34943 17629
rect 35069 17663 35127 17669
rect 35069 17629 35081 17663
rect 35115 17629 35127 17663
rect 35250 17660 35256 17672
rect 35211 17632 35256 17660
rect 35069 17623 35127 17629
rect 35250 17620 35256 17632
rect 35308 17620 35314 17672
rect 38930 17620 38936 17672
rect 38988 17660 38994 17672
rect 40313 17663 40371 17669
rect 40313 17660 40325 17663
rect 38988 17632 40325 17660
rect 38988 17620 38994 17632
rect 40313 17629 40325 17632
rect 40359 17629 40371 17663
rect 40313 17623 40371 17629
rect 32858 17592 32864 17604
rect 32508 17564 32864 17592
rect 32508 17524 32536 17564
rect 32858 17552 32864 17564
rect 32916 17552 32922 17604
rect 33042 17552 33048 17604
rect 33100 17592 33106 17604
rect 33100 17564 33732 17592
rect 33100 17552 33106 17564
rect 33704 17536 33732 17564
rect 33870 17552 33876 17604
rect 33928 17592 33934 17604
rect 33928 17564 34468 17592
rect 33928 17552 33934 17564
rect 30852 17496 32536 17524
rect 30745 17487 30803 17493
rect 33226 17484 33232 17536
rect 33284 17524 33290 17536
rect 33321 17527 33379 17533
rect 33321 17524 33333 17527
rect 33284 17496 33333 17524
rect 33284 17484 33290 17496
rect 33321 17493 33333 17496
rect 33367 17493 33379 17527
rect 33686 17524 33692 17536
rect 33647 17496 33692 17524
rect 33321 17487 33379 17493
rect 33686 17484 33692 17496
rect 33744 17484 33750 17536
rect 33781 17527 33839 17533
rect 33781 17493 33793 17527
rect 33827 17524 33839 17527
rect 34330 17524 34336 17536
rect 33827 17496 34336 17524
rect 33827 17493 33839 17496
rect 33781 17487 33839 17493
rect 34330 17484 34336 17496
rect 34388 17484 34394 17536
rect 34440 17524 34468 17564
rect 34514 17552 34520 17604
rect 34572 17592 34578 17604
rect 40420 17592 40448 17700
rect 40586 17669 40592 17672
rect 40580 17660 40592 17669
rect 40547 17632 40592 17660
rect 40580 17623 40592 17632
rect 40586 17620 40592 17623
rect 40644 17620 40650 17672
rect 47857 17663 47915 17669
rect 47857 17660 47869 17663
rect 41386 17632 47869 17660
rect 41386 17592 41414 17632
rect 47857 17629 47869 17632
rect 47903 17629 47915 17663
rect 48222 17660 48228 17672
rect 48183 17632 48228 17660
rect 47857 17623 47915 17629
rect 48222 17620 48228 17632
rect 48280 17620 48286 17672
rect 48314 17620 48320 17672
rect 48372 17660 48378 17672
rect 50724 17669 50752 17836
rect 52825 17833 52837 17836
rect 52871 17864 52883 17867
rect 55582 17864 55588 17876
rect 52871 17836 55588 17864
rect 52871 17833 52883 17836
rect 52825 17827 52883 17833
rect 55582 17824 55588 17836
rect 55640 17824 55646 17876
rect 57054 17824 57060 17876
rect 57112 17864 57118 17876
rect 58253 17867 58311 17873
rect 58253 17864 58265 17867
rect 57112 17836 58265 17864
rect 57112 17824 57118 17836
rect 58253 17833 58265 17836
rect 58299 17833 58311 17867
rect 58253 17827 58311 17833
rect 54570 17756 54576 17808
rect 54628 17796 54634 17808
rect 54628 17768 55720 17796
rect 54628 17756 54634 17768
rect 55692 17737 55720 17768
rect 55677 17731 55735 17737
rect 55677 17697 55689 17731
rect 55723 17697 55735 17731
rect 55677 17691 55735 17697
rect 56502 17688 56508 17740
rect 56560 17728 56566 17740
rect 56873 17731 56931 17737
rect 56873 17728 56885 17731
rect 56560 17700 56885 17728
rect 56560 17688 56566 17700
rect 56873 17697 56885 17700
rect 56919 17697 56931 17731
rect 56873 17691 56931 17697
rect 50433 17663 50491 17669
rect 50433 17660 50445 17663
rect 48372 17632 50445 17660
rect 48372 17620 48378 17632
rect 50433 17629 50445 17632
rect 50479 17629 50491 17663
rect 50433 17623 50491 17629
rect 50709 17663 50767 17669
rect 50709 17629 50721 17663
rect 50755 17629 50767 17663
rect 50709 17623 50767 17629
rect 50801 17663 50859 17669
rect 50801 17629 50813 17663
rect 50847 17629 50859 17663
rect 50801 17623 50859 17629
rect 43070 17592 43076 17604
rect 34572 17564 40356 17592
rect 40420 17564 41414 17592
rect 41616 17564 43076 17592
rect 34572 17552 34578 17564
rect 39114 17524 39120 17536
rect 34440 17496 39120 17524
rect 39114 17484 39120 17496
rect 39172 17484 39178 17536
rect 39209 17527 39267 17533
rect 39209 17493 39221 17527
rect 39255 17524 39267 17527
rect 39666 17524 39672 17536
rect 39255 17496 39672 17524
rect 39255 17493 39267 17496
rect 39209 17487 39267 17493
rect 39666 17484 39672 17496
rect 39724 17484 39730 17536
rect 40328 17524 40356 17564
rect 41616 17524 41644 17564
rect 43070 17552 43076 17564
rect 43128 17552 43134 17604
rect 47670 17552 47676 17604
rect 47728 17592 47734 17604
rect 48041 17595 48099 17601
rect 48041 17592 48053 17595
rect 47728 17564 48053 17592
rect 47728 17552 47734 17564
rect 48041 17561 48053 17564
rect 48087 17561 48099 17595
rect 48041 17555 48099 17561
rect 48133 17595 48191 17601
rect 48133 17561 48145 17595
rect 48179 17592 48191 17595
rect 49602 17592 49608 17604
rect 48179 17564 49608 17592
rect 48179 17561 48191 17564
rect 48133 17555 48191 17561
rect 49602 17552 49608 17564
rect 49660 17552 49666 17604
rect 50614 17592 50620 17604
rect 50575 17564 50620 17592
rect 50614 17552 50620 17564
rect 50672 17552 50678 17604
rect 50816 17592 50844 17623
rect 51074 17620 51080 17672
rect 51132 17660 51138 17672
rect 51445 17663 51503 17669
rect 51445 17660 51457 17663
rect 51132 17632 51457 17660
rect 51132 17620 51138 17632
rect 51445 17629 51457 17632
rect 51491 17629 51503 17663
rect 52454 17660 52460 17672
rect 51445 17623 51503 17629
rect 51644 17632 52460 17660
rect 51644 17592 51672 17632
rect 52454 17620 52460 17632
rect 52512 17620 52518 17672
rect 54570 17620 54576 17672
rect 54628 17660 54634 17672
rect 55493 17663 55551 17669
rect 55493 17660 55505 17663
rect 54628 17632 55505 17660
rect 54628 17620 54634 17632
rect 55493 17629 55505 17632
rect 55539 17629 55551 17663
rect 58894 17660 58900 17672
rect 55493 17623 55551 17629
rect 55600 17632 58900 17660
rect 51718 17601 51724 17604
rect 50816 17564 51672 17592
rect 51712 17555 51724 17601
rect 51776 17592 51782 17604
rect 51776 17564 51812 17592
rect 51718 17552 51724 17555
rect 51776 17552 51782 17564
rect 52362 17552 52368 17604
rect 52420 17592 52426 17604
rect 55600 17592 55628 17632
rect 58894 17620 58900 17632
rect 58952 17620 58958 17672
rect 52420 17564 55628 17592
rect 52420 17552 52426 17564
rect 56134 17552 56140 17604
rect 56192 17592 56198 17604
rect 57118 17595 57176 17601
rect 57118 17592 57130 17595
rect 56192 17564 57130 17592
rect 56192 17552 56198 17564
rect 57118 17561 57130 17564
rect 57164 17561 57176 17595
rect 57118 17555 57176 17561
rect 40328 17496 41644 17524
rect 41693 17527 41751 17533
rect 41693 17493 41705 17527
rect 41739 17524 41751 17527
rect 41874 17524 41880 17536
rect 41739 17496 41880 17524
rect 41739 17493 41751 17496
rect 41693 17487 41751 17493
rect 41874 17484 41880 17496
rect 41932 17484 41938 17536
rect 50985 17527 51043 17533
rect 50985 17493 50997 17527
rect 51031 17524 51043 17527
rect 51534 17524 51540 17536
rect 51031 17496 51540 17524
rect 51031 17493 51043 17496
rect 50985 17487 51043 17493
rect 51534 17484 51540 17496
rect 51592 17484 51598 17536
rect 53098 17484 53104 17536
rect 53156 17524 53162 17536
rect 58342 17524 58348 17536
rect 53156 17496 58348 17524
rect 53156 17484 53162 17496
rect 58342 17484 58348 17496
rect 58400 17484 58406 17536
rect 1104 17434 58880 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 58880 17434
rect 1104 17360 58880 17382
rect 13722 17320 13728 17332
rect 13683 17292 13728 17320
rect 13722 17280 13728 17292
rect 13780 17280 13786 17332
rect 15378 17280 15384 17332
rect 15436 17320 15442 17332
rect 16574 17320 16580 17332
rect 15436 17292 16580 17320
rect 15436 17280 15442 17292
rect 16574 17280 16580 17292
rect 16632 17280 16638 17332
rect 16666 17280 16672 17332
rect 16724 17320 16730 17332
rect 21266 17320 21272 17332
rect 16724 17292 21272 17320
rect 16724 17280 16730 17292
rect 21266 17280 21272 17292
rect 21324 17280 21330 17332
rect 22646 17280 22652 17332
rect 22704 17320 22710 17332
rect 23201 17323 23259 17329
rect 23201 17320 23213 17323
rect 22704 17292 23213 17320
rect 22704 17280 22710 17292
rect 23201 17289 23213 17292
rect 23247 17289 23259 17323
rect 23201 17283 23259 17289
rect 26329 17323 26387 17329
rect 26329 17289 26341 17323
rect 26375 17320 26387 17323
rect 27338 17320 27344 17332
rect 26375 17292 27344 17320
rect 26375 17289 26387 17292
rect 26329 17283 26387 17289
rect 9861 17255 9919 17261
rect 6748 17224 8340 17252
rect 1581 17187 1639 17193
rect 1581 17153 1593 17187
rect 1627 17184 1639 17187
rect 2406 17184 2412 17196
rect 1627 17156 2412 17184
rect 1627 17153 1639 17156
rect 1581 17147 1639 17153
rect 2406 17144 2412 17156
rect 2464 17144 2470 17196
rect 6748 17193 6776 17224
rect 6733 17187 6791 17193
rect 6733 17153 6745 17187
rect 6779 17153 6791 17187
rect 8202 17184 8208 17196
rect 8163 17156 8208 17184
rect 6733 17147 6791 17153
rect 8202 17144 8208 17156
rect 8260 17144 8266 17196
rect 8312 17184 8340 17224
rect 9861 17221 9873 17255
rect 9907 17252 9919 17255
rect 9907 17224 24716 17252
rect 9907 17221 9919 17224
rect 9861 17215 9919 17221
rect 12526 17184 12532 17196
rect 8312 17156 12434 17184
rect 12487 17156 12532 17184
rect 1762 17116 1768 17128
rect 1723 17088 1768 17116
rect 1762 17076 1768 17088
rect 1820 17076 1826 17128
rect 6825 17119 6883 17125
rect 6825 17085 6837 17119
rect 6871 17085 6883 17119
rect 6825 17079 6883 17085
rect 6840 16980 6868 17079
rect 7006 17076 7012 17128
rect 7064 17116 7070 17128
rect 7101 17119 7159 17125
rect 7101 17116 7113 17119
rect 7064 17088 7113 17116
rect 7064 17076 7070 17088
rect 7101 17085 7113 17088
rect 7147 17085 7159 17119
rect 7101 17079 7159 17085
rect 8481 17119 8539 17125
rect 8481 17085 8493 17119
rect 8527 17116 8539 17119
rect 9766 17116 9772 17128
rect 8527 17088 9772 17116
rect 8527 17085 8539 17088
rect 8481 17079 8539 17085
rect 9766 17076 9772 17088
rect 9824 17076 9830 17128
rect 12406 17116 12434 17156
rect 12526 17144 12532 17156
rect 12584 17144 12590 17196
rect 15841 17187 15899 17193
rect 15841 17153 15853 17187
rect 15887 17184 15899 17187
rect 16114 17184 16120 17196
rect 15887 17156 16120 17184
rect 15887 17153 15899 17156
rect 15841 17147 15899 17153
rect 16114 17144 16120 17156
rect 16172 17144 16178 17196
rect 17037 17187 17095 17193
rect 17681 17187 17739 17193
rect 17037 17153 17049 17187
rect 17083 17159 17163 17187
rect 17083 17153 17095 17159
rect 17037 17147 17095 17153
rect 16390 17116 16396 17128
rect 12406 17088 16396 17116
rect 16390 17076 16396 17088
rect 16448 17076 16454 17128
rect 16758 17076 16764 17128
rect 16816 17116 16822 17128
rect 16853 17119 16911 17125
rect 16853 17116 16865 17119
rect 16816 17088 16865 17116
rect 16816 17076 16822 17088
rect 16853 17085 16865 17088
rect 16899 17085 16911 17119
rect 17135 17116 17163 17159
rect 17681 17153 17693 17187
rect 17727 17184 17739 17187
rect 20714 17184 20720 17196
rect 17727 17156 20720 17184
rect 17727 17153 17739 17156
rect 17681 17147 17739 17153
rect 20714 17144 20720 17156
rect 20772 17144 20778 17196
rect 21082 17184 21088 17196
rect 21043 17156 21088 17184
rect 21082 17144 21088 17156
rect 21140 17144 21146 17196
rect 21266 17144 21272 17196
rect 21324 17184 21330 17196
rect 22005 17187 22063 17193
rect 22005 17184 22017 17187
rect 21324 17156 22017 17184
rect 21324 17144 21330 17156
rect 22005 17153 22017 17156
rect 22051 17153 22063 17187
rect 24578 17184 24584 17196
rect 22005 17147 22063 17153
rect 23400 17156 24584 17184
rect 17135 17088 20760 17116
rect 16853 17079 16911 17085
rect 16209 17051 16267 17057
rect 16209 17017 16221 17051
rect 16255 17048 16267 17051
rect 17221 17051 17279 17057
rect 16255 17020 17172 17048
rect 16255 17017 16267 17020
rect 16209 17011 16267 17017
rect 9582 16980 9588 16992
rect 6840 16952 9588 16980
rect 9582 16940 9588 16952
rect 9640 16940 9646 16992
rect 15010 16940 15016 16992
rect 15068 16980 15074 16992
rect 16301 16983 16359 16989
rect 16301 16980 16313 16983
rect 15068 16952 16313 16980
rect 15068 16940 15074 16952
rect 16301 16949 16313 16952
rect 16347 16949 16359 16983
rect 17144 16980 17172 17020
rect 17221 17017 17233 17051
rect 17267 17048 17279 17051
rect 20438 17048 20444 17060
rect 17267 17020 20444 17048
rect 17267 17017 17279 17020
rect 17221 17011 17279 17017
rect 20438 17008 20444 17020
rect 20496 17008 20502 17060
rect 20732 17057 20760 17088
rect 20990 17076 20996 17128
rect 21048 17116 21054 17128
rect 21177 17119 21235 17125
rect 21177 17116 21189 17119
rect 21048 17088 21189 17116
rect 21048 17076 21054 17088
rect 21177 17085 21189 17088
rect 21223 17085 21235 17119
rect 21177 17079 21235 17085
rect 21361 17119 21419 17125
rect 21361 17085 21373 17119
rect 21407 17116 21419 17119
rect 23400 17116 23428 17156
rect 24578 17144 24584 17156
rect 24636 17144 24642 17196
rect 21407 17088 23428 17116
rect 24688 17116 24716 17224
rect 25222 17212 25228 17264
rect 25280 17261 25286 17264
rect 25280 17255 25329 17261
rect 25280 17221 25283 17255
rect 25317 17221 25329 17255
rect 25280 17215 25329 17221
rect 25280 17212 25286 17215
rect 25406 17212 25412 17264
rect 25464 17252 25470 17264
rect 25866 17252 25872 17264
rect 25464 17224 25872 17252
rect 25464 17212 25470 17224
rect 25866 17212 25872 17224
rect 25924 17252 25930 17264
rect 26344 17252 26372 17283
rect 27338 17280 27344 17292
rect 27396 17280 27402 17332
rect 31846 17320 31852 17332
rect 27632 17292 31852 17320
rect 25924 17224 26372 17252
rect 25924 17212 25930 17224
rect 25130 17184 25136 17196
rect 25091 17156 25136 17184
rect 25130 17144 25136 17156
rect 25188 17144 25194 17196
rect 25958 17144 25964 17196
rect 26016 17184 26022 17196
rect 26145 17187 26203 17193
rect 26145 17184 26157 17187
rect 26016 17156 26157 17184
rect 26016 17144 26022 17156
rect 26145 17153 26157 17156
rect 26191 17153 26203 17187
rect 26145 17147 26203 17153
rect 26283 17187 26341 17193
rect 26283 17153 26295 17187
rect 26329 17184 26341 17187
rect 26418 17184 26424 17196
rect 26329 17156 26424 17184
rect 26329 17153 26341 17156
rect 26283 17147 26341 17153
rect 26418 17144 26424 17156
rect 26476 17144 26482 17196
rect 26510 17144 26516 17196
rect 26568 17184 26574 17196
rect 27249 17187 27307 17193
rect 26568 17156 26613 17184
rect 26568 17144 26574 17156
rect 27249 17153 27261 17187
rect 27295 17184 27307 17187
rect 27522 17184 27528 17196
rect 27295 17156 27528 17184
rect 27295 17153 27307 17156
rect 27249 17147 27307 17153
rect 27522 17144 27528 17156
rect 27580 17144 27586 17196
rect 27632 17116 27660 17292
rect 31846 17280 31852 17292
rect 31904 17280 31910 17332
rect 33686 17280 33692 17332
rect 33744 17320 33750 17332
rect 38746 17320 38752 17332
rect 33744 17292 38752 17320
rect 33744 17280 33750 17292
rect 38746 17280 38752 17292
rect 38804 17280 38810 17332
rect 51718 17320 51724 17332
rect 51679 17292 51724 17320
rect 51718 17280 51724 17292
rect 51776 17280 51782 17332
rect 52270 17280 52276 17332
rect 52328 17320 52334 17332
rect 54662 17320 54668 17332
rect 52328 17292 54668 17320
rect 52328 17280 52334 17292
rect 54662 17280 54668 17292
rect 54720 17280 54726 17332
rect 54754 17280 54760 17332
rect 54812 17320 54818 17332
rect 55674 17320 55680 17332
rect 54812 17292 55680 17320
rect 54812 17280 54818 17292
rect 27798 17252 27804 17264
rect 27759 17224 27804 17252
rect 27798 17212 27804 17224
rect 27856 17212 27862 17264
rect 28350 17252 28356 17264
rect 28000 17224 28356 17252
rect 27709 17187 27767 17193
rect 27709 17153 27721 17187
rect 27755 17153 27767 17187
rect 27890 17184 27896 17196
rect 27851 17156 27896 17184
rect 27709 17147 27767 17153
rect 24688 17088 27660 17116
rect 27724 17116 27752 17147
rect 27890 17144 27896 17156
rect 27948 17144 27954 17196
rect 28000 17116 28028 17224
rect 28350 17212 28356 17224
rect 28408 17212 28414 17264
rect 28902 17252 28908 17264
rect 28863 17224 28908 17252
rect 28902 17212 28908 17224
rect 28960 17212 28966 17264
rect 29362 17252 29368 17264
rect 29017 17224 29368 17252
rect 28718 17193 28724 17196
rect 28537 17187 28595 17193
rect 28537 17184 28549 17187
rect 27724 17088 28028 17116
rect 28092 17156 28549 17184
rect 21407 17085 21419 17088
rect 21361 17079 21419 17085
rect 20717 17051 20775 17057
rect 20717 17017 20729 17051
rect 20763 17017 20775 17051
rect 21192 17048 21220 17079
rect 28092 17057 28120 17156
rect 28537 17153 28549 17156
rect 28583 17153 28595 17187
rect 28537 17147 28595 17153
rect 28685 17187 28724 17193
rect 28685 17153 28697 17187
rect 28685 17147 28724 17153
rect 28718 17144 28724 17147
rect 28776 17144 28782 17196
rect 28810 17144 28816 17196
rect 28868 17184 28874 17196
rect 29017 17193 29045 17224
rect 29362 17212 29368 17224
rect 29420 17252 29426 17264
rect 29638 17252 29644 17264
rect 29420 17224 29644 17252
rect 29420 17212 29426 17224
rect 29638 17212 29644 17224
rect 29696 17212 29702 17264
rect 30742 17212 30748 17264
rect 30800 17252 30806 17264
rect 31754 17252 31760 17264
rect 30800 17224 31760 17252
rect 30800 17212 30806 17224
rect 31754 17212 31760 17224
rect 31812 17212 31818 17264
rect 32582 17212 32588 17264
rect 32640 17212 32646 17264
rect 35250 17252 35256 17264
rect 32784 17224 35256 17252
rect 29002 17187 29060 17193
rect 28868 17156 28913 17184
rect 28868 17144 28874 17156
rect 29002 17153 29014 17187
rect 29048 17153 29060 17187
rect 29733 17187 29791 17193
rect 29733 17184 29745 17187
rect 29002 17147 29060 17153
rect 29196 17156 29745 17184
rect 25961 17051 26019 17057
rect 21192 17020 25912 17048
rect 20717 17011 20775 17017
rect 18138 16980 18144 16992
rect 17144 16952 18144 16980
rect 16301 16943 16359 16949
rect 18138 16940 18144 16952
rect 18196 16940 18202 16992
rect 18874 16980 18880 16992
rect 18835 16952 18880 16980
rect 18874 16940 18880 16952
rect 18932 16940 18938 16992
rect 20349 16983 20407 16989
rect 20349 16949 20361 16983
rect 20395 16980 20407 16983
rect 20990 16980 20996 16992
rect 20395 16952 20996 16980
rect 20395 16949 20407 16952
rect 20349 16943 20407 16949
rect 20990 16940 20996 16952
rect 21048 16940 21054 16992
rect 23658 16940 23664 16992
rect 23716 16980 23722 16992
rect 24118 16980 24124 16992
rect 23716 16952 24124 16980
rect 23716 16940 23722 16952
rect 24118 16940 24124 16952
rect 24176 16940 24182 16992
rect 24857 16983 24915 16989
rect 24857 16949 24869 16983
rect 24903 16980 24915 16983
rect 25590 16980 25596 16992
rect 24903 16952 25596 16980
rect 24903 16949 24915 16952
rect 24857 16943 24915 16949
rect 25590 16940 25596 16952
rect 25648 16940 25654 16992
rect 25884 16980 25912 17020
rect 25961 17017 25973 17051
rect 26007 17048 26019 17051
rect 28077 17051 28135 17057
rect 26007 17020 28028 17048
rect 26007 17017 26019 17020
rect 25961 17011 26019 17017
rect 26878 16980 26884 16992
rect 25884 16952 26884 16980
rect 26878 16940 26884 16952
rect 26936 16940 26942 16992
rect 28000 16980 28028 17020
rect 28077 17017 28089 17051
rect 28123 17017 28135 17051
rect 28077 17011 28135 17017
rect 28534 17008 28540 17060
rect 28592 17048 28598 17060
rect 29086 17048 29092 17060
rect 28592 17020 29092 17048
rect 28592 17008 28598 17020
rect 29086 17008 29092 17020
rect 29144 17008 29150 17060
rect 29196 17057 29224 17156
rect 29733 17153 29745 17156
rect 29779 17153 29791 17187
rect 30006 17184 30012 17196
rect 29967 17156 30012 17184
rect 29733 17147 29791 17153
rect 30006 17144 30012 17156
rect 30064 17144 30070 17196
rect 32600 17184 32628 17212
rect 32784 17193 32812 17224
rect 35250 17212 35256 17224
rect 35308 17212 35314 17264
rect 35986 17212 35992 17264
rect 36044 17252 36050 17264
rect 36044 17224 37274 17252
rect 36044 17212 36050 17224
rect 33962 17193 33968 17196
rect 32324 17156 32628 17184
rect 32769 17187 32827 17193
rect 29270 17076 29276 17128
rect 29328 17116 29334 17128
rect 29825 17119 29883 17125
rect 29825 17116 29837 17119
rect 29328 17088 29837 17116
rect 29328 17076 29334 17088
rect 29825 17085 29837 17088
rect 29871 17085 29883 17119
rect 29825 17079 29883 17085
rect 30469 17119 30527 17125
rect 30469 17085 30481 17119
rect 30515 17116 30527 17119
rect 31202 17116 31208 17128
rect 30515 17088 31208 17116
rect 30515 17085 30527 17088
rect 30469 17079 30527 17085
rect 31202 17076 31208 17088
rect 31260 17076 31266 17128
rect 32324 17125 32352 17156
rect 32769 17153 32781 17187
rect 32815 17153 32827 17187
rect 32769 17147 32827 17153
rect 33956 17147 33968 17193
rect 34020 17184 34026 17196
rect 37246 17184 37274 17224
rect 38562 17212 38568 17264
rect 38620 17252 38626 17264
rect 38620 17224 38665 17252
rect 38620 17212 38626 17224
rect 40310 17212 40316 17264
rect 40368 17252 40374 17264
rect 40678 17252 40684 17264
rect 40368 17224 40684 17252
rect 40368 17212 40374 17224
rect 40678 17212 40684 17224
rect 40736 17212 40742 17264
rect 40954 17252 40960 17264
rect 40915 17224 40960 17252
rect 40954 17212 40960 17224
rect 41012 17212 41018 17264
rect 41046 17212 41052 17264
rect 41104 17252 41110 17264
rect 41104 17224 41149 17252
rect 41104 17212 41110 17224
rect 41322 17212 41328 17264
rect 41380 17252 41386 17264
rect 52362 17252 52368 17264
rect 41380 17224 52368 17252
rect 41380 17212 41386 17224
rect 52362 17212 52368 17224
rect 52420 17212 52426 17264
rect 52454 17212 52460 17264
rect 52512 17252 52518 17264
rect 54956 17261 54984 17292
rect 55674 17280 55680 17292
rect 55732 17280 55738 17332
rect 56134 17320 56140 17332
rect 56095 17292 56140 17320
rect 56134 17280 56140 17292
rect 56192 17280 56198 17332
rect 57054 17280 57060 17332
rect 57112 17280 57118 17332
rect 54941 17255 54999 17261
rect 52512 17224 54892 17252
rect 52512 17212 52518 17224
rect 51166 17184 51172 17196
rect 34020 17156 34056 17184
rect 37246 17156 51172 17184
rect 33962 17144 33968 17147
rect 34020 17144 34026 17156
rect 51166 17144 51172 17156
rect 51224 17144 51230 17196
rect 51350 17184 51356 17196
rect 51311 17156 51356 17184
rect 51350 17144 51356 17156
rect 51408 17144 51414 17196
rect 51534 17184 51540 17196
rect 51495 17156 51540 17184
rect 51534 17144 51540 17156
rect 51592 17144 51598 17196
rect 54116 17177 54174 17183
rect 54116 17143 54128 17177
rect 54162 17143 54174 17177
rect 54294 17144 54300 17196
rect 54352 17184 54358 17196
rect 54757 17187 54815 17193
rect 54757 17184 54769 17187
rect 54352 17156 54769 17184
rect 54352 17144 54358 17156
rect 54757 17153 54769 17156
rect 54803 17153 54815 17187
rect 54864 17184 54892 17224
rect 54941 17221 54953 17255
rect 54987 17221 54999 17255
rect 54941 17215 54999 17221
rect 55033 17255 55091 17261
rect 55033 17221 55045 17255
rect 55079 17252 55091 17255
rect 57072 17252 57100 17280
rect 55079 17224 57100 17252
rect 55079 17221 55091 17224
rect 55033 17215 55091 17221
rect 55125 17187 55183 17193
rect 55125 17184 55137 17187
rect 54864 17156 55137 17184
rect 54757 17147 54815 17153
rect 55125 17153 55137 17156
rect 55171 17153 55183 17187
rect 55125 17147 55183 17153
rect 55953 17187 56011 17193
rect 55953 17153 55965 17187
rect 55999 17153 56011 17187
rect 55953 17147 56011 17153
rect 54116 17137 54174 17143
rect 32309 17119 32367 17125
rect 32309 17085 32321 17119
rect 32355 17085 32367 17119
rect 32309 17079 32367 17085
rect 32398 17076 32404 17128
rect 32456 17116 32462 17128
rect 32493 17119 32551 17125
rect 32493 17116 32505 17119
rect 32456 17088 32505 17116
rect 32456 17076 32462 17088
rect 32493 17085 32505 17088
rect 32539 17085 32551 17119
rect 32493 17079 32551 17085
rect 32585 17119 32643 17125
rect 32585 17085 32597 17119
rect 32631 17085 32643 17119
rect 32585 17079 32643 17085
rect 32677 17119 32735 17125
rect 32677 17085 32689 17119
rect 32723 17116 32735 17119
rect 32858 17116 32864 17128
rect 32723 17088 32864 17116
rect 32723 17085 32735 17088
rect 32677 17079 32735 17085
rect 29181 17051 29239 17057
rect 29181 17017 29193 17051
rect 29227 17017 29239 17051
rect 29181 17011 29239 17017
rect 32122 17008 32128 17060
rect 32180 17048 32186 17060
rect 32600 17048 32628 17079
rect 32858 17076 32864 17088
rect 32916 17076 32922 17128
rect 33134 17076 33140 17128
rect 33192 17116 33198 17128
rect 33689 17119 33747 17125
rect 33689 17116 33701 17119
rect 33192 17088 33701 17116
rect 33192 17076 33198 17088
rect 33689 17085 33701 17088
rect 33735 17085 33747 17119
rect 33689 17079 33747 17085
rect 38657 17119 38715 17125
rect 38657 17085 38669 17119
rect 38703 17116 38715 17119
rect 38746 17116 38752 17128
rect 38703 17088 38752 17116
rect 38703 17085 38715 17088
rect 38657 17079 38715 17085
rect 38746 17076 38752 17088
rect 38804 17076 38810 17128
rect 38838 17076 38844 17128
rect 38896 17116 38902 17128
rect 41233 17119 41291 17125
rect 38896 17088 38941 17116
rect 38896 17076 38902 17088
rect 41233 17085 41245 17119
rect 41279 17116 41291 17119
rect 43898 17116 43904 17128
rect 41279 17088 43904 17116
rect 41279 17085 41291 17088
rect 41233 17079 41291 17085
rect 43898 17076 43904 17088
rect 43956 17076 43962 17128
rect 51442 17076 51448 17128
rect 51500 17116 51506 17128
rect 52086 17116 52092 17128
rect 51500 17088 52092 17116
rect 51500 17076 51506 17088
rect 52086 17076 52092 17088
rect 52144 17116 52150 17128
rect 53926 17116 53932 17128
rect 52144 17088 53932 17116
rect 52144 17076 52150 17088
rect 53926 17076 53932 17088
rect 53984 17076 53990 17128
rect 38470 17048 38476 17060
rect 32180 17020 32628 17048
rect 34624 17020 38476 17048
rect 32180 17008 32186 17020
rect 34624 16980 34652 17020
rect 38470 17008 38476 17020
rect 38528 17008 38534 17060
rect 39298 17008 39304 17060
rect 39356 17048 39362 17060
rect 39482 17048 39488 17060
rect 39356 17020 39488 17048
rect 39356 17008 39362 17020
rect 39482 17008 39488 17020
rect 39540 17008 39546 17060
rect 39758 17008 39764 17060
rect 39816 17048 39822 17060
rect 48314 17048 48320 17060
rect 39816 17020 48320 17048
rect 39816 17008 39822 17020
rect 48314 17008 48320 17020
rect 48372 17008 48378 17060
rect 54128 16992 54156 17137
rect 55766 17116 55772 17128
rect 55727 17088 55772 17116
rect 55766 17076 55772 17088
rect 55824 17076 55830 17128
rect 55309 17051 55367 17057
rect 55309 17017 55321 17051
rect 55355 17048 55367 17051
rect 55968 17048 55996 17147
rect 56042 17144 56048 17196
rect 56100 17184 56106 17196
rect 57057 17187 57115 17193
rect 57057 17184 57069 17187
rect 56100 17156 57069 17184
rect 56100 17144 56106 17156
rect 57057 17153 57069 17156
rect 57103 17153 57115 17187
rect 57057 17147 57115 17153
rect 57330 17116 57336 17128
rect 57291 17088 57336 17116
rect 57330 17076 57336 17088
rect 57388 17076 57394 17128
rect 55355 17020 55996 17048
rect 55355 17017 55367 17020
rect 55309 17011 55367 17017
rect 28000 16952 34652 16980
rect 35069 16983 35127 16989
rect 35069 16949 35081 16983
rect 35115 16980 35127 16983
rect 35342 16980 35348 16992
rect 35115 16952 35348 16980
rect 35115 16949 35127 16952
rect 35069 16943 35127 16949
rect 35342 16940 35348 16952
rect 35400 16940 35406 16992
rect 38194 16980 38200 16992
rect 38155 16952 38200 16980
rect 38194 16940 38200 16952
rect 38252 16940 38258 16992
rect 39114 16940 39120 16992
rect 39172 16980 39178 16992
rect 40034 16980 40040 16992
rect 39172 16952 40040 16980
rect 39172 16940 39178 16952
rect 40034 16940 40040 16952
rect 40092 16940 40098 16992
rect 40589 16983 40647 16989
rect 40589 16949 40601 16983
rect 40635 16980 40647 16983
rect 44174 16980 44180 16992
rect 40635 16952 44180 16980
rect 40635 16949 40647 16952
rect 40589 16943 40647 16949
rect 44174 16940 44180 16952
rect 44232 16940 44238 16992
rect 54110 16940 54116 16992
rect 54168 16940 54174 16992
rect 54294 16980 54300 16992
rect 54255 16952 54300 16980
rect 54294 16940 54300 16952
rect 54352 16940 54358 16992
rect 1104 16890 58880 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 58880 16890
rect 1104 16816 58880 16838
rect 14274 16776 14280 16788
rect 11072 16748 14280 16776
rect 1578 16668 1584 16720
rect 1636 16708 1642 16720
rect 1636 16680 11008 16708
rect 1636 16668 1642 16680
rect 9398 16640 9404 16652
rect 9324 16612 9404 16640
rect 1581 16575 1639 16581
rect 1581 16541 1593 16575
rect 1627 16572 1639 16575
rect 7558 16572 7564 16584
rect 1627 16544 7564 16572
rect 1627 16541 1639 16544
rect 1581 16535 1639 16541
rect 7558 16532 7564 16544
rect 7616 16532 7622 16584
rect 9122 16572 9128 16584
rect 9083 16544 9128 16572
rect 9122 16532 9128 16544
rect 9180 16532 9186 16584
rect 9324 16581 9352 16612
rect 9398 16600 9404 16612
rect 9456 16600 9462 16652
rect 9309 16575 9367 16581
rect 9309 16541 9321 16575
rect 9355 16541 9367 16575
rect 10980 16572 11008 16680
rect 11072 16649 11100 16748
rect 14274 16736 14280 16748
rect 14332 16736 14338 16788
rect 26326 16776 26332 16788
rect 14752 16748 25636 16776
rect 13173 16711 13231 16717
rect 13173 16708 13185 16711
rect 12406 16680 13185 16708
rect 11057 16643 11115 16649
rect 11057 16609 11069 16643
rect 11103 16609 11115 16643
rect 11057 16603 11115 16609
rect 12406 16572 12434 16680
rect 13173 16677 13185 16680
rect 13219 16677 13231 16711
rect 14752 16708 14780 16748
rect 13173 16671 13231 16677
rect 13465 16680 14780 16708
rect 16117 16711 16175 16717
rect 13465 16649 13493 16680
rect 16117 16677 16129 16711
rect 16163 16677 16175 16711
rect 16117 16671 16175 16677
rect 13449 16643 13507 16649
rect 13449 16609 13461 16643
rect 13495 16609 13507 16643
rect 13449 16603 13507 16609
rect 13633 16643 13691 16649
rect 13633 16609 13645 16643
rect 13679 16640 13691 16643
rect 16132 16640 16160 16671
rect 16758 16668 16764 16720
rect 16816 16708 16822 16720
rect 17126 16708 17132 16720
rect 16816 16680 17132 16708
rect 16816 16668 16822 16680
rect 17126 16668 17132 16680
rect 17184 16708 17190 16720
rect 17402 16708 17408 16720
rect 17184 16680 17408 16708
rect 17184 16668 17190 16680
rect 17402 16668 17408 16680
rect 17460 16668 17466 16720
rect 22741 16711 22799 16717
rect 22741 16677 22753 16711
rect 22787 16708 22799 16711
rect 24581 16711 24639 16717
rect 22787 16680 24532 16708
rect 22787 16677 22799 16680
rect 22741 16671 22799 16677
rect 22281 16643 22339 16649
rect 13679 16612 13860 16640
rect 16132 16612 16712 16640
rect 13679 16609 13691 16612
rect 13633 16603 13691 16609
rect 10980 16544 12434 16572
rect 9309 16535 9367 16541
rect 12802 16532 12808 16584
rect 12860 16572 12866 16584
rect 13354 16572 13360 16584
rect 12860 16544 13032 16572
rect 13315 16544 13360 16572
rect 12860 16532 12866 16544
rect 1854 16504 1860 16516
rect 1815 16476 1860 16504
rect 1854 16464 1860 16476
rect 1912 16464 1918 16516
rect 11324 16507 11382 16513
rect 11324 16473 11336 16507
rect 11370 16504 11382 16507
rect 12894 16504 12900 16516
rect 11370 16476 12900 16504
rect 11370 16473 11382 16476
rect 11324 16467 11382 16473
rect 12894 16464 12900 16476
rect 12952 16464 12958 16516
rect 13004 16504 13032 16544
rect 13354 16532 13360 16544
rect 13412 16532 13418 16584
rect 13541 16575 13599 16581
rect 13541 16541 13553 16575
rect 13587 16572 13599 16575
rect 13722 16572 13728 16584
rect 13587 16544 13728 16572
rect 13587 16541 13599 16544
rect 13541 16535 13599 16541
rect 13722 16532 13728 16544
rect 13780 16532 13786 16584
rect 13832 16504 13860 16612
rect 14274 16532 14280 16584
rect 14332 16572 14338 16584
rect 14737 16575 14795 16581
rect 14737 16572 14749 16575
rect 14332 16544 14749 16572
rect 14332 16532 14338 16544
rect 14737 16541 14749 16544
rect 14783 16572 14795 16575
rect 16574 16572 16580 16584
rect 14783 16544 15148 16572
rect 16535 16544 16580 16572
rect 14783 16541 14795 16544
rect 14737 16535 14795 16541
rect 15010 16513 15016 16516
rect 15004 16504 15016 16513
rect 13004 16476 13860 16504
rect 14971 16476 15016 16504
rect 15004 16467 15016 16476
rect 15010 16464 15016 16467
rect 15068 16464 15074 16516
rect 15120 16504 15148 16544
rect 16574 16532 16580 16544
rect 16632 16532 16638 16584
rect 16684 16572 16712 16612
rect 22281 16609 22293 16643
rect 22327 16640 22339 16643
rect 22462 16640 22468 16652
rect 22327 16612 22468 16640
rect 22327 16609 22339 16612
rect 22281 16603 22339 16609
rect 22462 16600 22468 16612
rect 22520 16600 22526 16652
rect 23382 16640 23388 16652
rect 23343 16612 23388 16640
rect 23382 16600 23388 16612
rect 23440 16600 23446 16652
rect 23566 16600 23572 16652
rect 23624 16640 23630 16652
rect 24504 16640 24532 16680
rect 24581 16677 24593 16711
rect 24627 16708 24639 16711
rect 24762 16708 24768 16720
rect 24627 16680 24768 16708
rect 24627 16677 24639 16680
rect 24581 16671 24639 16677
rect 24762 16668 24768 16680
rect 24820 16668 24826 16720
rect 23624 16612 24072 16640
rect 24504 16612 25544 16640
rect 23624 16600 23630 16612
rect 19981 16575 20039 16581
rect 16684 16544 19932 16572
rect 16850 16504 16856 16516
rect 15120 16476 16856 16504
rect 16850 16464 16856 16476
rect 16908 16464 16914 16516
rect 19904 16504 19932 16544
rect 19981 16541 19993 16575
rect 20027 16572 20039 16575
rect 20070 16572 20076 16584
rect 20027 16544 20076 16572
rect 20027 16541 20039 16544
rect 19981 16535 20039 16541
rect 20070 16532 20076 16544
rect 20128 16532 20134 16584
rect 22186 16532 22192 16584
rect 22244 16572 22250 16584
rect 22830 16572 22836 16584
rect 22888 16581 22894 16584
rect 22888 16575 22924 16581
rect 22244 16544 22836 16572
rect 22244 16532 22250 16544
rect 22830 16532 22836 16544
rect 22912 16541 22924 16575
rect 23198 16572 23204 16584
rect 22888 16535 22924 16541
rect 23032 16544 23204 16572
rect 22888 16532 22894 16535
rect 21082 16504 21088 16516
rect 19904 16476 21088 16504
rect 21082 16464 21088 16476
rect 21140 16464 21146 16516
rect 23032 16513 23060 16544
rect 23198 16532 23204 16544
rect 23256 16532 23262 16584
rect 23293 16575 23351 16581
rect 23293 16541 23305 16575
rect 23339 16541 23351 16575
rect 23842 16572 23848 16584
rect 23803 16544 23848 16572
rect 23293 16535 23351 16541
rect 22991 16507 23060 16513
rect 22991 16473 23003 16507
rect 23037 16476 23060 16507
rect 23308 16504 23336 16535
rect 23842 16532 23848 16544
rect 23900 16532 23906 16584
rect 24044 16572 24072 16612
rect 24486 16572 24492 16584
rect 24044 16544 24492 16572
rect 24486 16532 24492 16544
rect 24544 16572 24550 16584
rect 24765 16575 24823 16581
rect 24765 16572 24777 16575
rect 24544 16544 24777 16572
rect 24544 16532 24550 16544
rect 24765 16541 24777 16544
rect 24811 16541 24823 16575
rect 24765 16535 24823 16541
rect 24854 16532 24860 16584
rect 24912 16572 24918 16584
rect 25133 16575 25191 16581
rect 25133 16572 25145 16575
rect 24912 16544 25145 16572
rect 24912 16532 24918 16544
rect 25133 16541 25145 16544
rect 25179 16541 25191 16575
rect 25133 16535 25191 16541
rect 23308 16476 24992 16504
rect 23037 16473 23049 16476
rect 22991 16467 23049 16473
rect 9306 16436 9312 16448
rect 9267 16408 9312 16436
rect 9306 16396 9312 16408
rect 9364 16396 9370 16448
rect 12437 16439 12495 16445
rect 12437 16405 12449 16439
rect 12483 16436 12495 16439
rect 16390 16436 16396 16448
rect 12483 16408 16396 16436
rect 12483 16405 12495 16408
rect 12437 16399 12495 16405
rect 16390 16396 16396 16408
rect 16448 16396 16454 16448
rect 16574 16396 16580 16448
rect 16632 16436 16638 16448
rect 16942 16436 16948 16448
rect 16632 16408 16948 16436
rect 16632 16396 16638 16408
rect 16942 16396 16948 16408
rect 17000 16396 17006 16448
rect 17954 16436 17960 16448
rect 17915 16408 17960 16436
rect 17954 16396 17960 16408
rect 18012 16396 18018 16448
rect 18046 16396 18052 16448
rect 18104 16436 18110 16448
rect 22278 16436 22284 16448
rect 18104 16408 22284 16436
rect 18104 16396 18110 16408
rect 22278 16396 22284 16408
rect 22336 16396 22342 16448
rect 23382 16396 23388 16448
rect 23440 16436 23446 16448
rect 23937 16439 23995 16445
rect 23937 16436 23949 16439
rect 23440 16408 23949 16436
rect 23440 16396 23446 16408
rect 23937 16405 23949 16408
rect 23983 16405 23995 16439
rect 24854 16436 24860 16448
rect 24815 16408 24860 16436
rect 23937 16399 23995 16405
rect 24854 16396 24860 16408
rect 24912 16396 24918 16448
rect 24964 16445 24992 16476
rect 24949 16439 25007 16445
rect 24949 16405 24961 16439
rect 24995 16436 25007 16439
rect 25038 16436 25044 16448
rect 24995 16408 25044 16436
rect 24995 16405 25007 16408
rect 24949 16399 25007 16405
rect 25038 16396 25044 16408
rect 25096 16436 25102 16448
rect 25406 16436 25412 16448
rect 25096 16408 25412 16436
rect 25096 16396 25102 16408
rect 25406 16396 25412 16408
rect 25464 16396 25470 16448
rect 25516 16436 25544 16612
rect 25608 16572 25636 16748
rect 25700 16748 26332 16776
rect 25700 16649 25728 16748
rect 26326 16736 26332 16748
rect 26384 16736 26390 16788
rect 26878 16736 26884 16788
rect 26936 16776 26942 16788
rect 28626 16776 28632 16788
rect 26936 16748 28632 16776
rect 26936 16736 26942 16748
rect 28626 16736 28632 16748
rect 28684 16736 28690 16788
rect 33134 16776 33140 16788
rect 32968 16748 33140 16776
rect 31662 16708 31668 16720
rect 26712 16680 31668 16708
rect 25685 16643 25743 16649
rect 25685 16609 25697 16643
rect 25731 16609 25743 16643
rect 25685 16603 25743 16609
rect 26712 16572 26740 16680
rect 31662 16668 31668 16680
rect 31720 16668 31726 16720
rect 27062 16600 27068 16652
rect 27120 16640 27126 16652
rect 27985 16643 28043 16649
rect 27985 16640 27997 16643
rect 27120 16612 27997 16640
rect 27120 16600 27126 16612
rect 27985 16609 27997 16612
rect 28031 16609 28043 16643
rect 27985 16603 28043 16609
rect 28169 16643 28227 16649
rect 28169 16609 28181 16643
rect 28215 16640 28227 16643
rect 28258 16640 28264 16652
rect 28215 16612 28264 16640
rect 28215 16609 28227 16612
rect 28169 16603 28227 16609
rect 28258 16600 28264 16612
rect 28316 16600 28322 16652
rect 28442 16600 28448 16652
rect 28500 16640 28506 16652
rect 28721 16643 28779 16649
rect 28721 16640 28733 16643
rect 28500 16612 28733 16640
rect 28500 16600 28506 16612
rect 28721 16609 28733 16612
rect 28767 16609 28779 16643
rect 28721 16603 28779 16609
rect 30006 16600 30012 16652
rect 30064 16640 30070 16652
rect 32968 16649 32996 16748
rect 33134 16736 33140 16748
rect 33192 16736 33198 16788
rect 33594 16736 33600 16788
rect 33652 16776 33658 16788
rect 35342 16776 35348 16788
rect 33652 16748 35348 16776
rect 33652 16736 33658 16748
rect 35342 16736 35348 16748
rect 35400 16736 35406 16788
rect 37384 16748 38654 16776
rect 32493 16643 32551 16649
rect 32493 16640 32505 16643
rect 30064 16612 32505 16640
rect 30064 16600 30070 16612
rect 32493 16609 32505 16612
rect 32539 16609 32551 16643
rect 32493 16603 32551 16609
rect 32953 16643 33011 16649
rect 32953 16609 32965 16643
rect 32999 16609 33011 16643
rect 32953 16603 33011 16609
rect 25608 16544 26740 16572
rect 26786 16532 26792 16584
rect 26844 16572 26850 16584
rect 27890 16572 27896 16584
rect 26844 16544 27660 16572
rect 27851 16544 27896 16572
rect 26844 16532 26850 16544
rect 25952 16507 26010 16513
rect 25952 16473 25964 16507
rect 25998 16504 26010 16507
rect 27632 16504 27660 16544
rect 27890 16532 27896 16544
rect 27948 16532 27954 16584
rect 28902 16572 28908 16584
rect 28863 16544 28908 16572
rect 28902 16532 28908 16544
rect 28960 16532 28966 16584
rect 32508 16572 32536 16603
rect 36078 16600 36084 16652
rect 36136 16640 36142 16652
rect 36722 16640 36728 16652
rect 36136 16612 36728 16640
rect 36136 16600 36142 16612
rect 36722 16600 36728 16612
rect 36780 16600 36786 16652
rect 37384 16649 37412 16748
rect 38626 16708 38654 16748
rect 39666 16736 39672 16788
rect 39724 16776 39730 16788
rect 52270 16776 52276 16788
rect 39724 16748 52276 16776
rect 39724 16736 39730 16748
rect 52270 16736 52276 16748
rect 52328 16736 52334 16788
rect 52365 16779 52423 16785
rect 52365 16745 52377 16779
rect 52411 16776 52423 16779
rect 52454 16776 52460 16788
rect 52411 16748 52460 16776
rect 52411 16745 52423 16748
rect 52365 16739 52423 16745
rect 52454 16736 52460 16748
rect 52512 16736 52518 16788
rect 56502 16776 56508 16788
rect 53576 16748 56508 16776
rect 38930 16708 38936 16720
rect 38626 16680 38936 16708
rect 38930 16668 38936 16680
rect 38988 16668 38994 16720
rect 39482 16668 39488 16720
rect 39540 16708 39546 16720
rect 42886 16708 42892 16720
rect 39540 16680 40908 16708
rect 39540 16668 39546 16680
rect 37369 16643 37427 16649
rect 37369 16640 37381 16643
rect 37200 16612 37381 16640
rect 33042 16572 33048 16584
rect 32508 16544 33048 16572
rect 33042 16532 33048 16544
rect 33100 16532 33106 16584
rect 33226 16581 33232 16584
rect 33220 16572 33232 16581
rect 33187 16544 33232 16572
rect 33220 16535 33232 16544
rect 33226 16532 33232 16535
rect 33284 16532 33290 16584
rect 36354 16532 36360 16584
rect 36412 16572 36418 16584
rect 37200 16572 37228 16612
rect 37369 16609 37381 16612
rect 37415 16609 37427 16643
rect 37369 16603 37427 16609
rect 38746 16600 38752 16652
rect 38804 16640 38810 16652
rect 40497 16643 40555 16649
rect 40497 16640 40509 16643
rect 38804 16612 40509 16640
rect 38804 16600 38810 16612
rect 40497 16609 40509 16612
rect 40543 16609 40555 16643
rect 40880 16640 40908 16680
rect 41708 16680 42892 16708
rect 41509 16643 41567 16649
rect 41509 16640 41521 16643
rect 40497 16603 40555 16609
rect 40604 16612 40816 16640
rect 40880 16612 41521 16640
rect 36412 16544 37228 16572
rect 37636 16575 37694 16581
rect 36412 16532 36418 16544
rect 37636 16541 37648 16575
rect 37682 16572 37694 16575
rect 38194 16572 38200 16584
rect 37682 16544 38200 16572
rect 37682 16541 37694 16544
rect 37636 16535 37694 16541
rect 38194 16532 38200 16544
rect 38252 16532 38258 16584
rect 30374 16504 30380 16516
rect 25998 16476 27568 16504
rect 27632 16476 30380 16504
rect 25998 16473 26010 16476
rect 25952 16467 26010 16473
rect 26234 16436 26240 16448
rect 25516 16408 26240 16436
rect 26234 16396 26240 16408
rect 26292 16396 26298 16448
rect 27062 16436 27068 16448
rect 27023 16408 27068 16436
rect 27062 16396 27068 16408
rect 27120 16396 27126 16448
rect 27540 16445 27568 16476
rect 30374 16464 30380 16476
rect 30432 16464 30438 16516
rect 32125 16507 32183 16513
rect 32125 16473 32137 16507
rect 32171 16504 32183 16507
rect 32214 16504 32220 16516
rect 32171 16476 32220 16504
rect 32171 16473 32183 16476
rect 32125 16467 32183 16473
rect 32214 16464 32220 16476
rect 32272 16464 32278 16516
rect 32309 16507 32367 16513
rect 32309 16473 32321 16507
rect 32355 16504 32367 16507
rect 32490 16504 32496 16516
rect 32355 16476 32496 16504
rect 32355 16473 32367 16476
rect 32309 16467 32367 16473
rect 32490 16464 32496 16476
rect 32548 16464 32554 16516
rect 36538 16504 36544 16516
rect 36499 16476 36544 16504
rect 36538 16464 36544 16476
rect 36596 16464 36602 16516
rect 27525 16439 27583 16445
rect 27525 16405 27537 16439
rect 27571 16405 27583 16439
rect 27525 16399 27583 16405
rect 28258 16396 28264 16448
rect 28316 16436 28322 16448
rect 28718 16436 28724 16448
rect 28316 16408 28724 16436
rect 28316 16396 28322 16408
rect 28718 16396 28724 16408
rect 28776 16396 28782 16448
rect 29086 16436 29092 16448
rect 29047 16408 29092 16436
rect 29086 16396 29092 16408
rect 29144 16396 29150 16448
rect 34330 16436 34336 16448
rect 34291 16408 34336 16436
rect 34330 16396 34336 16408
rect 34388 16396 34394 16448
rect 36173 16439 36231 16445
rect 36173 16405 36185 16439
rect 36219 16436 36231 16439
rect 36446 16436 36452 16448
rect 36219 16408 36452 16436
rect 36219 16405 36231 16408
rect 36173 16399 36231 16405
rect 36446 16396 36452 16408
rect 36504 16396 36510 16448
rect 36633 16439 36691 16445
rect 36633 16405 36645 16439
rect 36679 16436 36691 16439
rect 36722 16436 36728 16448
rect 36679 16408 36728 16436
rect 36679 16405 36691 16408
rect 36633 16399 36691 16405
rect 36722 16396 36728 16408
rect 36780 16396 36786 16448
rect 38378 16396 38384 16448
rect 38436 16436 38442 16448
rect 38654 16436 38660 16448
rect 38436 16408 38660 16436
rect 38436 16396 38442 16408
rect 38654 16396 38660 16408
rect 38712 16436 38718 16448
rect 38749 16439 38807 16445
rect 38749 16436 38761 16439
rect 38712 16408 38761 16436
rect 38712 16396 38718 16408
rect 38749 16405 38761 16408
rect 38795 16405 38807 16439
rect 40604 16436 40632 16612
rect 40788 16581 40816 16612
rect 41509 16609 41521 16612
rect 41555 16609 41567 16643
rect 41509 16603 41567 16609
rect 40681 16575 40739 16581
rect 40681 16541 40693 16575
rect 40727 16541 40739 16575
rect 40681 16535 40739 16541
rect 40773 16575 40831 16581
rect 40773 16541 40785 16575
rect 40819 16541 40831 16575
rect 40773 16535 40831 16541
rect 40696 16504 40724 16535
rect 40862 16532 40868 16584
rect 40920 16572 40926 16584
rect 40957 16575 41015 16581
rect 40957 16572 40969 16575
rect 40920 16544 40969 16572
rect 40920 16532 40926 16544
rect 40957 16541 40969 16544
rect 41003 16541 41015 16575
rect 40957 16535 41015 16541
rect 41046 16532 41052 16584
rect 41104 16572 41110 16584
rect 41708 16581 41736 16680
rect 42886 16668 42892 16680
rect 42944 16668 42950 16720
rect 41892 16612 42288 16640
rect 41693 16575 41751 16581
rect 41693 16572 41705 16575
rect 41104 16544 41149 16572
rect 41248 16544 41705 16572
rect 41104 16532 41110 16544
rect 41248 16516 41276 16544
rect 41693 16541 41705 16544
rect 41739 16541 41751 16575
rect 41693 16535 41751 16541
rect 41785 16575 41843 16581
rect 41785 16541 41797 16575
rect 41831 16572 41843 16575
rect 41892 16572 41920 16612
rect 41831 16544 41920 16572
rect 41969 16575 42027 16581
rect 41831 16541 41843 16544
rect 41785 16535 41843 16541
rect 41969 16541 41981 16575
rect 42015 16541 42027 16575
rect 41969 16535 42027 16541
rect 41230 16504 41236 16516
rect 40696 16476 41236 16504
rect 41230 16464 41236 16476
rect 41288 16464 41294 16516
rect 41322 16464 41328 16516
rect 41380 16504 41386 16516
rect 41414 16504 41420 16516
rect 41380 16476 41420 16504
rect 41380 16464 41386 16476
rect 41414 16464 41420 16476
rect 41472 16464 41478 16516
rect 41984 16504 42012 16535
rect 42058 16532 42064 16584
rect 42116 16572 42122 16584
rect 42260 16572 42288 16612
rect 42702 16600 42708 16652
rect 42760 16640 42766 16652
rect 44726 16640 44732 16652
rect 42760 16612 44732 16640
rect 42760 16600 42766 16612
rect 44726 16600 44732 16612
rect 44784 16600 44790 16652
rect 45186 16640 45192 16652
rect 45147 16612 45192 16640
rect 45186 16600 45192 16612
rect 45244 16600 45250 16652
rect 50614 16600 50620 16652
rect 50672 16640 50678 16652
rect 50982 16640 50988 16652
rect 50672 16612 50988 16640
rect 50672 16600 50678 16612
rect 50982 16600 50988 16612
rect 51040 16600 51046 16652
rect 52472 16640 52500 16736
rect 53576 16649 53604 16748
rect 56502 16736 56508 16748
rect 56560 16736 56566 16788
rect 54662 16668 54668 16720
rect 54720 16708 54726 16720
rect 58526 16708 58532 16720
rect 54720 16680 58532 16708
rect 54720 16668 54726 16680
rect 58526 16668 58532 16680
rect 58584 16668 58590 16720
rect 53009 16643 53067 16649
rect 52472 16612 52960 16640
rect 47118 16572 47124 16584
rect 42116 16544 42161 16572
rect 42260 16544 47124 16572
rect 42116 16532 42122 16544
rect 47118 16532 47124 16544
rect 47176 16532 47182 16584
rect 51350 16572 51356 16584
rect 51311 16544 51356 16572
rect 51350 16532 51356 16544
rect 51408 16532 51414 16584
rect 51534 16572 51540 16584
rect 51495 16544 51540 16572
rect 51534 16532 51540 16544
rect 51592 16532 51598 16584
rect 52932 16581 52960 16612
rect 53009 16609 53021 16643
rect 53055 16640 53067 16643
rect 53561 16643 53619 16649
rect 53055 16612 53512 16640
rect 53055 16609 53067 16612
rect 53009 16603 53067 16609
rect 52181 16575 52239 16581
rect 52181 16541 52193 16575
rect 52227 16572 52239 16575
rect 52917 16575 52975 16581
rect 52227 16544 52868 16572
rect 52227 16541 52239 16544
rect 52181 16535 52239 16541
rect 43162 16504 43168 16516
rect 41984 16476 43168 16504
rect 43162 16464 43168 16476
rect 43220 16464 43226 16516
rect 45456 16507 45514 16513
rect 45456 16473 45468 16507
rect 45502 16504 45514 16507
rect 46382 16504 46388 16516
rect 45502 16476 46388 16504
rect 45502 16473 45514 16476
rect 45456 16467 45514 16473
rect 46382 16464 46388 16476
rect 46440 16464 46446 16516
rect 47578 16464 47584 16516
rect 47636 16504 47642 16516
rect 52196 16504 52224 16535
rect 47636 16476 52224 16504
rect 47636 16464 47642 16476
rect 40862 16436 40868 16448
rect 40604 16408 40868 16436
rect 38749 16399 38807 16405
rect 40862 16396 40868 16408
rect 40920 16396 40926 16448
rect 46566 16436 46572 16448
rect 46527 16408 46572 16436
rect 46566 16396 46572 16408
rect 46624 16396 46630 16448
rect 51718 16436 51724 16448
rect 51679 16408 51724 16436
rect 51718 16396 51724 16408
rect 51776 16396 51782 16448
rect 52840 16436 52868 16544
rect 52917 16541 52929 16575
rect 52963 16541 52975 16575
rect 53098 16572 53104 16584
rect 53059 16544 53104 16572
rect 52917 16535 52975 16541
rect 53098 16532 53104 16544
rect 53156 16532 53162 16584
rect 53484 16504 53512 16612
rect 53561 16609 53573 16643
rect 53607 16609 53619 16643
rect 53561 16603 53619 16609
rect 53828 16575 53886 16581
rect 53828 16541 53840 16575
rect 53874 16572 53886 16575
rect 54294 16572 54300 16584
rect 53874 16544 54300 16572
rect 53874 16541 53886 16544
rect 53828 16535 53886 16541
rect 54294 16532 54300 16544
rect 54352 16532 54358 16584
rect 57974 16572 57980 16584
rect 57935 16544 57980 16572
rect 57974 16532 57980 16544
rect 58032 16532 58038 16584
rect 54570 16504 54576 16516
rect 53484 16476 54576 16504
rect 54570 16464 54576 16476
rect 54628 16464 54634 16516
rect 57054 16504 57060 16516
rect 54680 16476 56180 16504
rect 57015 16476 57060 16504
rect 54680 16436 54708 16476
rect 52840 16408 54708 16436
rect 54941 16439 54999 16445
rect 54941 16405 54953 16439
rect 54987 16436 54999 16439
rect 55214 16436 55220 16448
rect 54987 16408 55220 16436
rect 54987 16405 54999 16408
rect 54941 16399 54999 16405
rect 55214 16396 55220 16408
rect 55272 16436 55278 16448
rect 56042 16436 56048 16448
rect 55272 16408 56048 16436
rect 55272 16396 55278 16408
rect 56042 16396 56048 16408
rect 56100 16396 56106 16448
rect 56152 16436 56180 16476
rect 57054 16464 57060 16476
rect 57112 16464 57118 16516
rect 56962 16436 56968 16448
rect 56152 16408 56968 16436
rect 56962 16396 56968 16408
rect 57020 16396 57026 16448
rect 57146 16436 57152 16448
rect 57107 16408 57152 16436
rect 57146 16396 57152 16408
rect 57204 16396 57210 16448
rect 58066 16436 58072 16448
rect 58027 16408 58072 16436
rect 58066 16396 58072 16408
rect 58124 16396 58130 16448
rect 1104 16346 58880 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 58880 16346
rect 1104 16272 58880 16294
rect 13630 16192 13636 16244
rect 13688 16232 13694 16244
rect 15105 16235 15163 16241
rect 15105 16232 15117 16235
rect 13688 16204 15117 16232
rect 13688 16192 13694 16204
rect 15105 16201 15117 16204
rect 15151 16201 15163 16235
rect 15105 16195 15163 16201
rect 16209 16235 16267 16241
rect 16209 16201 16221 16235
rect 16255 16232 16267 16235
rect 16666 16232 16672 16244
rect 16255 16204 16672 16232
rect 16255 16201 16267 16204
rect 16209 16195 16267 16201
rect 16666 16192 16672 16204
rect 16724 16192 16730 16244
rect 19426 16192 19432 16244
rect 19484 16232 19490 16244
rect 19705 16235 19763 16241
rect 19705 16232 19717 16235
rect 19484 16204 19717 16232
rect 19484 16192 19490 16204
rect 19705 16201 19717 16204
rect 19751 16201 19763 16235
rect 19705 16195 19763 16201
rect 20438 16192 20444 16244
rect 20496 16232 20502 16244
rect 20496 16204 21772 16232
rect 20496 16192 20502 16204
rect 7558 16124 7564 16176
rect 7616 16164 7622 16176
rect 13078 16164 13084 16176
rect 7616 16136 13084 16164
rect 7616 16124 7622 16136
rect 13078 16124 13084 16136
rect 13136 16124 13142 16176
rect 14274 16164 14280 16176
rect 13188 16136 14280 16164
rect 1581 16099 1639 16105
rect 1581 16065 1593 16099
rect 1627 16096 1639 16099
rect 10134 16096 10140 16108
rect 1627 16068 2452 16096
rect 10095 16068 10140 16096
rect 1627 16065 1639 16068
rect 1581 16059 1639 16065
rect 2424 16040 2452 16068
rect 10134 16056 10140 16068
rect 10192 16056 10198 16108
rect 11882 16096 11888 16108
rect 11843 16068 11888 16096
rect 11882 16056 11888 16068
rect 11940 16056 11946 16108
rect 13188 16105 13216 16136
rect 14274 16124 14280 16136
rect 14332 16124 14338 16176
rect 17865 16167 17923 16173
rect 14384 16136 15516 16164
rect 13446 16105 13452 16108
rect 13173 16099 13231 16105
rect 13173 16065 13185 16099
rect 13219 16065 13231 16099
rect 13440 16096 13452 16105
rect 13407 16068 13452 16096
rect 13173 16059 13231 16065
rect 13440 16059 13452 16068
rect 13446 16056 13452 16059
rect 13504 16056 13510 16108
rect 13722 16056 13728 16108
rect 13780 16096 13786 16108
rect 14384 16096 14412 16136
rect 15378 16096 15384 16108
rect 13780 16068 14412 16096
rect 15339 16068 15384 16096
rect 13780 16056 13786 16068
rect 15378 16056 15384 16068
rect 15436 16056 15442 16108
rect 15488 16105 15516 16136
rect 17865 16133 17877 16167
rect 17911 16164 17923 16167
rect 19334 16164 19340 16176
rect 17911 16136 19340 16164
rect 17911 16133 17923 16136
rect 17865 16127 17923 16133
rect 19334 16124 19340 16136
rect 19392 16124 19398 16176
rect 21744 16164 21772 16204
rect 21818 16192 21824 16244
rect 21876 16232 21882 16244
rect 21876 16204 23888 16232
rect 21876 16192 21882 16204
rect 22250 16167 22308 16173
rect 22250 16164 22262 16167
rect 21284 16136 21680 16164
rect 21744 16136 22262 16164
rect 15473 16099 15531 16105
rect 15473 16065 15485 16099
rect 15519 16065 15531 16099
rect 16114 16096 16120 16108
rect 16075 16068 16120 16096
rect 15473 16059 15531 16065
rect 16114 16056 16120 16068
rect 16172 16056 16178 16108
rect 16298 16096 16304 16108
rect 16259 16068 16304 16096
rect 16298 16056 16304 16068
rect 16356 16056 16362 16108
rect 17678 16096 17684 16108
rect 17639 16068 17684 16096
rect 17678 16056 17684 16068
rect 17736 16056 17742 16108
rect 18509 16099 18567 16105
rect 18509 16065 18521 16099
rect 18555 16096 18567 16099
rect 19242 16096 19248 16108
rect 18555 16068 19248 16096
rect 18555 16065 18567 16068
rect 18509 16059 18567 16065
rect 19242 16056 19248 16068
rect 19300 16056 19306 16108
rect 21174 16096 21180 16108
rect 19352 16068 21180 16096
rect 1762 16028 1768 16040
rect 1723 16000 1768 16028
rect 1762 15988 1768 16000
rect 1820 15988 1826 16040
rect 2406 16028 2412 16040
rect 2367 16000 2412 16028
rect 2406 15988 2412 16000
rect 2464 15988 2470 16040
rect 9953 16031 10011 16037
rect 9953 15997 9965 16031
rect 9999 16028 10011 16031
rect 10042 16028 10048 16040
rect 9999 16000 10048 16028
rect 9999 15997 10011 16000
rect 9953 15991 10011 15997
rect 10042 15988 10048 16000
rect 10100 15988 10106 16040
rect 11977 16031 12035 16037
rect 11977 15997 11989 16031
rect 12023 16028 12035 16031
rect 12618 16028 12624 16040
rect 12023 16000 12624 16028
rect 12023 15997 12035 16000
rect 11977 15991 12035 15997
rect 12618 15988 12624 16000
rect 12676 15988 12682 16040
rect 15289 16031 15347 16037
rect 15289 15997 15301 16031
rect 15335 16028 15347 16031
rect 15335 16000 15424 16028
rect 15335 15997 15347 16000
rect 15289 15991 15347 15997
rect 15396 15960 15424 16000
rect 15562 15988 15568 16040
rect 15620 16028 15626 16040
rect 17957 16031 18015 16037
rect 15620 16000 15665 16028
rect 15620 15988 15626 16000
rect 17957 15997 17969 16031
rect 18003 16028 18015 16031
rect 19352 16028 19380 16068
rect 21174 16056 21180 16068
rect 21232 16056 21238 16108
rect 21284 16105 21312 16136
rect 21269 16099 21327 16105
rect 21269 16065 21281 16099
rect 21315 16065 21327 16099
rect 21450 16096 21456 16108
rect 21411 16068 21456 16096
rect 21269 16059 21327 16065
rect 21450 16056 21456 16068
rect 21508 16056 21514 16108
rect 21652 16096 21680 16136
rect 22250 16133 22262 16136
rect 22296 16133 22308 16167
rect 22250 16127 22308 16133
rect 22830 16124 22836 16176
rect 22888 16164 22894 16176
rect 23566 16164 23572 16176
rect 22888 16136 23572 16164
rect 22888 16124 22894 16136
rect 23566 16124 23572 16136
rect 23624 16124 23630 16176
rect 23382 16096 23388 16108
rect 21652 16068 23388 16096
rect 23382 16056 23388 16068
rect 23440 16056 23446 16108
rect 23860 16105 23888 16204
rect 24118 16192 24124 16244
rect 24176 16232 24182 16244
rect 27062 16232 27068 16244
rect 24176 16204 27068 16232
rect 24176 16192 24182 16204
rect 27062 16192 27068 16204
rect 27120 16192 27126 16244
rect 27249 16235 27307 16241
rect 27249 16201 27261 16235
rect 27295 16232 27307 16235
rect 28902 16232 28908 16244
rect 27295 16204 28908 16232
rect 27295 16201 27307 16204
rect 27249 16195 27307 16201
rect 28902 16192 28908 16204
rect 28960 16192 28966 16244
rect 30374 16192 30380 16244
rect 30432 16232 30438 16244
rect 37182 16232 37188 16244
rect 30432 16204 37188 16232
rect 30432 16192 30438 16204
rect 37182 16192 37188 16204
rect 37240 16192 37246 16244
rect 39482 16232 39488 16244
rect 37476 16204 39488 16232
rect 24210 16124 24216 16176
rect 24268 16164 24274 16176
rect 26786 16164 26792 16176
rect 24268 16136 26792 16164
rect 24268 16124 24274 16136
rect 26786 16124 26792 16136
rect 26844 16124 26850 16176
rect 27709 16167 27767 16173
rect 27709 16133 27721 16167
rect 27755 16164 27767 16167
rect 27890 16164 27896 16176
rect 27755 16136 27896 16164
rect 27755 16133 27767 16136
rect 27709 16127 27767 16133
rect 27890 16124 27896 16136
rect 27948 16124 27954 16176
rect 29270 16164 29276 16176
rect 28460 16136 29276 16164
rect 23845 16099 23903 16105
rect 23845 16065 23857 16099
rect 23891 16096 23903 16099
rect 27617 16099 27675 16105
rect 27617 16096 27629 16099
rect 23891 16068 27629 16096
rect 23891 16065 23903 16068
rect 23845 16059 23903 16065
rect 27617 16065 27629 16068
rect 27663 16096 27675 16099
rect 28258 16096 28264 16108
rect 27663 16068 28264 16096
rect 27663 16065 27675 16068
rect 27617 16059 27675 16065
rect 28258 16056 28264 16068
rect 28316 16056 28322 16108
rect 28460 16105 28488 16136
rect 29270 16124 29276 16136
rect 29328 16164 29334 16176
rect 29454 16164 29460 16176
rect 29328 16136 29460 16164
rect 29328 16124 29334 16136
rect 29454 16124 29460 16136
rect 29512 16124 29518 16176
rect 30466 16164 30472 16176
rect 30427 16136 30472 16164
rect 30466 16124 30472 16136
rect 30524 16124 30530 16176
rect 37476 16173 37504 16204
rect 39482 16192 39488 16204
rect 39540 16192 39546 16244
rect 40405 16235 40463 16241
rect 40405 16201 40417 16235
rect 40451 16232 40463 16235
rect 41046 16232 41052 16244
rect 40451 16204 41052 16232
rect 40451 16201 40463 16204
rect 40405 16195 40463 16201
rect 41046 16192 41052 16204
rect 41104 16192 41110 16244
rect 42058 16192 42064 16244
rect 42116 16232 42122 16244
rect 43162 16232 43168 16244
rect 42116 16204 43024 16232
rect 43123 16204 43168 16232
rect 42116 16192 42122 16204
rect 37461 16167 37519 16173
rect 37461 16133 37473 16167
rect 37507 16133 37519 16167
rect 37461 16127 37519 16133
rect 38473 16167 38531 16173
rect 38473 16133 38485 16167
rect 38519 16164 38531 16167
rect 38746 16164 38752 16176
rect 38519 16136 38752 16164
rect 38519 16133 38531 16136
rect 38473 16127 38531 16133
rect 38746 16124 38752 16136
rect 38804 16124 38810 16176
rect 38838 16124 38844 16176
rect 38896 16164 38902 16176
rect 39025 16167 39083 16173
rect 39025 16164 39037 16167
rect 38896 16136 39037 16164
rect 38896 16124 38902 16136
rect 39025 16133 39037 16136
rect 39071 16133 39083 16167
rect 40126 16164 40132 16176
rect 40087 16136 40132 16164
rect 39025 16127 39083 16133
rect 40126 16124 40132 16136
rect 40184 16124 40190 16176
rect 42150 16164 42156 16176
rect 40696 16136 42156 16164
rect 28445 16099 28503 16105
rect 28445 16065 28457 16099
rect 28491 16065 28503 16099
rect 28445 16059 28503 16065
rect 28712 16099 28770 16105
rect 28712 16065 28724 16099
rect 28758 16096 28770 16099
rect 29730 16096 29736 16108
rect 28758 16068 29736 16096
rect 28758 16065 28770 16068
rect 28712 16059 28770 16065
rect 29730 16056 29736 16068
rect 29788 16056 29794 16108
rect 30285 16099 30343 16105
rect 30285 16065 30297 16099
rect 30331 16096 30343 16099
rect 30374 16096 30380 16108
rect 30331 16068 30380 16096
rect 30331 16065 30343 16068
rect 30285 16059 30343 16065
rect 30374 16056 30380 16068
rect 30432 16056 30438 16108
rect 32398 16096 32404 16108
rect 32359 16068 32404 16096
rect 32398 16056 32404 16068
rect 32456 16056 32462 16108
rect 32582 16096 32588 16108
rect 32543 16068 32588 16096
rect 32582 16056 32588 16068
rect 32640 16056 32646 16108
rect 32674 16056 32680 16108
rect 32732 16096 32738 16108
rect 32861 16099 32919 16105
rect 32732 16068 32777 16096
rect 32732 16056 32738 16068
rect 32861 16065 32873 16099
rect 32907 16065 32919 16099
rect 32861 16059 32919 16065
rect 32953 16099 33011 16105
rect 32953 16065 32965 16099
rect 32999 16065 33011 16099
rect 32953 16059 33011 16065
rect 18003 16000 19380 16028
rect 18003 15997 18015 16000
rect 17957 15991 18015 15997
rect 19426 15988 19432 16040
rect 19484 16028 19490 16040
rect 21818 16028 21824 16040
rect 19484 16000 21824 16028
rect 19484 15988 19490 16000
rect 21818 15988 21824 16000
rect 21876 15988 21882 16040
rect 22002 16028 22008 16040
rect 21963 16000 22008 16028
rect 22002 15988 22008 16000
rect 22060 15988 22066 16040
rect 24854 15988 24860 16040
rect 24912 16028 24918 16040
rect 27706 16028 27712 16040
rect 24912 16000 27712 16028
rect 24912 15988 24918 16000
rect 27706 15988 27712 16000
rect 27764 15988 27770 16040
rect 27893 16031 27951 16037
rect 27893 15997 27905 16031
rect 27939 16028 27951 16031
rect 27982 16028 27988 16040
rect 27939 16000 27988 16028
rect 27939 15997 27951 16000
rect 27893 15991 27951 15997
rect 27982 15988 27988 16000
rect 28040 15988 28046 16040
rect 29546 15988 29552 16040
rect 29604 16028 29610 16040
rect 30653 16031 30711 16037
rect 30653 16028 30665 16031
rect 29604 16000 30665 16028
rect 29604 15988 29610 16000
rect 30653 15997 30665 16000
rect 30699 15997 30711 16031
rect 30653 15991 30711 15997
rect 31294 15988 31300 16040
rect 31352 16028 31358 16040
rect 32876 16028 32904 16059
rect 31352 16000 32904 16028
rect 32968 16028 32996 16059
rect 33042 16056 33048 16108
rect 33100 16096 33106 16108
rect 37645 16099 37703 16105
rect 37645 16096 37657 16099
rect 33100 16068 37657 16096
rect 33100 16056 33106 16068
rect 37645 16065 37657 16068
rect 37691 16096 37703 16099
rect 38657 16099 38715 16105
rect 38657 16096 38669 16099
rect 37691 16068 38669 16096
rect 37691 16065 37703 16068
rect 37645 16059 37703 16065
rect 38657 16065 38669 16068
rect 38703 16065 38715 16099
rect 38657 16059 38715 16065
rect 39758 16056 39764 16108
rect 39816 16096 39822 16108
rect 39853 16099 39911 16105
rect 39853 16096 39865 16099
rect 39816 16068 39865 16096
rect 39816 16056 39822 16068
rect 39853 16065 39865 16068
rect 39899 16065 39911 16099
rect 39853 16059 39911 16065
rect 40037 16099 40095 16105
rect 40037 16065 40049 16099
rect 40083 16065 40095 16099
rect 40037 16059 40095 16065
rect 40221 16099 40279 16105
rect 40221 16065 40233 16099
rect 40267 16096 40279 16099
rect 40586 16096 40592 16108
rect 40267 16068 40592 16096
rect 40267 16065 40279 16068
rect 40221 16059 40279 16065
rect 36998 16028 37004 16040
rect 32968 16000 37004 16028
rect 31352 15988 31358 16000
rect 36998 15988 37004 16000
rect 37056 15988 37062 16040
rect 38838 15988 38844 16040
rect 38896 16028 38902 16040
rect 40052 16028 40080 16059
rect 40586 16056 40592 16068
rect 40644 16056 40650 16108
rect 40696 16028 40724 16136
rect 41509 16099 41567 16105
rect 41509 16065 41521 16099
rect 41555 16096 41567 16099
rect 41690 16096 41696 16108
rect 41555 16068 41696 16096
rect 41555 16065 41567 16068
rect 41509 16059 41567 16065
rect 41690 16056 41696 16068
rect 41748 16056 41754 16108
rect 41984 16105 42012 16136
rect 42150 16124 42156 16136
rect 42208 16164 42214 16176
rect 42886 16164 42892 16176
rect 42208 16136 42748 16164
rect 42847 16136 42892 16164
rect 42208 16124 42214 16136
rect 41877 16099 41935 16105
rect 41877 16065 41889 16099
rect 41923 16065 41935 16099
rect 41877 16059 41935 16065
rect 41969 16099 42027 16105
rect 41969 16065 41981 16099
rect 42015 16065 42027 16099
rect 41969 16059 42027 16065
rect 42613 16099 42671 16105
rect 42613 16065 42625 16099
rect 42659 16065 42671 16099
rect 42720 16096 42748 16136
rect 42886 16124 42892 16136
rect 42944 16124 42950 16176
rect 42996 16164 43024 16204
rect 43162 16192 43168 16204
rect 43220 16192 43226 16244
rect 45370 16192 45376 16244
rect 45428 16232 45434 16244
rect 45465 16235 45523 16241
rect 45465 16232 45477 16235
rect 45428 16204 45477 16232
rect 45428 16192 45434 16204
rect 45465 16201 45477 16204
rect 45511 16201 45523 16235
rect 46382 16232 46388 16244
rect 46343 16204 46388 16232
rect 45465 16195 45523 16201
rect 46382 16192 46388 16204
rect 46440 16192 46446 16244
rect 46566 16192 46572 16244
rect 46624 16232 46630 16244
rect 46845 16235 46903 16241
rect 46845 16232 46857 16235
rect 46624 16204 46857 16232
rect 46624 16192 46630 16204
rect 46845 16201 46857 16204
rect 46891 16201 46903 16235
rect 46845 16195 46903 16201
rect 48133 16235 48191 16241
rect 48133 16201 48145 16235
rect 48179 16232 48191 16235
rect 53742 16232 53748 16244
rect 48179 16204 53748 16232
rect 48179 16201 48191 16204
rect 48133 16195 48191 16201
rect 53742 16192 53748 16204
rect 53800 16192 53806 16244
rect 54110 16232 54116 16244
rect 54071 16204 54116 16232
rect 54110 16192 54116 16204
rect 54168 16192 54174 16244
rect 54754 16232 54760 16244
rect 54715 16204 54760 16232
rect 54754 16192 54760 16204
rect 54812 16192 54818 16244
rect 51252 16167 51310 16173
rect 42996 16136 51212 16164
rect 42797 16099 42855 16105
rect 42797 16096 42809 16099
rect 42720 16068 42809 16096
rect 42613 16059 42671 16065
rect 42797 16065 42809 16068
rect 42843 16065 42855 16099
rect 42797 16059 42855 16065
rect 42981 16099 43039 16105
rect 42981 16065 42993 16099
rect 43027 16065 43039 16099
rect 44174 16096 44180 16108
rect 44135 16068 44180 16096
rect 42981 16059 43039 16065
rect 41598 16028 41604 16040
rect 38896 16000 40724 16028
rect 41559 16000 41604 16028
rect 38896 15988 38902 16000
rect 41598 15988 41604 16000
rect 41656 15988 41662 16040
rect 41892 16028 41920 16059
rect 42518 16028 42524 16040
rect 41892 16000 42524 16028
rect 42518 15988 42524 16000
rect 42576 15988 42582 16040
rect 14108 15932 15424 15960
rect 9858 15852 9864 15904
rect 9916 15892 9922 15904
rect 10321 15895 10379 15901
rect 10321 15892 10333 15895
rect 9916 15864 10333 15892
rect 9916 15852 9922 15864
rect 10321 15861 10333 15864
rect 10367 15861 10379 15895
rect 12250 15892 12256 15904
rect 12211 15864 12256 15892
rect 10321 15855 10379 15861
rect 12250 15852 12256 15864
rect 12308 15852 12314 15904
rect 13354 15852 13360 15904
rect 13412 15892 13418 15904
rect 14108 15892 14136 15932
rect 13412 15864 14136 15892
rect 14553 15895 14611 15901
rect 13412 15852 13418 15864
rect 14553 15861 14565 15895
rect 14599 15892 14611 15895
rect 14918 15892 14924 15904
rect 14599 15864 14924 15892
rect 14599 15861 14611 15864
rect 14553 15855 14611 15861
rect 14918 15852 14924 15864
rect 14976 15852 14982 15904
rect 15396 15892 15424 15932
rect 16850 15920 16856 15972
rect 16908 15960 16914 15972
rect 17405 15963 17463 15969
rect 17405 15960 17417 15963
rect 16908 15932 17417 15960
rect 16908 15920 16914 15932
rect 17405 15929 17417 15932
rect 17451 15929 17463 15963
rect 20898 15960 20904 15972
rect 17405 15923 17463 15929
rect 17512 15932 20904 15960
rect 17512 15892 17540 15932
rect 20898 15920 20904 15932
rect 20956 15920 20962 15972
rect 21082 15920 21088 15972
rect 21140 15960 21146 15972
rect 21140 15932 21404 15960
rect 21140 15920 21146 15932
rect 15396 15864 17540 15892
rect 17862 15852 17868 15904
rect 17920 15892 17926 15904
rect 19610 15892 19616 15904
rect 17920 15864 19616 15892
rect 17920 15852 17926 15864
rect 19610 15852 19616 15864
rect 19668 15852 19674 15904
rect 20070 15852 20076 15904
rect 20128 15892 20134 15904
rect 21269 15895 21327 15901
rect 21269 15892 21281 15895
rect 20128 15864 21281 15892
rect 20128 15852 20134 15864
rect 21269 15861 21281 15864
rect 21315 15861 21327 15895
rect 21376 15892 21404 15932
rect 23474 15920 23480 15972
rect 23532 15960 23538 15972
rect 24026 15960 24032 15972
rect 23532 15932 24032 15960
rect 23532 15920 23538 15932
rect 24026 15920 24032 15932
rect 24084 15920 24090 15972
rect 29454 15920 29460 15972
rect 29512 15960 29518 15972
rect 42058 15960 42064 15972
rect 29512 15932 42064 15960
rect 29512 15920 29518 15932
rect 42058 15920 42064 15932
rect 42116 15920 42122 15972
rect 23385 15895 23443 15901
rect 23385 15892 23397 15895
rect 21376 15864 23397 15892
rect 21269 15855 21327 15861
rect 23385 15861 23397 15864
rect 23431 15861 23443 15895
rect 23385 15855 23443 15861
rect 23566 15852 23572 15904
rect 23624 15892 23630 15904
rect 25041 15895 25099 15901
rect 25041 15892 25053 15895
rect 23624 15864 25053 15892
rect 23624 15852 23630 15864
rect 25041 15861 25053 15864
rect 25087 15861 25099 15895
rect 25041 15855 25099 15861
rect 27706 15852 27712 15904
rect 27764 15892 27770 15904
rect 29825 15895 29883 15901
rect 29825 15892 29837 15895
rect 27764 15864 29837 15892
rect 27764 15852 27770 15864
rect 29825 15861 29837 15864
rect 29871 15892 29883 15895
rect 30006 15892 30012 15904
rect 29871 15864 30012 15892
rect 29871 15861 29883 15864
rect 29825 15855 29883 15861
rect 30006 15852 30012 15864
rect 30064 15852 30070 15904
rect 31018 15852 31024 15904
rect 31076 15892 31082 15904
rect 35986 15892 35992 15904
rect 31076 15864 35992 15892
rect 31076 15852 31082 15864
rect 35986 15852 35992 15864
rect 36044 15852 36050 15904
rect 37182 15852 37188 15904
rect 37240 15892 37246 15904
rect 37737 15895 37795 15901
rect 37737 15892 37749 15895
rect 37240 15864 37749 15892
rect 37240 15852 37246 15864
rect 37737 15861 37749 15864
rect 37783 15861 37795 15895
rect 40954 15892 40960 15904
rect 40915 15864 40960 15892
rect 37737 15855 37795 15861
rect 40954 15852 40960 15864
rect 41012 15852 41018 15904
rect 42628 15892 42656 16059
rect 42886 15988 42892 16040
rect 42944 16028 42950 16040
rect 42996 16028 43024 16059
rect 44174 16056 44180 16068
rect 44232 16056 44238 16108
rect 46750 16096 46756 16108
rect 46711 16068 46756 16096
rect 46750 16056 46756 16068
rect 46808 16056 46814 16108
rect 51074 16096 51080 16108
rect 46952 16068 48360 16096
rect 42944 16000 43024 16028
rect 42944 15988 42950 16000
rect 43254 15988 43260 16040
rect 43312 16028 43318 16040
rect 46566 16028 46572 16040
rect 43312 16000 46572 16028
rect 43312 15988 43318 16000
rect 46566 15988 46572 16000
rect 46624 16028 46630 16040
rect 46952 16037 46980 16068
rect 46937 16031 46995 16037
rect 46937 16028 46949 16031
rect 46624 16000 46949 16028
rect 46624 15988 46630 16000
rect 46937 15997 46949 16000
rect 46983 15997 46995 16031
rect 48222 16028 48228 16040
rect 48183 16000 48228 16028
rect 46937 15991 46995 15997
rect 48222 15988 48228 16000
rect 48280 15988 48286 16040
rect 48332 16037 48360 16068
rect 51000 16068 51080 16096
rect 51000 16037 51028 16068
rect 51074 16056 51080 16068
rect 51132 16056 51138 16108
rect 51184 16096 51212 16136
rect 51252 16133 51264 16167
rect 51298 16164 51310 16167
rect 51718 16164 51724 16176
rect 51298 16136 51724 16164
rect 51298 16133 51310 16136
rect 51252 16127 51310 16133
rect 51718 16124 51724 16136
rect 51776 16124 51782 16176
rect 53837 16167 53895 16173
rect 53837 16133 53849 16167
rect 53883 16164 53895 16167
rect 55214 16164 55220 16176
rect 53883 16136 55220 16164
rect 53883 16133 53895 16136
rect 53837 16127 53895 16133
rect 55214 16124 55220 16136
rect 55272 16124 55278 16176
rect 53561 16099 53619 16105
rect 53561 16096 53573 16099
rect 51184 16068 53573 16096
rect 53561 16065 53573 16068
rect 53607 16065 53619 16099
rect 53561 16059 53619 16065
rect 53745 16099 53803 16105
rect 53745 16065 53757 16099
rect 53791 16065 53803 16099
rect 53926 16096 53932 16108
rect 53887 16068 53932 16096
rect 53745 16059 53803 16065
rect 48317 16031 48375 16037
rect 48317 15997 48329 16031
rect 48363 15997 48375 16031
rect 48317 15991 48375 15997
rect 50985 16031 51043 16037
rect 50985 15997 50997 16031
rect 51031 15997 51043 16031
rect 50985 15991 51043 15997
rect 53760 16028 53788 16059
rect 53926 16056 53932 16068
rect 53984 16096 53990 16108
rect 54386 16096 54392 16108
rect 53984 16068 54392 16096
rect 53984 16056 53990 16068
rect 54386 16056 54392 16068
rect 54444 16056 54450 16108
rect 54570 16096 54576 16108
rect 54531 16068 54576 16096
rect 54570 16056 54576 16068
rect 54628 16056 54634 16108
rect 54754 16028 54760 16040
rect 53760 16000 54760 16028
rect 48130 15920 48136 15972
rect 48188 15960 48194 15972
rect 51000 15960 51028 15991
rect 53760 15960 53788 16000
rect 54754 15988 54760 16000
rect 54812 15988 54818 16040
rect 48188 15932 51028 15960
rect 51920 15932 53788 15960
rect 48188 15920 48194 15932
rect 47210 15892 47216 15904
rect 42628 15864 47216 15892
rect 47210 15852 47216 15864
rect 47268 15852 47274 15904
rect 47762 15892 47768 15904
rect 47723 15864 47768 15892
rect 47762 15852 47768 15864
rect 47820 15852 47826 15904
rect 51166 15852 51172 15904
rect 51224 15892 51230 15904
rect 51920 15892 51948 15932
rect 52362 15892 52368 15904
rect 51224 15864 51948 15892
rect 52323 15864 52368 15892
rect 51224 15852 51230 15864
rect 52362 15852 52368 15864
rect 52420 15852 52426 15904
rect 53742 15852 53748 15904
rect 53800 15892 53806 15904
rect 58618 15892 58624 15904
rect 53800 15864 58624 15892
rect 53800 15852 53806 15864
rect 58618 15852 58624 15864
rect 58676 15852 58682 15904
rect 1104 15802 58880 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 58880 15802
rect 1104 15728 58880 15750
rect 13078 15648 13084 15700
rect 13136 15688 13142 15700
rect 13173 15691 13231 15697
rect 13173 15688 13185 15691
rect 13136 15660 13185 15688
rect 13136 15648 13142 15660
rect 13173 15657 13185 15660
rect 13219 15657 13231 15691
rect 24854 15688 24860 15700
rect 13173 15651 13231 15657
rect 13464 15660 24860 15688
rect 13354 15552 13360 15564
rect 13315 15524 13360 15552
rect 13354 15512 13360 15524
rect 13412 15512 13418 15564
rect 13464 15561 13492 15660
rect 24854 15648 24860 15660
rect 24912 15648 24918 15700
rect 25133 15691 25191 15697
rect 25133 15657 25145 15691
rect 25179 15688 25191 15691
rect 29454 15688 29460 15700
rect 25179 15660 29460 15688
rect 25179 15657 25191 15660
rect 25133 15651 25191 15657
rect 29454 15648 29460 15660
rect 29512 15648 29518 15700
rect 29730 15688 29736 15700
rect 29691 15660 29736 15688
rect 29730 15648 29736 15660
rect 29788 15648 29794 15700
rect 30024 15660 30420 15688
rect 16298 15580 16304 15632
rect 16356 15620 16362 15632
rect 19429 15623 19487 15629
rect 19429 15620 19441 15623
rect 16356 15592 19441 15620
rect 16356 15580 16362 15592
rect 19429 15589 19441 15592
rect 19475 15589 19487 15623
rect 19429 15583 19487 15589
rect 19981 15623 20039 15629
rect 19981 15589 19993 15623
rect 20027 15620 20039 15623
rect 20254 15620 20260 15632
rect 20027 15592 20260 15620
rect 20027 15589 20039 15592
rect 19981 15583 20039 15589
rect 13449 15555 13507 15561
rect 13449 15521 13461 15555
rect 13495 15521 13507 15555
rect 13449 15515 13507 15521
rect 13541 15555 13599 15561
rect 13541 15521 13553 15555
rect 13587 15552 13599 15555
rect 13722 15552 13728 15564
rect 13587 15524 13728 15552
rect 13587 15521 13599 15524
rect 13541 15515 13599 15521
rect 9858 15484 9864 15496
rect 9819 15456 9864 15484
rect 9858 15444 9864 15456
rect 9916 15444 9922 15496
rect 11606 15444 11612 15496
rect 11664 15484 11670 15496
rect 13556 15484 13584 15515
rect 13722 15512 13728 15524
rect 13780 15512 13786 15564
rect 14274 15552 14280 15564
rect 14235 15524 14280 15552
rect 14274 15512 14280 15524
rect 14332 15512 14338 15564
rect 14642 15512 14648 15564
rect 14700 15552 14706 15564
rect 15562 15552 15568 15564
rect 14700 15524 15568 15552
rect 14700 15512 14706 15524
rect 15562 15512 15568 15524
rect 15620 15512 15626 15564
rect 15933 15555 15991 15561
rect 15933 15521 15945 15555
rect 15979 15552 15991 15555
rect 18046 15552 18052 15564
rect 15979 15524 18052 15552
rect 15979 15521 15991 15524
rect 15933 15515 15991 15521
rect 18046 15512 18052 15524
rect 18104 15512 18110 15564
rect 19444 15552 19472 15583
rect 20254 15580 20260 15592
rect 20312 15580 20318 15632
rect 21450 15580 21456 15632
rect 21508 15620 21514 15632
rect 23474 15620 23480 15632
rect 21508 15592 23480 15620
rect 21508 15580 21514 15592
rect 23474 15580 23480 15592
rect 23532 15580 23538 15632
rect 26237 15623 26295 15629
rect 26237 15589 26249 15623
rect 26283 15589 26295 15623
rect 26237 15583 26295 15589
rect 23566 15552 23572 15564
rect 19444 15524 23572 15552
rect 23566 15512 23572 15524
rect 23624 15512 23630 15564
rect 24596 15524 25728 15552
rect 11664 15456 13584 15484
rect 13633 15487 13691 15493
rect 11664 15444 11670 15456
rect 13633 15453 13645 15487
rect 13679 15453 13691 15487
rect 13633 15447 13691 15453
rect 14553 15487 14611 15493
rect 14553 15453 14565 15487
rect 14599 15484 14611 15487
rect 15194 15484 15200 15496
rect 14599 15456 15200 15484
rect 14599 15453 14611 15456
rect 14553 15447 14611 15453
rect 12710 15376 12716 15428
rect 12768 15416 12774 15428
rect 13648 15416 13676 15447
rect 15194 15444 15200 15456
rect 15252 15444 15258 15496
rect 16577 15487 16635 15493
rect 16577 15453 16589 15487
rect 16623 15453 16635 15487
rect 16577 15447 16635 15453
rect 12768 15388 13676 15416
rect 16592 15416 16620 15447
rect 16666 15444 16672 15496
rect 16724 15484 16730 15496
rect 16724 15456 19564 15484
rect 16724 15444 16730 15456
rect 19242 15416 19248 15428
rect 16592 15388 19248 15416
rect 12768 15376 12774 15388
rect 19242 15376 19248 15388
rect 19300 15376 19306 15428
rect 19536 15416 19564 15456
rect 19610 15444 19616 15496
rect 19668 15484 19674 15496
rect 19797 15487 19855 15493
rect 19668 15456 19713 15484
rect 19668 15444 19674 15456
rect 19797 15453 19809 15487
rect 19843 15484 19855 15487
rect 20162 15484 20168 15496
rect 19843 15456 20168 15484
rect 19843 15453 19855 15456
rect 19797 15447 19855 15453
rect 20162 15444 20168 15456
rect 20220 15444 20226 15496
rect 21082 15484 21088 15496
rect 21043 15456 21088 15484
rect 21082 15444 21088 15456
rect 21140 15444 21146 15496
rect 23385 15487 23443 15493
rect 23385 15484 23397 15487
rect 22066 15456 23397 15484
rect 22066 15416 22094 15456
rect 23385 15453 23397 15456
rect 23431 15484 23443 15487
rect 23845 15487 23903 15493
rect 23845 15484 23857 15487
rect 23431 15456 23857 15484
rect 23431 15453 23443 15456
rect 23385 15447 23443 15453
rect 23845 15453 23857 15456
rect 23891 15453 23903 15487
rect 23845 15447 23903 15453
rect 24486 15444 24492 15496
rect 24544 15484 24550 15496
rect 24596 15493 24624 15524
rect 24581 15487 24639 15493
rect 24581 15484 24593 15487
rect 24544 15456 24593 15484
rect 24544 15444 24550 15456
rect 24581 15453 24593 15456
rect 24627 15453 24639 15487
rect 24857 15487 24915 15493
rect 24857 15484 24869 15487
rect 24581 15447 24639 15453
rect 24688 15456 24869 15484
rect 19536 15388 22094 15416
rect 23198 15376 23204 15428
rect 23256 15416 23262 15428
rect 24688 15416 24716 15456
rect 24857 15453 24869 15456
rect 24903 15453 24915 15487
rect 24857 15447 24915 15453
rect 24946 15444 24952 15496
rect 25004 15493 25010 15496
rect 25700 15493 25728 15524
rect 25004 15484 25012 15493
rect 25685 15487 25743 15493
rect 25004 15456 25268 15484
rect 25004 15447 25012 15456
rect 25004 15444 25010 15447
rect 23256 15388 24716 15416
rect 23256 15376 23262 15388
rect 24762 15376 24768 15428
rect 24820 15416 24826 15428
rect 24820 15388 24865 15416
rect 24820 15376 24826 15388
rect 10226 15308 10232 15360
rect 10284 15348 10290 15360
rect 11057 15351 11115 15357
rect 11057 15348 11069 15351
rect 10284 15320 11069 15348
rect 10284 15308 10290 15320
rect 11057 15317 11069 15320
rect 11103 15317 11115 15351
rect 11057 15311 11115 15317
rect 11882 15308 11888 15360
rect 11940 15348 11946 15360
rect 17218 15348 17224 15360
rect 11940 15320 17224 15348
rect 11940 15308 11946 15320
rect 17218 15308 17224 15320
rect 17276 15348 17282 15360
rect 17957 15351 18015 15357
rect 17957 15348 17969 15351
rect 17276 15320 17969 15348
rect 17276 15308 17282 15320
rect 17957 15317 17969 15320
rect 18003 15317 18015 15351
rect 17957 15311 18015 15317
rect 18414 15308 18420 15360
rect 18472 15348 18478 15360
rect 19150 15348 19156 15360
rect 18472 15320 19156 15348
rect 18472 15308 18478 15320
rect 19150 15308 19156 15320
rect 19208 15348 19214 15360
rect 19705 15351 19763 15357
rect 19705 15348 19717 15351
rect 19208 15320 19717 15348
rect 19208 15308 19214 15320
rect 19705 15317 19717 15320
rect 19751 15317 19763 15351
rect 19705 15311 19763 15317
rect 20070 15308 20076 15360
rect 20128 15348 20134 15360
rect 22646 15348 22652 15360
rect 20128 15320 22652 15348
rect 20128 15308 20134 15320
rect 22646 15308 22652 15320
rect 22704 15348 22710 15360
rect 23382 15348 23388 15360
rect 22704 15320 23388 15348
rect 22704 15308 22710 15320
rect 23382 15308 23388 15320
rect 23440 15308 23446 15360
rect 23474 15308 23480 15360
rect 23532 15348 23538 15360
rect 23937 15351 23995 15357
rect 23937 15348 23949 15351
rect 23532 15320 23949 15348
rect 23532 15308 23538 15320
rect 23937 15317 23949 15320
rect 23983 15348 23995 15351
rect 25130 15348 25136 15360
rect 23983 15320 25136 15348
rect 23983 15317 23995 15320
rect 23937 15311 23995 15317
rect 25130 15308 25136 15320
rect 25188 15308 25194 15360
rect 25240 15348 25268 15456
rect 25685 15453 25697 15487
rect 25731 15453 25743 15487
rect 25685 15447 25743 15453
rect 26105 15487 26163 15493
rect 26105 15453 26117 15487
rect 26151 15453 26163 15487
rect 26252 15484 26280 15583
rect 28442 15580 28448 15632
rect 28500 15620 28506 15632
rect 30024 15620 30052 15660
rect 28500 15592 30052 15620
rect 30392 15620 30420 15660
rect 31662 15648 31668 15700
rect 31720 15688 31726 15700
rect 41322 15688 41328 15700
rect 31720 15660 41328 15688
rect 31720 15648 31726 15660
rect 41322 15648 41328 15660
rect 41380 15648 41386 15700
rect 41690 15688 41696 15700
rect 41651 15660 41696 15688
rect 41690 15648 41696 15660
rect 41748 15648 41754 15700
rect 42518 15648 42524 15700
rect 42576 15688 42582 15700
rect 47394 15688 47400 15700
rect 42576 15660 47400 15688
rect 42576 15648 42582 15660
rect 47394 15648 47400 15660
rect 47452 15648 47458 15700
rect 51534 15688 51540 15700
rect 51495 15660 51540 15688
rect 51534 15648 51540 15660
rect 51592 15648 51598 15700
rect 30392 15592 32352 15620
rect 28500 15580 28506 15592
rect 26326 15512 26332 15564
rect 26384 15552 26390 15564
rect 27338 15552 27344 15564
rect 26384 15524 27344 15552
rect 26384 15512 26390 15524
rect 27338 15512 27344 15524
rect 27396 15512 27402 15564
rect 28718 15512 28724 15564
rect 28776 15552 28782 15564
rect 28902 15552 28908 15564
rect 28776 15524 28908 15552
rect 28776 15512 28782 15524
rect 28902 15512 28908 15524
rect 28960 15552 28966 15564
rect 30285 15555 30343 15561
rect 30285 15552 30297 15555
rect 28960 15524 30297 15552
rect 28960 15512 28966 15524
rect 30285 15521 30297 15524
rect 30331 15521 30343 15555
rect 30285 15515 30343 15521
rect 31662 15484 31668 15496
rect 26252 15456 31668 15484
rect 26105 15447 26163 15453
rect 25314 15376 25320 15428
rect 25372 15416 25378 15428
rect 25869 15419 25927 15425
rect 25869 15416 25881 15419
rect 25372 15388 25881 15416
rect 25372 15376 25378 15388
rect 25869 15385 25881 15388
rect 25915 15385 25927 15419
rect 25869 15379 25927 15385
rect 25958 15376 25964 15428
rect 26016 15416 26022 15428
rect 26016 15388 26061 15416
rect 26016 15376 26022 15388
rect 26120 15348 26148 15447
rect 31662 15444 31668 15456
rect 31720 15444 31726 15496
rect 32122 15484 32128 15496
rect 32083 15456 32128 15484
rect 32122 15444 32128 15456
rect 32180 15444 32186 15496
rect 32324 15493 32352 15592
rect 46750 15580 46756 15632
rect 46808 15620 46814 15632
rect 58802 15620 58808 15632
rect 46808 15592 58808 15620
rect 46808 15580 46814 15592
rect 58802 15580 58808 15592
rect 58860 15580 58866 15632
rect 41414 15512 41420 15564
rect 41472 15552 41478 15564
rect 53926 15552 53932 15564
rect 41472 15524 51028 15552
rect 41472 15512 41478 15524
rect 32309 15487 32367 15493
rect 32309 15453 32321 15487
rect 32355 15484 32367 15487
rect 34146 15484 34152 15496
rect 32355 15456 34152 15484
rect 32355 15453 32367 15456
rect 32309 15447 32367 15453
rect 34146 15444 34152 15456
rect 34204 15444 34210 15496
rect 36354 15484 36360 15496
rect 36315 15456 36360 15484
rect 36354 15444 36360 15456
rect 36412 15444 36418 15496
rect 36446 15444 36452 15496
rect 36504 15484 36510 15496
rect 36613 15487 36671 15493
rect 36613 15484 36625 15487
rect 36504 15456 36625 15484
rect 36504 15444 36510 15456
rect 36613 15453 36625 15456
rect 36659 15453 36671 15487
rect 41046 15484 41052 15496
rect 41007 15456 41052 15484
rect 36613 15447 36671 15453
rect 41046 15444 41052 15456
rect 41104 15444 41110 15496
rect 41142 15487 41200 15493
rect 41142 15453 41154 15487
rect 41188 15453 41200 15487
rect 41142 15447 41200 15453
rect 27608 15419 27666 15425
rect 27608 15385 27620 15419
rect 27654 15416 27666 15419
rect 29086 15416 29092 15428
rect 27654 15388 29092 15416
rect 27654 15385 27666 15388
rect 27608 15379 27666 15385
rect 29086 15376 29092 15388
rect 29144 15376 29150 15428
rect 29270 15376 29276 15428
rect 29328 15416 29334 15428
rect 29730 15416 29736 15428
rect 29328 15388 29736 15416
rect 29328 15376 29334 15388
rect 29730 15376 29736 15388
rect 29788 15376 29794 15428
rect 30006 15376 30012 15428
rect 30064 15416 30070 15428
rect 30193 15419 30251 15425
rect 30193 15416 30205 15419
rect 30064 15388 30205 15416
rect 30064 15376 30070 15388
rect 30193 15385 30205 15388
rect 30239 15385 30251 15419
rect 31110 15416 31116 15428
rect 30193 15379 30251 15385
rect 30300 15388 31116 15416
rect 27522 15348 27528 15360
rect 25240 15320 27528 15348
rect 27522 15308 27528 15320
rect 27580 15308 27586 15360
rect 28258 15308 28264 15360
rect 28316 15348 28322 15360
rect 28721 15351 28779 15357
rect 28721 15348 28733 15351
rect 28316 15320 28733 15348
rect 28316 15308 28322 15320
rect 28721 15317 28733 15320
rect 28767 15317 28779 15351
rect 28721 15311 28779 15317
rect 30101 15351 30159 15357
rect 30101 15317 30113 15351
rect 30147 15348 30159 15351
rect 30300 15348 30328 15388
rect 31110 15376 31116 15388
rect 31168 15376 31174 15428
rect 34330 15416 34336 15428
rect 31864 15388 34336 15416
rect 30147 15320 30328 15348
rect 30147 15317 30159 15320
rect 30101 15311 30159 15317
rect 30466 15308 30472 15360
rect 30524 15348 30530 15360
rect 31864 15348 31892 15388
rect 34330 15376 34336 15388
rect 34388 15376 34394 15428
rect 40126 15376 40132 15428
rect 40184 15416 40190 15428
rect 41156 15416 41184 15447
rect 41230 15444 41236 15496
rect 41288 15484 41294 15496
rect 41325 15487 41383 15493
rect 41325 15484 41337 15487
rect 41288 15456 41337 15484
rect 41288 15444 41294 15456
rect 41325 15453 41337 15456
rect 41371 15453 41383 15487
rect 41325 15447 41383 15453
rect 41555 15487 41613 15493
rect 41555 15453 41567 15487
rect 41601 15484 41613 15487
rect 42426 15484 42432 15496
rect 41601 15456 42432 15484
rect 41601 15453 41613 15456
rect 41555 15447 41613 15453
rect 40184 15388 41184 15416
rect 41417 15419 41475 15425
rect 40184 15376 40190 15388
rect 41417 15385 41429 15419
rect 41463 15416 41475 15419
rect 41782 15416 41788 15428
rect 41463 15388 41788 15416
rect 41463 15385 41475 15388
rect 41417 15379 41475 15385
rect 41782 15376 41788 15388
rect 41840 15376 41846 15428
rect 30524 15320 31892 15348
rect 30524 15308 30530 15320
rect 36722 15308 36728 15360
rect 36780 15348 36786 15360
rect 37737 15351 37795 15357
rect 37737 15348 37749 15351
rect 36780 15320 37749 15348
rect 36780 15308 36786 15320
rect 37737 15317 37749 15320
rect 37783 15317 37795 15351
rect 37737 15311 37795 15317
rect 40586 15308 40592 15360
rect 40644 15348 40650 15360
rect 41892 15348 41920 15456
rect 42426 15444 42432 15456
rect 42484 15444 42490 15496
rect 44174 15444 44180 15496
rect 44232 15484 44238 15496
rect 51000 15493 51028 15524
rect 51368 15524 53932 15552
rect 46845 15487 46903 15493
rect 46845 15484 46857 15487
rect 44232 15456 46857 15484
rect 44232 15444 44238 15456
rect 46845 15453 46857 15456
rect 46891 15453 46903 15487
rect 46845 15447 46903 15453
rect 50985 15487 51043 15493
rect 50985 15453 50997 15487
rect 51031 15453 51043 15487
rect 51166 15484 51172 15496
rect 51127 15456 51172 15484
rect 50985 15447 51043 15453
rect 51166 15444 51172 15456
rect 51224 15444 51230 15496
rect 51368 15493 51396 15524
rect 53926 15512 53932 15524
rect 53984 15512 53990 15564
rect 51353 15487 51411 15493
rect 51353 15453 51365 15487
rect 51399 15453 51411 15487
rect 51353 15447 51411 15453
rect 52362 15444 52368 15496
rect 52420 15484 52426 15496
rect 57885 15487 57943 15493
rect 57885 15484 57897 15487
rect 52420 15456 57897 15484
rect 52420 15444 52426 15456
rect 57885 15453 57897 15456
rect 57931 15453 57943 15487
rect 57885 15447 57943 15453
rect 51261 15419 51319 15425
rect 51261 15385 51273 15419
rect 51307 15416 51319 15419
rect 52380 15416 52408 15444
rect 58158 15416 58164 15428
rect 51307 15388 52408 15416
rect 58119 15388 58164 15416
rect 51307 15385 51319 15388
rect 51261 15379 51319 15385
rect 58158 15376 58164 15388
rect 58216 15376 58222 15428
rect 48130 15348 48136 15360
rect 40644 15320 41920 15348
rect 48091 15320 48136 15348
rect 40644 15308 40650 15320
rect 48130 15308 48136 15320
rect 48188 15308 48194 15360
rect 1104 15258 58880 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 58880 15258
rect 1104 15184 58880 15206
rect 12894 15104 12900 15156
rect 12952 15144 12958 15156
rect 13449 15147 13507 15153
rect 13449 15144 13461 15147
rect 12952 15116 13461 15144
rect 12952 15104 12958 15116
rect 13449 15113 13461 15116
rect 13495 15113 13507 15147
rect 13449 15107 13507 15113
rect 15749 15147 15807 15153
rect 15749 15113 15761 15147
rect 15795 15144 15807 15147
rect 15795 15116 18092 15144
rect 15795 15113 15807 15116
rect 15749 15107 15807 15113
rect 14550 15076 14556 15088
rect 2746 15048 14556 15076
rect 1581 15011 1639 15017
rect 1581 14977 1593 15011
rect 1627 15008 1639 15011
rect 2746 15008 2774 15048
rect 14550 15036 14556 15048
rect 14608 15036 14614 15088
rect 14734 15036 14740 15088
rect 14792 15076 14798 15088
rect 15838 15076 15844 15088
rect 14792 15048 15844 15076
rect 14792 15036 14798 15048
rect 15838 15036 15844 15048
rect 15896 15036 15902 15088
rect 16390 15036 16396 15088
rect 16448 15076 16454 15088
rect 17120 15079 17178 15085
rect 16448 15048 16988 15076
rect 16448 15036 16454 15048
rect 1627 14980 2774 15008
rect 8849 15011 8907 15017
rect 1627 14977 1639 14980
rect 1581 14971 1639 14977
rect 8849 14977 8861 15011
rect 8895 15008 8907 15011
rect 9766 15008 9772 15020
rect 8895 14980 9772 15008
rect 8895 14977 8907 14980
rect 8849 14971 8907 14977
rect 9766 14968 9772 14980
rect 9824 14968 9830 15020
rect 12250 15008 12256 15020
rect 12211 14980 12256 15008
rect 12250 14968 12256 14980
rect 12308 14968 12314 15020
rect 12618 14968 12624 15020
rect 12676 15008 12682 15020
rect 16022 15011 16028 15020
rect 15948 15008 16028 15011
rect 12676 14980 16028 15008
rect 12676 14968 12682 14980
rect 16022 14968 16028 14980
rect 16080 14968 16086 15020
rect 16117 15011 16175 15017
rect 16117 14977 16129 15011
rect 16163 14977 16175 15011
rect 16117 14971 16175 14977
rect 16209 15011 16267 15017
rect 16209 14977 16221 15011
rect 16255 15008 16267 15011
rect 16666 15008 16672 15020
rect 16255 14980 16672 15008
rect 16255 14977 16267 14980
rect 16209 14971 16267 14977
rect 1762 14940 1768 14952
rect 1723 14912 1768 14940
rect 1762 14900 1768 14912
rect 1820 14900 1826 14952
rect 15930 14900 15936 14952
rect 15988 14940 15994 14952
rect 16132 14940 16160 14971
rect 16666 14968 16672 14980
rect 16724 14968 16730 15020
rect 16850 15008 16856 15020
rect 16811 14980 16856 15008
rect 16850 14968 16856 14980
rect 16908 14968 16914 15020
rect 16960 15008 16988 15048
rect 17120 15045 17132 15079
rect 17166 15076 17178 15079
rect 17954 15076 17960 15088
rect 17166 15048 17960 15076
rect 17166 15045 17178 15048
rect 17120 15039 17178 15045
rect 17954 15036 17960 15048
rect 18012 15036 18018 15088
rect 18064 15008 18092 15116
rect 18138 15104 18144 15156
rect 18196 15144 18202 15156
rect 20165 15147 20223 15153
rect 20165 15144 20177 15147
rect 18196 15116 20177 15144
rect 18196 15104 18202 15116
rect 20165 15113 20177 15116
rect 20211 15113 20223 15147
rect 20165 15107 20223 15113
rect 22002 15104 22008 15156
rect 22060 15144 22066 15156
rect 22060 15116 24808 15144
rect 22060 15104 22066 15116
rect 18322 15036 18328 15088
rect 18380 15076 18386 15088
rect 20070 15076 20076 15088
rect 18380 15048 20076 15076
rect 18380 15036 18386 15048
rect 20070 15036 20076 15048
rect 20128 15036 20134 15088
rect 24780 15076 24808 15116
rect 25498 15104 25504 15156
rect 25556 15144 25562 15156
rect 26050 15144 26056 15156
rect 25556 15116 26056 15144
rect 25556 15104 25562 15116
rect 26050 15104 26056 15116
rect 26108 15144 26114 15156
rect 28258 15144 28264 15156
rect 26108 15116 28120 15144
rect 26108 15104 26114 15116
rect 26326 15076 26332 15088
rect 24780 15048 26332 15076
rect 24780 15020 24808 15048
rect 26326 15036 26332 15048
rect 26384 15036 26390 15088
rect 27522 15036 27528 15088
rect 27580 15076 27586 15088
rect 28092 15085 28120 15116
rect 28184 15116 28264 15144
rect 28184 15085 28212 15116
rect 28258 15104 28264 15116
rect 28316 15104 28322 15156
rect 28902 15104 28908 15156
rect 28960 15144 28966 15156
rect 29822 15144 29828 15156
rect 28960 15116 29828 15144
rect 28960 15104 28966 15116
rect 29822 15104 29828 15116
rect 29880 15144 29886 15156
rect 29880 15116 30420 15144
rect 29880 15104 29886 15116
rect 28077 15079 28135 15085
rect 27580 15048 28028 15076
rect 27580 15036 27586 15048
rect 18969 15011 19027 15017
rect 18969 15008 18981 15011
rect 16960 14980 18000 15008
rect 18064 14980 18981 15008
rect 16758 14940 16764 14952
rect 15988 14912 16033 14940
rect 16132 14912 16764 14940
rect 15988 14900 15994 14912
rect 16758 14900 16764 14912
rect 16816 14900 16822 14952
rect 17972 14940 18000 14980
rect 18969 14977 18981 14980
rect 19015 14977 19027 15011
rect 22005 15011 22063 15017
rect 22005 15008 22017 15011
rect 18969 14971 19027 14977
rect 19076 14980 22017 15008
rect 19076 14940 19104 14980
rect 22005 14977 22017 14980
rect 22051 15008 22063 15011
rect 24302 15008 24308 15020
rect 22051 14980 24308 15008
rect 22051 14977 22063 14980
rect 22005 14971 22063 14977
rect 24302 14968 24308 14980
rect 24360 14968 24366 15020
rect 24762 15008 24768 15020
rect 24675 14980 24768 15008
rect 24762 14968 24768 14980
rect 24820 14968 24826 15020
rect 25032 15011 25090 15017
rect 25032 14977 25044 15011
rect 25078 15008 25090 15011
rect 27614 15008 27620 15020
rect 25078 14980 27620 15008
rect 25078 14977 25090 14980
rect 25032 14971 25090 14977
rect 27614 14968 27620 14980
rect 27672 14968 27678 15020
rect 27890 15008 27896 15020
rect 27851 14980 27896 15008
rect 27890 14968 27896 14980
rect 27948 14968 27954 15020
rect 28000 15008 28028 15048
rect 28077 15045 28089 15079
rect 28123 15045 28135 15079
rect 28077 15039 28135 15045
rect 28169 15079 28227 15085
rect 28169 15045 28181 15079
rect 28215 15045 28227 15079
rect 28169 15039 28227 15045
rect 29270 15036 29276 15088
rect 29328 15076 29334 15088
rect 30392 15076 30420 15116
rect 30466 15104 30472 15156
rect 30524 15144 30530 15156
rect 32582 15144 32588 15156
rect 30524 15116 32588 15144
rect 30524 15104 30530 15116
rect 32582 15104 32588 15116
rect 32640 15104 32646 15156
rect 32674 15104 32680 15156
rect 32732 15144 32738 15156
rect 33873 15147 33931 15153
rect 33873 15144 33885 15147
rect 32732 15116 33885 15144
rect 32732 15104 32738 15116
rect 33873 15113 33885 15116
rect 33919 15144 33931 15147
rect 38657 15147 38715 15153
rect 33919 15116 36492 15144
rect 33919 15113 33931 15116
rect 33873 15107 33931 15113
rect 31938 15076 31944 15088
rect 29328 15048 30328 15076
rect 30392 15048 31944 15076
rect 29328 15036 29334 15048
rect 28266 15011 28324 15017
rect 28266 15008 28278 15011
rect 28000 14980 28278 15008
rect 28266 14977 28278 14980
rect 28312 14977 28324 15011
rect 28266 14971 28324 14977
rect 28626 14968 28632 15020
rect 28684 15008 28690 15020
rect 29181 15011 29239 15017
rect 29181 15008 29193 15011
rect 28684 14980 29193 15008
rect 28684 14968 28690 14980
rect 29181 14977 29193 14980
rect 29227 15008 29239 15011
rect 29822 15008 29828 15020
rect 29227 14980 29828 15008
rect 29227 14977 29239 14980
rect 29181 14971 29239 14977
rect 29822 14968 29828 14980
rect 29880 14968 29886 15020
rect 29917 15011 29975 15017
rect 29917 14977 29929 15011
rect 29963 15008 29975 15011
rect 30098 15008 30104 15020
rect 29963 14980 30104 15008
rect 29963 14977 29975 14980
rect 29917 14971 29975 14977
rect 17972 14912 19104 14940
rect 19242 14900 19248 14952
rect 19300 14940 19306 14952
rect 23109 14943 23167 14949
rect 23109 14940 23121 14943
rect 19300 14912 23121 14940
rect 19300 14900 19306 14912
rect 23109 14909 23121 14912
rect 23155 14909 23167 14943
rect 23109 14903 23167 14909
rect 25866 14900 25872 14952
rect 25924 14940 25930 14952
rect 27706 14940 27712 14952
rect 25924 14912 27712 14940
rect 25924 14900 25930 14912
rect 27706 14900 27712 14912
rect 27764 14900 27770 14952
rect 27982 14900 27988 14952
rect 28040 14940 28046 14952
rect 29932 14940 29960 14971
rect 30098 14968 30104 14980
rect 30156 14968 30162 15020
rect 28040 14912 29960 14940
rect 28040 14900 28046 14912
rect 30006 14900 30012 14952
rect 30064 14940 30070 14952
rect 30193 14943 30251 14949
rect 30193 14940 30205 14943
rect 30064 14912 30205 14940
rect 30064 14900 30070 14912
rect 30193 14909 30205 14912
rect 30239 14909 30251 14943
rect 30300 14940 30328 15048
rect 31938 15036 31944 15048
rect 31996 15036 32002 15088
rect 36354 15076 36360 15088
rect 34440 15048 36360 15076
rect 32030 14968 32036 15020
rect 32088 15008 32094 15020
rect 34440 15017 34468 15048
rect 36354 15036 36360 15048
rect 36412 15036 36418 15088
rect 36464 15076 36492 15116
rect 38657 15113 38669 15147
rect 38703 15144 38715 15147
rect 38930 15144 38936 15156
rect 38703 15116 38936 15144
rect 38703 15113 38715 15116
rect 38657 15107 38715 15113
rect 38930 15104 38936 15116
rect 38988 15104 38994 15156
rect 57698 15076 57704 15088
rect 36464 15048 57704 15076
rect 57698 15036 57704 15048
rect 57756 15036 57762 15088
rect 34698 15017 34704 15020
rect 32585 15011 32643 15017
rect 32585 15008 32597 15011
rect 32088 14980 32597 15008
rect 32088 14968 32094 14980
rect 32585 14977 32597 14980
rect 32631 14977 32643 15011
rect 32585 14971 32643 14977
rect 34425 15011 34483 15017
rect 34425 14977 34437 15011
rect 34471 14977 34483 15011
rect 34425 14971 34483 14977
rect 34692 14971 34704 15017
rect 34756 15008 34762 15020
rect 38654 15011 38712 15017
rect 34756 14980 34792 15008
rect 34698 14968 34704 14971
rect 34756 14968 34762 14980
rect 38654 14977 38666 15011
rect 38700 15008 38712 15011
rect 40310 15008 40316 15020
rect 38700 14980 40316 15008
rect 38700 14977 38712 14980
rect 38654 14971 38712 14977
rect 40310 14968 40316 14980
rect 40368 14968 40374 15020
rect 42889 15011 42947 15017
rect 42889 14977 42901 15011
rect 42935 15008 42947 15011
rect 43530 15008 43536 15020
rect 42935 14980 43536 15008
rect 42935 14977 42947 14980
rect 42889 14971 42947 14977
rect 43530 14968 43536 14980
rect 43588 14968 43594 15020
rect 31754 14940 31760 14952
rect 30300 14912 31760 14940
rect 30193 14903 30251 14909
rect 31754 14900 31760 14912
rect 31812 14900 31818 14952
rect 32309 14943 32367 14949
rect 32309 14909 32321 14943
rect 32355 14940 32367 14943
rect 33226 14940 33232 14952
rect 32355 14912 33232 14940
rect 32355 14909 32367 14912
rect 32309 14903 32367 14909
rect 33226 14900 33232 14912
rect 33284 14900 33290 14952
rect 38746 14900 38752 14952
rect 38804 14940 38810 14952
rect 39117 14943 39175 14949
rect 39117 14940 39129 14943
rect 38804 14912 39129 14940
rect 38804 14900 38810 14912
rect 39117 14909 39129 14912
rect 39163 14909 39175 14943
rect 39117 14903 39175 14909
rect 41138 14900 41144 14952
rect 41196 14940 41202 14952
rect 43073 14943 43131 14949
rect 43073 14940 43085 14943
rect 41196 14912 43085 14940
rect 41196 14900 41202 14912
rect 43073 14909 43085 14912
rect 43119 14940 43131 14943
rect 43162 14940 43168 14952
rect 43119 14912 43168 14940
rect 43119 14909 43131 14912
rect 43073 14903 43131 14909
rect 43162 14900 43168 14912
rect 43220 14900 43226 14952
rect 44358 14900 44364 14952
rect 44416 14940 44422 14952
rect 54846 14940 54852 14952
rect 44416 14912 54852 14940
rect 44416 14900 44422 14912
rect 54846 14900 54852 14912
rect 54904 14900 54910 14952
rect 1578 14832 1584 14884
rect 1636 14872 1642 14884
rect 15654 14872 15660 14884
rect 1636 14844 15660 14872
rect 1636 14832 1642 14844
rect 15654 14832 15660 14844
rect 15712 14832 15718 14884
rect 18233 14875 18291 14881
rect 18233 14841 18245 14875
rect 18279 14872 18291 14875
rect 19426 14872 19432 14884
rect 18279 14844 19432 14872
rect 18279 14841 18291 14844
rect 18233 14835 18291 14841
rect 19426 14832 19432 14844
rect 19484 14832 19490 14884
rect 28445 14875 28503 14881
rect 28445 14841 28457 14875
rect 28491 14872 28503 14875
rect 31018 14872 31024 14884
rect 28491 14844 31024 14872
rect 28491 14841 28503 14844
rect 28445 14835 28503 14841
rect 31018 14832 31024 14844
rect 31076 14832 31082 14884
rect 33502 14832 33508 14884
rect 33560 14872 33566 14884
rect 33560 14844 34468 14872
rect 33560 14832 33566 14844
rect 9674 14764 9680 14816
rect 9732 14804 9738 14816
rect 10045 14807 10103 14813
rect 10045 14804 10057 14807
rect 9732 14776 10057 14804
rect 9732 14764 9738 14776
rect 10045 14773 10057 14776
rect 10091 14773 10103 14807
rect 10045 14767 10103 14773
rect 15930 14764 15936 14816
rect 15988 14804 15994 14816
rect 18414 14804 18420 14816
rect 15988 14776 18420 14804
rect 15988 14764 15994 14776
rect 18414 14764 18420 14776
rect 18472 14764 18478 14816
rect 19518 14764 19524 14816
rect 19576 14804 19582 14816
rect 20622 14804 20628 14816
rect 19576 14776 20628 14804
rect 19576 14764 19582 14776
rect 20622 14764 20628 14776
rect 20680 14764 20686 14816
rect 24026 14764 24032 14816
rect 24084 14804 24090 14816
rect 24946 14804 24952 14816
rect 24084 14776 24952 14804
rect 24084 14764 24090 14776
rect 24946 14764 24952 14776
rect 25004 14764 25010 14816
rect 25406 14764 25412 14816
rect 25464 14804 25470 14816
rect 25958 14804 25964 14816
rect 25464 14776 25964 14804
rect 25464 14764 25470 14776
rect 25958 14764 25964 14776
rect 26016 14804 26022 14816
rect 26145 14807 26203 14813
rect 26145 14804 26157 14807
rect 26016 14776 26157 14804
rect 26016 14764 26022 14776
rect 26145 14773 26157 14776
rect 26191 14773 26203 14807
rect 26145 14767 26203 14773
rect 26326 14764 26332 14816
rect 26384 14804 26390 14816
rect 28902 14804 28908 14816
rect 26384 14776 28908 14804
rect 26384 14764 26390 14776
rect 28902 14764 28908 14776
rect 28960 14764 28966 14816
rect 29086 14764 29092 14816
rect 29144 14804 29150 14816
rect 29273 14807 29331 14813
rect 29273 14804 29285 14807
rect 29144 14776 29285 14804
rect 29144 14764 29150 14776
rect 29273 14773 29285 14776
rect 29319 14804 29331 14807
rect 29638 14804 29644 14816
rect 29319 14776 29644 14804
rect 29319 14773 29331 14776
rect 29273 14767 29331 14773
rect 29638 14764 29644 14776
rect 29696 14764 29702 14816
rect 32582 14764 32588 14816
rect 32640 14804 32646 14816
rect 34330 14804 34336 14816
rect 32640 14776 34336 14804
rect 32640 14764 32646 14776
rect 34330 14764 34336 14776
rect 34388 14764 34394 14816
rect 34440 14804 34468 14844
rect 35360 14844 39160 14872
rect 35360 14804 35388 14844
rect 34440 14776 35388 14804
rect 35805 14807 35863 14813
rect 35805 14773 35817 14807
rect 35851 14804 35863 14807
rect 35894 14804 35900 14816
rect 35851 14776 35900 14804
rect 35851 14773 35863 14776
rect 35805 14767 35863 14773
rect 35894 14764 35900 14776
rect 35952 14764 35958 14816
rect 38470 14804 38476 14816
rect 38431 14776 38476 14804
rect 38470 14764 38476 14776
rect 38528 14764 38534 14816
rect 38562 14764 38568 14816
rect 38620 14804 38626 14816
rect 39025 14807 39083 14813
rect 39025 14804 39037 14807
rect 38620 14776 39037 14804
rect 38620 14764 38626 14776
rect 39025 14773 39037 14776
rect 39071 14773 39083 14807
rect 39132 14804 39160 14844
rect 39482 14832 39488 14884
rect 39540 14872 39546 14884
rect 48314 14872 48320 14884
rect 39540 14844 48320 14872
rect 39540 14832 39546 14844
rect 48314 14832 48320 14844
rect 48372 14832 48378 14884
rect 41046 14804 41052 14816
rect 39132 14776 41052 14804
rect 39025 14767 39083 14773
rect 41046 14764 41052 14776
rect 41104 14764 41110 14816
rect 41598 14764 41604 14816
rect 41656 14804 41662 14816
rect 52454 14804 52460 14816
rect 41656 14776 52460 14804
rect 41656 14764 41662 14776
rect 52454 14764 52460 14776
rect 52512 14764 52518 14816
rect 1104 14714 58880 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 58880 14714
rect 1104 14640 58880 14662
rect 14550 14560 14556 14612
rect 14608 14600 14614 14612
rect 14608 14572 15240 14600
rect 14608 14560 14614 14572
rect 15212 14532 15240 14572
rect 19426 14560 19432 14612
rect 19484 14600 19490 14612
rect 22833 14603 22891 14609
rect 22833 14600 22845 14603
rect 19484 14572 22845 14600
rect 19484 14560 19490 14572
rect 22833 14569 22845 14572
rect 22879 14569 22891 14603
rect 27614 14600 27620 14612
rect 22833 14563 22891 14569
rect 24780 14572 27476 14600
rect 27575 14572 27620 14600
rect 19518 14532 19524 14544
rect 15212 14504 19524 14532
rect 19518 14492 19524 14504
rect 19576 14492 19582 14544
rect 20806 14492 20812 14544
rect 20864 14532 20870 14544
rect 24394 14532 24400 14544
rect 20864 14504 24400 14532
rect 20864 14492 20870 14504
rect 24394 14492 24400 14504
rect 24452 14492 24458 14544
rect 2406 14464 2412 14476
rect 1596 14436 2412 14464
rect 1596 14405 1624 14436
rect 2406 14424 2412 14436
rect 2464 14424 2470 14476
rect 8294 14424 8300 14476
rect 8352 14464 8358 14476
rect 9306 14464 9312 14476
rect 8352 14436 9312 14464
rect 8352 14424 8358 14436
rect 9306 14424 9312 14436
rect 9364 14424 9370 14476
rect 9585 14467 9643 14473
rect 9585 14433 9597 14467
rect 9631 14464 9643 14467
rect 10226 14464 10232 14476
rect 9631 14436 10232 14464
rect 9631 14433 9643 14436
rect 9585 14427 9643 14433
rect 10226 14424 10232 14436
rect 10284 14424 10290 14476
rect 14274 14464 14280 14476
rect 14235 14436 14280 14464
rect 14274 14424 14280 14436
rect 14332 14424 14338 14476
rect 15654 14424 15660 14476
rect 15712 14464 15718 14476
rect 19242 14464 19248 14476
rect 15712 14436 19248 14464
rect 15712 14424 15718 14436
rect 19242 14424 19248 14436
rect 19300 14424 19306 14476
rect 21818 14464 21824 14476
rect 21100 14436 21824 14464
rect 1581 14399 1639 14405
rect 1581 14365 1593 14399
rect 1627 14365 1639 14399
rect 1581 14359 1639 14365
rect 11146 14356 11152 14408
rect 11204 14396 11210 14408
rect 11425 14399 11483 14405
rect 11425 14396 11437 14399
rect 11204 14368 11437 14396
rect 11204 14356 11210 14368
rect 11425 14365 11437 14368
rect 11471 14365 11483 14399
rect 11425 14359 11483 14365
rect 14553 14399 14611 14405
rect 14553 14365 14565 14399
rect 14599 14396 14611 14399
rect 15378 14396 15384 14408
rect 14599 14368 15384 14396
rect 14599 14365 14611 14368
rect 14553 14359 14611 14365
rect 15378 14356 15384 14368
rect 15436 14356 15442 14408
rect 16577 14399 16635 14405
rect 16577 14365 16589 14399
rect 16623 14396 16635 14399
rect 18046 14396 18052 14408
rect 16623 14368 18052 14396
rect 16623 14365 16635 14368
rect 16577 14359 16635 14365
rect 18046 14356 18052 14368
rect 18104 14356 18110 14408
rect 19705 14399 19763 14405
rect 19705 14365 19717 14399
rect 19751 14396 19763 14399
rect 19794 14396 19800 14408
rect 19751 14368 19800 14396
rect 19751 14365 19763 14368
rect 19705 14359 19763 14365
rect 19794 14356 19800 14368
rect 19852 14396 19858 14408
rect 21100 14396 21128 14436
rect 21818 14424 21824 14436
rect 21876 14464 21882 14476
rect 22002 14464 22008 14476
rect 21876 14436 22008 14464
rect 21876 14424 21882 14436
rect 22002 14424 22008 14436
rect 22060 14424 22066 14476
rect 21634 14396 21640 14408
rect 19852 14368 21128 14396
rect 21595 14368 21640 14396
rect 19852 14356 19858 14368
rect 21634 14356 21640 14368
rect 21692 14396 21698 14408
rect 24780 14396 24808 14572
rect 25041 14535 25099 14541
rect 25041 14501 25053 14535
rect 25087 14532 25099 14535
rect 27448 14532 27476 14572
rect 27614 14560 27620 14572
rect 27672 14560 27678 14612
rect 27706 14560 27712 14612
rect 27764 14600 27770 14612
rect 29270 14600 29276 14612
rect 27764 14572 29276 14600
rect 27764 14560 27770 14572
rect 29270 14560 29276 14572
rect 29328 14560 29334 14612
rect 31110 14600 31116 14612
rect 29656 14572 31116 14600
rect 29656 14544 29684 14572
rect 31110 14560 31116 14572
rect 31168 14560 31174 14612
rect 31757 14603 31815 14609
rect 31757 14569 31769 14603
rect 31803 14600 31815 14603
rect 32030 14600 32036 14612
rect 31803 14572 32036 14600
rect 31803 14569 31815 14572
rect 31757 14563 31815 14569
rect 32030 14560 32036 14572
rect 32088 14560 32094 14612
rect 35250 14560 35256 14612
rect 35308 14600 35314 14612
rect 39393 14603 39451 14609
rect 35308 14572 38976 14600
rect 35308 14560 35314 14572
rect 29638 14532 29644 14544
rect 25087 14504 27292 14532
rect 27448 14504 29644 14532
rect 25087 14501 25099 14504
rect 25041 14495 25099 14501
rect 24854 14424 24860 14476
rect 24912 14464 24918 14476
rect 25685 14467 25743 14473
rect 25685 14464 25697 14467
rect 24912 14436 25697 14464
rect 24912 14424 24918 14436
rect 25685 14433 25697 14436
rect 25731 14464 25743 14467
rect 26142 14464 26148 14476
rect 25731 14436 26148 14464
rect 25731 14433 25743 14436
rect 25685 14427 25743 14433
rect 26142 14424 26148 14436
rect 26200 14424 26206 14476
rect 26418 14464 26424 14476
rect 26252 14436 26424 14464
rect 21692 14368 24808 14396
rect 25501 14399 25559 14405
rect 21692 14356 21698 14368
rect 25501 14365 25513 14399
rect 25547 14396 25559 14399
rect 25866 14396 25872 14408
rect 25547 14368 25872 14396
rect 25547 14365 25559 14368
rect 25501 14359 25559 14365
rect 1854 14328 1860 14340
rect 1815 14300 1860 14328
rect 1854 14288 1860 14300
rect 1912 14288 1918 14340
rect 10965 14331 11023 14337
rect 10965 14297 10977 14331
rect 11011 14328 11023 14331
rect 12434 14328 12440 14340
rect 11011 14300 12440 14328
rect 11011 14297 11023 14300
rect 10965 14291 11023 14297
rect 12434 14288 12440 14300
rect 12492 14288 12498 14340
rect 16758 14288 16764 14340
rect 16816 14328 16822 14340
rect 17586 14328 17592 14340
rect 16816 14300 17592 14328
rect 16816 14288 16822 14300
rect 17586 14288 17592 14300
rect 17644 14328 17650 14340
rect 19610 14328 19616 14340
rect 17644 14300 19616 14328
rect 17644 14288 17650 14300
rect 19610 14288 19616 14300
rect 19668 14288 19674 14340
rect 19972 14331 20030 14337
rect 19972 14297 19984 14331
rect 20018 14297 20030 14331
rect 19972 14291 20030 14297
rect 11974 14220 11980 14272
rect 12032 14260 12038 14272
rect 12621 14263 12679 14269
rect 12621 14260 12633 14263
rect 12032 14232 12633 14260
rect 12032 14220 12038 14232
rect 12621 14229 12633 14232
rect 12667 14229 12679 14263
rect 15654 14260 15660 14272
rect 15615 14232 15660 14260
rect 12621 14223 12679 14229
rect 15654 14220 15660 14232
rect 15712 14220 15718 14272
rect 17770 14260 17776 14272
rect 17731 14232 17776 14260
rect 17770 14220 17776 14232
rect 17828 14220 17834 14272
rect 19996 14260 20024 14291
rect 21450 14288 21456 14340
rect 21508 14328 21514 14340
rect 23842 14328 23848 14340
rect 21508 14300 23848 14328
rect 21508 14288 21514 14300
rect 23842 14288 23848 14300
rect 23900 14288 23906 14340
rect 24302 14288 24308 14340
rect 24360 14328 24366 14340
rect 25406 14328 25412 14340
rect 24360 14300 25412 14328
rect 24360 14288 24366 14300
rect 25406 14288 25412 14300
rect 25464 14288 25470 14340
rect 20898 14260 20904 14272
rect 19996 14232 20904 14260
rect 20898 14220 20904 14232
rect 20956 14220 20962 14272
rect 21082 14260 21088 14272
rect 21043 14232 21088 14260
rect 21082 14220 21088 14232
rect 21140 14220 21146 14272
rect 22922 14220 22928 14272
rect 22980 14260 22986 14272
rect 25516 14260 25544 14359
rect 25866 14356 25872 14368
rect 25924 14356 25930 14408
rect 26252 14405 26280 14436
rect 26418 14424 26424 14436
rect 26476 14424 26482 14476
rect 27154 14464 27160 14476
rect 26528 14436 27160 14464
rect 26528 14405 26556 14436
rect 27154 14424 27160 14436
rect 27212 14424 27218 14476
rect 27264 14464 27292 14504
rect 29638 14492 29644 14504
rect 29696 14492 29702 14544
rect 30742 14492 30748 14544
rect 30800 14532 30806 14544
rect 35986 14532 35992 14544
rect 30800 14504 33548 14532
rect 30800 14492 30806 14504
rect 28813 14467 28871 14473
rect 27264 14436 27384 14464
rect 26237 14399 26295 14405
rect 26237 14365 26249 14399
rect 26283 14365 26295 14399
rect 26237 14359 26295 14365
rect 26513 14399 26571 14405
rect 26513 14365 26525 14399
rect 26559 14365 26571 14399
rect 26513 14359 26571 14365
rect 26602 14356 26608 14408
rect 26660 14396 26666 14408
rect 27246 14396 27252 14408
rect 26660 14368 26753 14396
rect 27207 14368 27252 14396
rect 26660 14356 26666 14368
rect 27246 14356 27252 14368
rect 27304 14356 27310 14408
rect 27356 14396 27384 14436
rect 28813 14433 28825 14467
rect 28859 14464 28871 14467
rect 29086 14464 29092 14476
rect 28859 14436 29092 14464
rect 28859 14433 28871 14436
rect 28813 14427 28871 14433
rect 29086 14424 29092 14436
rect 29144 14424 29150 14476
rect 32769 14467 32827 14473
rect 32769 14464 32781 14467
rect 31772 14436 32352 14464
rect 27433 14399 27491 14405
rect 27433 14396 27445 14399
rect 27356 14368 27445 14396
rect 27433 14365 27445 14368
rect 27479 14365 27491 14399
rect 27433 14359 27491 14365
rect 28997 14399 29055 14405
rect 28997 14365 29009 14399
rect 29043 14396 29055 14399
rect 29270 14396 29276 14408
rect 29043 14368 29276 14396
rect 29043 14365 29055 14368
rect 28997 14359 29055 14365
rect 29270 14356 29276 14368
rect 29328 14356 29334 14408
rect 29730 14396 29736 14408
rect 29691 14368 29736 14396
rect 29730 14356 29736 14368
rect 29788 14356 29794 14408
rect 31772 14405 31800 14436
rect 31757 14399 31815 14405
rect 31757 14365 31769 14399
rect 31803 14365 31815 14399
rect 31757 14359 31815 14365
rect 31941 14399 31999 14405
rect 31941 14365 31953 14399
rect 31987 14365 31999 14399
rect 32324 14396 32352 14436
rect 32508 14436 32781 14464
rect 32508 14396 32536 14436
rect 32769 14433 32781 14436
rect 32815 14433 32827 14467
rect 33410 14464 33416 14476
rect 32769 14427 32827 14433
rect 32968 14436 33416 14464
rect 32674 14396 32680 14408
rect 32324 14368 32536 14396
rect 32635 14368 32680 14396
rect 31941 14359 31999 14365
rect 26326 14288 26332 14340
rect 26384 14328 26390 14340
rect 26421 14331 26479 14337
rect 26421 14328 26433 14331
rect 26384 14300 26433 14328
rect 26384 14288 26390 14300
rect 26421 14297 26433 14300
rect 26467 14297 26479 14331
rect 26620 14328 26648 14356
rect 27982 14328 27988 14340
rect 26620 14300 27988 14328
rect 26421 14291 26479 14297
rect 27982 14288 27988 14300
rect 28040 14288 28046 14340
rect 29181 14331 29239 14337
rect 29181 14297 29193 14331
rect 29227 14328 29239 14331
rect 29978 14331 30036 14337
rect 29978 14328 29990 14331
rect 29227 14300 29990 14328
rect 29227 14297 29239 14300
rect 29181 14291 29239 14297
rect 29978 14297 29990 14300
rect 30024 14297 30036 14331
rect 29978 14291 30036 14297
rect 30190 14288 30196 14340
rect 30248 14328 30254 14340
rect 31956 14328 31984 14359
rect 32674 14356 32680 14368
rect 32732 14356 32738 14408
rect 32968 14405 32996 14436
rect 33410 14424 33416 14436
rect 33468 14424 33474 14476
rect 32953 14399 33011 14405
rect 32953 14365 32965 14399
rect 32999 14365 33011 14399
rect 32953 14359 33011 14365
rect 33042 14356 33048 14408
rect 33100 14396 33106 14408
rect 33137 14399 33195 14405
rect 33137 14396 33149 14399
rect 33100 14368 33149 14396
rect 33100 14356 33106 14368
rect 33137 14365 33149 14368
rect 33183 14365 33195 14399
rect 33520 14396 33548 14504
rect 34256 14504 35992 14532
rect 34256 14405 34284 14504
rect 35986 14492 35992 14504
rect 36044 14492 36050 14544
rect 38948 14532 38976 14572
rect 39393 14569 39405 14603
rect 39439 14600 39451 14603
rect 39482 14600 39488 14612
rect 39439 14572 39488 14600
rect 39439 14569 39451 14572
rect 39393 14563 39451 14569
rect 39482 14560 39488 14572
rect 39540 14560 39546 14612
rect 40218 14600 40224 14612
rect 39592 14572 40224 14600
rect 39592 14532 39620 14572
rect 40218 14560 40224 14572
rect 40276 14560 40282 14612
rect 40310 14560 40316 14612
rect 40368 14600 40374 14612
rect 41417 14603 41475 14609
rect 41417 14600 41429 14603
rect 40368 14572 41429 14600
rect 40368 14560 40374 14572
rect 41417 14569 41429 14572
rect 41463 14600 41475 14603
rect 44358 14600 44364 14612
rect 41463 14572 44364 14600
rect 41463 14569 41475 14572
rect 41417 14563 41475 14569
rect 44358 14560 44364 14572
rect 44416 14560 44422 14612
rect 44542 14600 44548 14612
rect 44455 14572 44548 14600
rect 44542 14560 44548 14572
rect 44600 14600 44606 14612
rect 48133 14603 48191 14609
rect 44600 14572 47716 14600
rect 44600 14560 44606 14572
rect 38948 14504 39620 14532
rect 47688 14532 47716 14572
rect 48133 14569 48145 14603
rect 48179 14600 48191 14603
rect 48222 14600 48228 14612
rect 48179 14572 48228 14600
rect 48179 14569 48191 14572
rect 48133 14563 48191 14569
rect 48222 14560 48228 14572
rect 48280 14560 48286 14612
rect 48314 14560 48320 14612
rect 48372 14600 48378 14612
rect 56594 14600 56600 14612
rect 48372 14572 56600 14600
rect 48372 14560 48378 14572
rect 56594 14560 56600 14572
rect 56652 14560 56658 14612
rect 56778 14532 56784 14544
rect 47688 14504 56784 14532
rect 56778 14492 56784 14504
rect 56836 14492 56842 14544
rect 34606 14424 34612 14476
rect 34664 14464 34670 14476
rect 35066 14464 35072 14476
rect 34664 14436 35072 14464
rect 34664 14424 34670 14436
rect 35066 14424 35072 14436
rect 35124 14424 35130 14476
rect 35158 14424 35164 14476
rect 35216 14464 35222 14476
rect 35529 14467 35587 14473
rect 35529 14464 35541 14467
rect 35216 14436 35541 14464
rect 35216 14424 35222 14436
rect 35529 14433 35541 14436
rect 35575 14464 35587 14467
rect 35618 14464 35624 14476
rect 35575 14436 35624 14464
rect 35575 14433 35587 14436
rect 35529 14427 35587 14433
rect 35618 14424 35624 14436
rect 35676 14424 35682 14476
rect 37461 14467 37519 14473
rect 37461 14433 37473 14467
rect 37507 14464 37519 14467
rect 37507 14436 37872 14464
rect 37507 14433 37519 14436
rect 37461 14427 37519 14433
rect 33597 14399 33655 14405
rect 33597 14396 33609 14399
rect 33520 14368 33609 14396
rect 33137 14359 33195 14365
rect 33597 14365 33609 14368
rect 33643 14365 33655 14399
rect 33597 14359 33655 14365
rect 34241 14399 34299 14405
rect 34241 14365 34253 14399
rect 34287 14365 34299 14399
rect 37366 14396 37372 14408
rect 34241 14359 34299 14365
rect 34348 14368 35664 14396
rect 37327 14368 37372 14396
rect 34348 14328 34376 14368
rect 35345 14331 35403 14337
rect 35345 14328 35357 14331
rect 30248 14300 34376 14328
rect 34808 14300 35357 14328
rect 30248 14288 30254 14300
rect 22980 14232 25544 14260
rect 22980 14220 22986 14232
rect 25682 14220 25688 14272
rect 25740 14260 25746 14272
rect 26789 14263 26847 14269
rect 26789 14260 26801 14263
rect 25740 14232 26801 14260
rect 25740 14220 25746 14232
rect 26789 14229 26801 14232
rect 26835 14229 26847 14263
rect 26789 14223 26847 14229
rect 27154 14220 27160 14272
rect 27212 14260 27218 14272
rect 31662 14260 31668 14272
rect 27212 14232 31668 14260
rect 27212 14220 27218 14232
rect 31662 14220 31668 14232
rect 31720 14220 31726 14272
rect 31754 14220 31760 14272
rect 31812 14260 31818 14272
rect 33502 14260 33508 14272
rect 31812 14232 33508 14260
rect 31812 14220 31818 14232
rect 33502 14220 33508 14232
rect 33560 14220 33566 14272
rect 33594 14220 33600 14272
rect 33652 14260 33658 14272
rect 34808 14260 34836 14300
rect 35345 14297 35357 14300
rect 35391 14297 35403 14331
rect 35636 14328 35664 14368
rect 37366 14356 37372 14368
rect 37424 14356 37430 14408
rect 37553 14399 37611 14405
rect 37553 14365 37565 14399
rect 37599 14365 37611 14399
rect 37553 14359 37611 14365
rect 37568 14328 37596 14359
rect 35636 14300 37596 14328
rect 37844 14328 37872 14436
rect 41046 14424 41052 14476
rect 41104 14464 41110 14476
rect 41104 14436 46244 14464
rect 41104 14424 41110 14436
rect 38013 14399 38071 14405
rect 38013 14365 38025 14399
rect 38059 14396 38071 14399
rect 39942 14396 39948 14408
rect 38059 14368 39948 14396
rect 38059 14365 38071 14368
rect 38013 14359 38071 14365
rect 39942 14356 39948 14368
rect 40000 14396 40006 14408
rect 40037 14399 40095 14405
rect 40037 14396 40049 14399
rect 40000 14368 40049 14396
rect 40000 14356 40006 14368
rect 40037 14365 40049 14368
rect 40083 14396 40095 14399
rect 42981 14399 43039 14405
rect 42981 14396 42993 14399
rect 40083 14368 42993 14396
rect 40083 14365 40095 14368
rect 40037 14359 40095 14365
rect 42981 14365 42993 14368
rect 43027 14396 43039 14399
rect 43070 14396 43076 14408
rect 43027 14368 43076 14396
rect 43027 14365 43039 14368
rect 42981 14359 43039 14365
rect 43070 14356 43076 14368
rect 43128 14356 43134 14408
rect 43254 14396 43260 14408
rect 43215 14368 43260 14396
rect 43254 14356 43260 14368
rect 43312 14356 43318 14408
rect 38258 14331 38316 14337
rect 38258 14328 38270 14331
rect 37844 14300 38270 14328
rect 35345 14291 35403 14297
rect 33652 14232 34836 14260
rect 33652 14220 33658 14232
rect 34882 14220 34888 14272
rect 34940 14260 34946 14272
rect 34940 14232 34985 14260
rect 34940 14220 34946 14232
rect 35066 14220 35072 14272
rect 35124 14260 35130 14272
rect 35253 14263 35311 14269
rect 35253 14260 35265 14263
rect 35124 14232 35265 14260
rect 35124 14220 35130 14232
rect 35253 14229 35265 14232
rect 35299 14229 35311 14263
rect 35360 14260 35388 14291
rect 35894 14260 35900 14272
rect 35360 14232 35900 14260
rect 35253 14223 35311 14229
rect 35894 14220 35900 14232
rect 35952 14220 35958 14272
rect 37568 14260 37596 14300
rect 38258 14297 38270 14300
rect 38304 14297 38316 14331
rect 38258 14291 38316 14297
rect 39114 14288 39120 14340
rect 39172 14328 39178 14340
rect 40282 14331 40340 14337
rect 40282 14328 40294 14331
rect 39172 14300 40294 14328
rect 39172 14288 39178 14300
rect 40282 14297 40294 14300
rect 40328 14297 40340 14331
rect 40282 14291 40340 14297
rect 41782 14260 41788 14272
rect 37568 14232 41788 14260
rect 41782 14220 41788 14232
rect 41840 14220 41846 14272
rect 46216 14260 46244 14436
rect 46753 14399 46811 14405
rect 46753 14365 46765 14399
rect 46799 14396 46811 14399
rect 48130 14396 48136 14408
rect 46799 14368 48136 14396
rect 46799 14365 46811 14368
rect 46753 14359 46811 14365
rect 48130 14356 48136 14368
rect 48188 14356 48194 14408
rect 57974 14396 57980 14408
rect 57935 14368 57980 14396
rect 57974 14356 57980 14368
rect 58032 14356 58038 14408
rect 47020 14331 47078 14337
rect 47020 14297 47032 14331
rect 47066 14328 47078 14331
rect 47762 14328 47768 14340
rect 47066 14300 47768 14328
rect 47066 14297 47078 14300
rect 47020 14291 47078 14297
rect 47762 14288 47768 14300
rect 47820 14288 47826 14340
rect 58069 14263 58127 14269
rect 58069 14260 58081 14263
rect 46216 14232 58081 14260
rect 58069 14229 58081 14232
rect 58115 14229 58127 14263
rect 58069 14223 58127 14229
rect 1104 14170 58880 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 58880 14170
rect 1104 14096 58880 14118
rect 10042 14056 10048 14068
rect 10003 14028 10048 14056
rect 10042 14016 10048 14028
rect 10100 14016 10106 14068
rect 13081 14059 13139 14065
rect 13081 14025 13093 14059
rect 13127 14056 13139 14059
rect 18233 14059 18291 14065
rect 13127 14028 18184 14056
rect 13127 14025 13139 14028
rect 13081 14019 13139 14025
rect 14274 13988 14280 14000
rect 11716 13960 14280 13988
rect 1578 13920 1584 13932
rect 1539 13892 1584 13920
rect 1578 13880 1584 13892
rect 1636 13880 1642 13932
rect 8846 13920 8852 13932
rect 8807 13892 8852 13920
rect 8846 13880 8852 13892
rect 8904 13880 8910 13932
rect 9306 13880 9312 13932
rect 9364 13920 9370 13932
rect 11716 13929 11744 13960
rect 14274 13948 14280 13960
rect 14332 13948 14338 14000
rect 17120 13991 17178 13997
rect 17120 13957 17132 13991
rect 17166 13988 17178 13991
rect 17770 13988 17776 14000
rect 17166 13960 17776 13988
rect 17166 13957 17178 13960
rect 17120 13951 17178 13957
rect 17770 13948 17776 13960
rect 17828 13948 17834 14000
rect 18156 13988 18184 14028
rect 18233 14025 18245 14059
rect 18279 14056 18291 14059
rect 21082 14056 21088 14068
rect 18279 14028 21088 14056
rect 18279 14025 18291 14028
rect 18233 14019 18291 14025
rect 21082 14016 21088 14028
rect 21140 14056 21146 14068
rect 24213 14059 24271 14065
rect 24213 14056 24225 14059
rect 21140 14028 24225 14056
rect 21140 14016 21146 14028
rect 24213 14025 24225 14028
rect 24259 14025 24271 14059
rect 24213 14019 24271 14025
rect 24394 14016 24400 14068
rect 24452 14056 24458 14068
rect 25133 14059 25191 14065
rect 25133 14056 25145 14059
rect 24452 14028 25145 14056
rect 24452 14016 24458 14028
rect 25133 14025 25145 14028
rect 25179 14056 25191 14059
rect 26418 14056 26424 14068
rect 25179 14028 26424 14056
rect 25179 14025 25191 14028
rect 25133 14019 25191 14025
rect 26418 14016 26424 14028
rect 26476 14016 26482 14068
rect 27433 14059 27491 14065
rect 27433 14025 27445 14059
rect 27479 14056 27491 14059
rect 28074 14056 28080 14068
rect 27479 14028 28080 14056
rect 27479 14025 27491 14028
rect 27433 14019 27491 14025
rect 28074 14016 28080 14028
rect 28132 14016 28138 14068
rect 29270 14056 29276 14068
rect 29231 14028 29276 14056
rect 29270 14016 29276 14028
rect 29328 14016 29334 14068
rect 31754 14056 31760 14068
rect 29380 14028 31760 14056
rect 21634 13988 21640 14000
rect 18156 13960 21640 13988
rect 21634 13948 21640 13960
rect 21692 13948 21698 14000
rect 23014 13988 23020 14000
rect 22940 13960 23020 13988
rect 11974 13929 11980 13932
rect 11701 13923 11759 13929
rect 11701 13920 11713 13923
rect 9364 13892 11713 13920
rect 9364 13880 9370 13892
rect 11701 13889 11713 13892
rect 11747 13889 11759 13923
rect 11968 13920 11980 13929
rect 11935 13892 11980 13920
rect 11701 13883 11759 13889
rect 11968 13883 11980 13892
rect 11974 13880 11980 13883
rect 12032 13880 12038 13932
rect 13722 13920 13728 13932
rect 13683 13892 13728 13920
rect 13722 13880 13728 13892
rect 13780 13880 13786 13932
rect 16850 13920 16856 13932
rect 16811 13892 16856 13920
rect 16850 13880 16856 13892
rect 16908 13880 16914 13932
rect 19153 13923 19211 13929
rect 19153 13889 19165 13923
rect 19199 13920 19211 13923
rect 20714 13920 20720 13932
rect 19199 13892 20720 13920
rect 19199 13889 19211 13892
rect 19153 13883 19211 13889
rect 20714 13880 20720 13892
rect 20772 13880 20778 13932
rect 21450 13920 21456 13932
rect 21411 13892 21456 13920
rect 21450 13880 21456 13892
rect 21508 13880 21514 13932
rect 21818 13920 21824 13932
rect 21779 13892 21824 13920
rect 21818 13880 21824 13892
rect 21876 13880 21882 13932
rect 22088 13923 22146 13929
rect 22088 13889 22100 13923
rect 22134 13920 22146 13923
rect 22370 13920 22376 13932
rect 22134 13892 22376 13920
rect 22134 13889 22146 13892
rect 22088 13883 22146 13889
rect 22370 13880 22376 13892
rect 22428 13880 22434 13932
rect 1762 13852 1768 13864
rect 1723 13824 1768 13852
rect 1762 13812 1768 13824
rect 1820 13812 1826 13864
rect 15194 13852 15200 13864
rect 15155 13824 15200 13852
rect 15194 13812 15200 13824
rect 15252 13812 15258 13864
rect 18230 13812 18236 13864
rect 18288 13852 18294 13864
rect 20806 13852 20812 13864
rect 18288 13824 20812 13852
rect 18288 13812 18294 13824
rect 20806 13812 20812 13824
rect 20864 13812 20870 13864
rect 21818 13784 21824 13796
rect 2746 13756 10180 13784
rect 1578 13676 1584 13728
rect 1636 13716 1642 13728
rect 2746 13716 2774 13756
rect 1636 13688 2774 13716
rect 10152 13716 10180 13756
rect 17788 13756 21824 13784
rect 17788 13716 17816 13756
rect 21818 13744 21824 13756
rect 21876 13744 21882 13796
rect 10152 13688 17816 13716
rect 1636 13676 1642 13688
rect 17954 13676 17960 13728
rect 18012 13716 18018 13728
rect 19426 13716 19432 13728
rect 18012 13688 19432 13716
rect 18012 13676 18018 13688
rect 19426 13676 19432 13688
rect 19484 13676 19490 13728
rect 22186 13676 22192 13728
rect 22244 13716 22250 13728
rect 22940 13716 22968 13960
rect 23014 13948 23020 13960
rect 23072 13948 23078 14000
rect 23934 13948 23940 14000
rect 23992 13988 23998 14000
rect 29380 13988 29408 14028
rect 31754 14016 31760 14028
rect 31812 14016 31818 14068
rect 32122 14016 32128 14068
rect 32180 14056 32186 14068
rect 32401 14059 32459 14065
rect 32401 14056 32413 14059
rect 32180 14028 32413 14056
rect 32180 14016 32186 14028
rect 32401 14025 32413 14028
rect 32447 14056 32459 14059
rect 33042 14056 33048 14068
rect 32447 14028 33048 14056
rect 32447 14025 32459 14028
rect 32401 14019 32459 14025
rect 33042 14016 33048 14028
rect 33100 14016 33106 14068
rect 34514 14016 34520 14068
rect 34572 14056 34578 14068
rect 35618 14056 35624 14068
rect 34572 14028 35624 14056
rect 34572 14016 34578 14028
rect 35618 14016 35624 14028
rect 35676 14016 35682 14068
rect 37366 14016 37372 14068
rect 37424 14056 37430 14068
rect 37921 14059 37979 14065
rect 37921 14056 37933 14059
rect 37424 14028 37933 14056
rect 37424 14016 37430 14028
rect 37921 14025 37933 14028
rect 37967 14025 37979 14059
rect 37921 14019 37979 14025
rect 38105 14059 38163 14065
rect 38105 14025 38117 14059
rect 38151 14056 38163 14059
rect 38930 14056 38936 14068
rect 38151 14028 38936 14056
rect 38151 14025 38163 14028
rect 38105 14019 38163 14025
rect 32030 13988 32036 14000
rect 23992 13960 25544 13988
rect 23992 13948 23998 13960
rect 23566 13920 23572 13932
rect 23479 13892 23572 13920
rect 23566 13880 23572 13892
rect 23624 13920 23630 13932
rect 23624 13892 24164 13920
rect 23624 13880 23630 13892
rect 23014 13812 23020 13864
rect 23072 13852 23078 13864
rect 24136 13852 24164 13892
rect 24946 13880 24952 13932
rect 25004 13920 25010 13932
rect 25308 13923 25366 13929
rect 25308 13920 25320 13923
rect 25004 13892 25320 13920
rect 25004 13880 25010 13892
rect 25308 13889 25320 13892
rect 25354 13889 25366 13923
rect 25308 13883 25366 13889
rect 25409 13923 25467 13929
rect 25409 13889 25421 13923
rect 25455 13889 25467 13923
rect 25516 13926 25544 13960
rect 26068 13960 29408 13988
rect 31128 13960 32036 13988
rect 25593 13926 25651 13929
rect 25516 13923 25651 13926
rect 25516 13898 25605 13923
rect 25409 13883 25467 13889
rect 25593 13889 25605 13898
rect 25639 13889 25651 13923
rect 25593 13883 25651 13889
rect 24305 13855 24363 13861
rect 24305 13852 24317 13855
rect 23072 13824 23888 13852
rect 24136 13824 24317 13852
rect 23072 13812 23078 13824
rect 23198 13784 23204 13796
rect 23159 13756 23204 13784
rect 23198 13744 23204 13756
rect 23256 13744 23262 13796
rect 23860 13793 23888 13824
rect 24305 13821 24317 13824
rect 24351 13852 24363 13855
rect 24394 13852 24400 13864
rect 24351 13824 24400 13852
rect 24351 13821 24363 13824
rect 24305 13815 24363 13821
rect 24394 13812 24400 13824
rect 24452 13812 24458 13864
rect 24489 13855 24547 13861
rect 24489 13821 24501 13855
rect 24535 13852 24547 13855
rect 24854 13852 24860 13864
rect 24535 13824 24860 13852
rect 24535 13821 24547 13824
rect 24489 13815 24547 13821
rect 24854 13812 24860 13824
rect 24912 13812 24918 13864
rect 23845 13787 23903 13793
rect 23845 13753 23857 13787
rect 23891 13753 23903 13787
rect 25323 13784 25351 13883
rect 25424 13852 25452 13883
rect 25682 13880 25688 13932
rect 25740 13920 25746 13932
rect 25740 13892 25785 13920
rect 25740 13880 25746 13892
rect 26068 13852 26096 13960
rect 26145 13923 26203 13929
rect 26145 13889 26157 13923
rect 26191 13889 26203 13923
rect 26145 13883 26203 13889
rect 25424 13824 26096 13852
rect 25958 13784 25964 13796
rect 25323 13756 25964 13784
rect 23845 13747 23903 13753
rect 25958 13744 25964 13756
rect 26016 13744 26022 13796
rect 26160 13784 26188 13883
rect 26510 13880 26516 13932
rect 26568 13920 26574 13932
rect 27341 13923 27399 13929
rect 27341 13920 27353 13923
rect 26568 13892 27353 13920
rect 26568 13880 26574 13892
rect 27341 13889 27353 13892
rect 27387 13889 27399 13923
rect 27522 13920 27528 13932
rect 27483 13892 27528 13920
rect 27341 13883 27399 13889
rect 27522 13880 27528 13892
rect 27580 13880 27586 13932
rect 29638 13920 29644 13932
rect 29599 13892 29644 13920
rect 29638 13880 29644 13892
rect 29696 13880 29702 13932
rect 31128 13929 31156 13960
rect 32030 13948 32036 13960
rect 32088 13948 32094 14000
rect 33410 13948 33416 14000
rect 33468 13988 33474 14000
rect 38120 13988 38148 14019
rect 38930 14016 38936 14028
rect 38988 14016 38994 14068
rect 39114 14056 39120 14068
rect 39075 14028 39120 14056
rect 39114 14016 39120 14028
rect 39172 14016 39178 14068
rect 42794 14016 42800 14068
rect 42852 14056 42858 14068
rect 44082 14056 44088 14068
rect 42852 14028 44088 14056
rect 42852 14016 42858 14028
rect 44082 14016 44088 14028
rect 44140 14016 44146 14068
rect 39482 13988 39488 14000
rect 33468 13960 38148 13988
rect 38396 13960 39488 13988
rect 33468 13948 33474 13960
rect 31113 13923 31171 13929
rect 31113 13889 31125 13923
rect 31159 13889 31171 13923
rect 31113 13883 31171 13889
rect 31205 13923 31263 13929
rect 31205 13889 31217 13923
rect 31251 13920 31263 13923
rect 31294 13920 31300 13932
rect 31251 13892 31300 13920
rect 31251 13889 31263 13892
rect 31205 13883 31263 13889
rect 31294 13880 31300 13892
rect 31352 13880 31358 13932
rect 31478 13920 31484 13932
rect 31439 13892 31484 13920
rect 31478 13880 31484 13892
rect 31536 13880 31542 13932
rect 31665 13923 31723 13929
rect 31665 13889 31677 13923
rect 31711 13920 31723 13923
rect 31846 13920 31852 13932
rect 31711 13892 31852 13920
rect 31711 13889 31723 13892
rect 31665 13883 31723 13889
rect 31846 13880 31852 13892
rect 31904 13880 31910 13932
rect 31938 13880 31944 13932
rect 31996 13920 32002 13932
rect 32585 13923 32643 13929
rect 32585 13920 32597 13923
rect 31996 13892 32597 13920
rect 31996 13880 32002 13892
rect 32585 13889 32597 13892
rect 32631 13920 32643 13923
rect 32674 13920 32680 13932
rect 32631 13892 32680 13920
rect 32631 13889 32643 13892
rect 32585 13883 32643 13889
rect 32674 13880 32680 13892
rect 32732 13880 32738 13932
rect 32769 13923 32827 13929
rect 32769 13889 32781 13923
rect 32815 13889 32827 13923
rect 32769 13883 32827 13889
rect 34885 13923 34943 13929
rect 34885 13889 34897 13923
rect 34931 13920 34943 13923
rect 35710 13920 35716 13932
rect 34931 13892 35716 13920
rect 34931 13889 34943 13892
rect 34885 13883 34943 13889
rect 26418 13852 26424 13864
rect 26331 13824 26424 13852
rect 26418 13812 26424 13824
rect 26476 13852 26482 13864
rect 27246 13852 27252 13864
rect 26476 13824 27252 13852
rect 26476 13812 26482 13824
rect 27246 13812 27252 13824
rect 27304 13812 27310 13864
rect 29362 13812 29368 13864
rect 29420 13852 29426 13864
rect 29733 13855 29791 13861
rect 29733 13852 29745 13855
rect 29420 13824 29745 13852
rect 29420 13812 29426 13824
rect 29733 13821 29745 13824
rect 29779 13821 29791 13855
rect 29733 13815 29791 13821
rect 29825 13855 29883 13861
rect 29825 13821 29837 13855
rect 29871 13852 29883 13855
rect 30006 13852 30012 13864
rect 29871 13824 30012 13852
rect 29871 13821 29883 13824
rect 29825 13815 29883 13821
rect 28626 13784 28632 13796
rect 26160 13756 28632 13784
rect 26160 13716 26188 13756
rect 28626 13744 28632 13756
rect 28684 13744 28690 13796
rect 28994 13744 29000 13796
rect 29052 13784 29058 13796
rect 29840 13784 29868 13815
rect 30006 13812 30012 13824
rect 30064 13812 30070 13864
rect 32398 13812 32404 13864
rect 32456 13852 32462 13864
rect 32784 13852 32812 13883
rect 35710 13880 35716 13892
rect 35768 13880 35774 13932
rect 36814 13880 36820 13932
rect 36872 13920 36878 13932
rect 37366 13920 37372 13932
rect 36872 13892 37372 13920
rect 36872 13880 36878 13892
rect 37366 13880 37372 13892
rect 37424 13880 37430 13932
rect 38102 13923 38160 13929
rect 38102 13889 38114 13923
rect 38148 13920 38160 13923
rect 38396 13920 38424 13960
rect 39482 13948 39488 13960
rect 39540 13948 39546 14000
rect 41598 13988 41604 14000
rect 41386 13960 41604 13988
rect 38148 13892 38424 13920
rect 38148 13889 38160 13892
rect 38102 13883 38160 13889
rect 38470 13880 38476 13932
rect 38528 13920 38534 13932
rect 39025 13923 39083 13929
rect 39025 13920 39037 13923
rect 38528 13892 39037 13920
rect 38528 13880 38534 13892
rect 39025 13889 39037 13892
rect 39071 13889 39083 13923
rect 39025 13883 39083 13889
rect 39209 13923 39267 13929
rect 39209 13889 39221 13923
rect 39255 13920 39267 13923
rect 41386 13920 41414 13960
rect 41598 13948 41604 13960
rect 41656 13948 41662 14000
rect 41785 13991 41843 13997
rect 41785 13957 41797 13991
rect 41831 13988 41843 13991
rect 41831 13960 43208 13988
rect 41831 13957 41843 13960
rect 41785 13951 41843 13957
rect 41506 13920 41512 13932
rect 39255 13892 41414 13920
rect 41467 13892 41512 13920
rect 39255 13889 39267 13892
rect 39209 13883 39267 13889
rect 41506 13880 41512 13892
rect 41564 13880 41570 13932
rect 41690 13920 41696 13932
rect 41651 13892 41696 13920
rect 41690 13880 41696 13892
rect 41748 13880 41754 13932
rect 41877 13923 41935 13929
rect 41877 13889 41889 13923
rect 41923 13920 41935 13923
rect 42794 13920 42800 13932
rect 41923 13892 42800 13920
rect 41923 13889 41935 13892
rect 41877 13883 41935 13889
rect 42794 13880 42800 13892
rect 42852 13880 42858 13932
rect 43070 13920 43076 13932
rect 43031 13892 43076 13920
rect 43070 13880 43076 13892
rect 43128 13880 43134 13932
rect 43180 13920 43208 13960
rect 43180 13892 44772 13920
rect 32456 13824 32812 13852
rect 32456 13812 32462 13824
rect 34606 13812 34612 13864
rect 34664 13852 34670 13864
rect 34977 13855 35035 13861
rect 34977 13852 34989 13855
rect 34664 13824 34989 13852
rect 34664 13812 34670 13824
rect 34977 13821 34989 13824
rect 35023 13821 35035 13855
rect 35158 13852 35164 13864
rect 35119 13824 35164 13852
rect 34977 13815 35035 13821
rect 35158 13812 35164 13824
rect 35216 13812 35222 13864
rect 38565 13855 38623 13861
rect 38565 13821 38577 13855
rect 38611 13852 38623 13855
rect 38654 13852 38660 13864
rect 38611 13824 38660 13852
rect 38611 13821 38623 13824
rect 38565 13815 38623 13821
rect 38654 13812 38660 13824
rect 38712 13812 38718 13864
rect 43346 13852 43352 13864
rect 43307 13824 43352 13852
rect 43346 13812 43352 13824
rect 43404 13812 43410 13864
rect 44744 13861 44772 13892
rect 44729 13855 44787 13861
rect 44729 13821 44741 13855
rect 44775 13852 44787 13855
rect 57238 13852 57244 13864
rect 44775 13824 57244 13852
rect 44775 13821 44787 13824
rect 44729 13815 44787 13821
rect 57238 13812 57244 13824
rect 57296 13812 57302 13864
rect 29052 13756 29868 13784
rect 30561 13787 30619 13793
rect 29052 13744 29058 13756
rect 30561 13753 30573 13787
rect 30607 13784 30619 13787
rect 30650 13784 30656 13796
rect 30607 13756 30656 13784
rect 30607 13753 30619 13756
rect 30561 13747 30619 13753
rect 30650 13744 30656 13756
rect 30708 13744 30714 13796
rect 38473 13787 38531 13793
rect 38473 13784 38485 13787
rect 31726 13756 38485 13784
rect 22244 13688 26188 13716
rect 22244 13676 22250 13688
rect 26234 13676 26240 13728
rect 26292 13716 26298 13728
rect 31726 13716 31754 13756
rect 38473 13753 38485 13756
rect 38519 13753 38531 13787
rect 38473 13747 38531 13753
rect 41386 13756 42196 13784
rect 34514 13716 34520 13728
rect 26292 13688 31754 13716
rect 34475 13688 34520 13716
rect 26292 13676 26298 13688
rect 34514 13676 34520 13688
rect 34572 13676 34578 13728
rect 34698 13676 34704 13728
rect 34756 13716 34762 13728
rect 41386 13716 41414 13756
rect 42058 13716 42064 13728
rect 34756 13688 41414 13716
rect 42019 13688 42064 13716
rect 34756 13676 34762 13688
rect 42058 13676 42064 13688
rect 42116 13676 42122 13728
rect 42168 13716 42196 13756
rect 49050 13744 49056 13796
rect 49108 13784 49114 13796
rect 55214 13784 55220 13796
rect 49108 13756 55220 13784
rect 49108 13744 49114 13756
rect 55214 13744 55220 13756
rect 55272 13744 55278 13796
rect 43530 13716 43536 13728
rect 42168 13688 43536 13716
rect 43530 13676 43536 13688
rect 43588 13676 43594 13728
rect 1104 13626 58880 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 58880 13626
rect 1104 13552 58880 13574
rect 16022 13472 16028 13524
rect 16080 13512 16086 13524
rect 17310 13512 17316 13524
rect 16080 13484 17316 13512
rect 16080 13472 16086 13484
rect 17310 13472 17316 13484
rect 17368 13512 17374 13524
rect 17862 13512 17868 13524
rect 17368 13484 17868 13512
rect 17368 13472 17374 13484
rect 17862 13472 17868 13484
rect 17920 13512 17926 13524
rect 18874 13512 18880 13524
rect 17920 13484 18880 13512
rect 17920 13472 17926 13484
rect 18874 13472 18880 13484
rect 18932 13472 18938 13524
rect 19334 13472 19340 13524
rect 19392 13512 19398 13524
rect 19521 13515 19579 13521
rect 19521 13512 19533 13515
rect 19392 13484 19533 13512
rect 19392 13472 19398 13484
rect 19521 13481 19533 13484
rect 19567 13481 19579 13515
rect 19521 13475 19579 13481
rect 19794 13472 19800 13524
rect 19852 13512 19858 13524
rect 19852 13484 20300 13512
rect 19852 13472 19858 13484
rect 18414 13404 18420 13456
rect 18472 13444 18478 13456
rect 20272 13444 20300 13484
rect 20714 13472 20720 13524
rect 20772 13512 20778 13524
rect 22189 13515 22247 13521
rect 22189 13512 22201 13515
rect 20772 13484 22201 13512
rect 20772 13472 20778 13484
rect 22189 13481 22201 13484
rect 22235 13481 22247 13515
rect 22189 13475 22247 13481
rect 23934 13472 23940 13524
rect 23992 13512 23998 13524
rect 26418 13512 26424 13524
rect 23992 13484 26424 13512
rect 23992 13472 23998 13484
rect 26418 13472 26424 13484
rect 26476 13472 26482 13524
rect 27338 13512 27344 13524
rect 27299 13484 27344 13512
rect 27338 13472 27344 13484
rect 27396 13472 27402 13524
rect 27890 13472 27896 13524
rect 27948 13512 27954 13524
rect 28261 13515 28319 13521
rect 28261 13512 28273 13515
rect 27948 13484 28273 13512
rect 27948 13472 27954 13484
rect 28261 13481 28273 13484
rect 28307 13481 28319 13515
rect 28261 13475 28319 13481
rect 31570 13472 31576 13524
rect 31628 13512 31634 13524
rect 38194 13512 38200 13524
rect 31628 13484 38200 13512
rect 31628 13472 31634 13484
rect 38194 13472 38200 13484
rect 38252 13472 38258 13524
rect 38286 13472 38292 13524
rect 38344 13512 38350 13524
rect 38344 13484 43208 13512
rect 38344 13472 38350 13484
rect 35802 13444 35808 13456
rect 18472 13416 20208 13444
rect 20272 13416 35808 13444
rect 18472 13404 18478 13416
rect 9306 13376 9312 13388
rect 9267 13348 9312 13376
rect 9306 13336 9312 13348
rect 9364 13336 9370 13388
rect 9585 13379 9643 13385
rect 9585 13345 9597 13379
rect 9631 13376 9643 13379
rect 9674 13376 9680 13388
rect 9631 13348 9680 13376
rect 9631 13345 9643 13348
rect 9585 13339 9643 13345
rect 9674 13336 9680 13348
rect 9732 13336 9738 13388
rect 14274 13376 14280 13388
rect 14235 13348 14280 13376
rect 14274 13336 14280 13348
rect 14332 13336 14338 13388
rect 16298 13336 16304 13388
rect 16356 13376 16362 13388
rect 16356 13348 16896 13376
rect 16356 13336 16362 13348
rect 1578 13308 1584 13320
rect 1539 13280 1584 13308
rect 1578 13268 1584 13280
rect 1636 13268 1642 13320
rect 11422 13308 11428 13320
rect 11383 13280 11428 13308
rect 11422 13268 11428 13280
rect 11480 13268 11486 13320
rect 13538 13268 13544 13320
rect 13596 13308 13602 13320
rect 14553 13311 14611 13317
rect 14553 13308 14565 13311
rect 13596 13280 14565 13308
rect 13596 13268 13602 13280
rect 14553 13277 14565 13280
rect 14599 13277 14611 13311
rect 14553 13271 14611 13277
rect 16577 13311 16635 13317
rect 16577 13277 16589 13311
rect 16623 13308 16635 13311
rect 16758 13308 16764 13320
rect 16623 13280 16764 13308
rect 16623 13277 16635 13280
rect 16577 13271 16635 13277
rect 16758 13268 16764 13280
rect 16816 13268 16822 13320
rect 16868 13308 16896 13348
rect 17218 13336 17224 13388
rect 17276 13376 17282 13388
rect 17862 13376 17868 13388
rect 17276 13348 17868 13376
rect 17276 13336 17282 13348
rect 17862 13336 17868 13348
rect 17920 13336 17926 13388
rect 18138 13376 18144 13388
rect 18099 13348 18144 13376
rect 18138 13336 18144 13348
rect 18196 13336 18202 13388
rect 19981 13379 20039 13385
rect 19981 13345 19993 13379
rect 20027 13376 20039 13379
rect 20070 13376 20076 13388
rect 20027 13348 20076 13376
rect 20027 13345 20039 13348
rect 19981 13339 20039 13345
rect 20070 13336 20076 13348
rect 20128 13336 20134 13388
rect 20180 13376 20208 13416
rect 35802 13404 35808 13416
rect 35860 13404 35866 13456
rect 38930 13404 38936 13456
rect 38988 13444 38994 13456
rect 42797 13447 42855 13453
rect 38988 13416 42656 13444
rect 38988 13404 38994 13416
rect 23474 13376 23480 13388
rect 20180 13348 23480 13376
rect 23474 13336 23480 13348
rect 23532 13336 23538 13388
rect 25038 13376 25044 13388
rect 24999 13348 25044 13376
rect 25038 13336 25044 13348
rect 25096 13336 25102 13388
rect 31570 13376 31576 13388
rect 25976 13348 31576 13376
rect 20993 13311 21051 13317
rect 16868 13280 20944 13308
rect 1854 13240 1860 13252
rect 1815 13212 1860 13240
rect 1854 13200 1860 13212
rect 1912 13200 1918 13252
rect 10965 13243 11023 13249
rect 10965 13209 10977 13243
rect 11011 13240 11023 13243
rect 19426 13240 19432 13252
rect 11011 13212 14412 13240
rect 11011 13209 11023 13212
rect 10965 13203 11023 13209
rect 11238 13132 11244 13184
rect 11296 13172 11302 13184
rect 12621 13175 12679 13181
rect 12621 13172 12633 13175
rect 11296 13144 12633 13172
rect 11296 13132 11302 13144
rect 12621 13141 12633 13144
rect 12667 13141 12679 13175
rect 14384 13172 14412 13212
rect 15212 13212 19432 13240
rect 15212 13172 15240 13212
rect 19426 13200 19432 13212
rect 19484 13200 19490 13252
rect 20073 13243 20131 13249
rect 20073 13209 20085 13243
rect 20119 13209 20131 13243
rect 20916 13240 20944 13280
rect 20993 13277 21005 13311
rect 21039 13308 21051 13311
rect 21082 13308 21088 13320
rect 21039 13280 21088 13308
rect 21039 13277 21051 13280
rect 20993 13271 21051 13277
rect 21082 13268 21088 13280
rect 21140 13268 21146 13320
rect 23842 13308 23848 13320
rect 21192 13280 23848 13308
rect 21192 13240 21220 13280
rect 23842 13268 23848 13280
rect 23900 13268 23906 13320
rect 24026 13308 24032 13320
rect 23987 13280 24032 13308
rect 24026 13268 24032 13280
rect 24084 13268 24090 13320
rect 24670 13308 24676 13320
rect 24228 13280 24676 13308
rect 20916 13212 21220 13240
rect 20073 13203 20131 13209
rect 14384 13144 15240 13172
rect 12621 13135 12679 13141
rect 15562 13132 15568 13184
rect 15620 13172 15626 13184
rect 15657 13175 15715 13181
rect 15657 13172 15669 13175
rect 15620 13144 15669 13172
rect 15620 13132 15626 13144
rect 15657 13141 15669 13144
rect 15703 13141 15715 13175
rect 15657 13135 15715 13141
rect 15930 13132 15936 13184
rect 15988 13172 15994 13184
rect 19794 13172 19800 13184
rect 15988 13144 19800 13172
rect 15988 13132 15994 13144
rect 19794 13132 19800 13144
rect 19852 13132 19858 13184
rect 19978 13172 19984 13184
rect 19939 13144 19984 13172
rect 19978 13132 19984 13144
rect 20036 13132 20042 13184
rect 20088 13172 20116 13203
rect 23382 13200 23388 13252
rect 23440 13240 23446 13252
rect 23937 13243 23995 13249
rect 23937 13240 23949 13243
rect 23440 13212 23949 13240
rect 23440 13200 23446 13212
rect 23937 13209 23949 13212
rect 23983 13209 23995 13243
rect 23937 13203 23995 13209
rect 21082 13172 21088 13184
rect 20088 13144 21088 13172
rect 21082 13132 21088 13144
rect 21140 13132 21146 13184
rect 22002 13132 22008 13184
rect 22060 13172 22066 13184
rect 24228 13172 24256 13280
rect 24670 13268 24676 13280
rect 24728 13308 24734 13320
rect 24765 13311 24823 13317
rect 24765 13308 24777 13311
rect 24728 13280 24777 13308
rect 24728 13268 24734 13280
rect 24765 13277 24777 13280
rect 24811 13277 24823 13311
rect 24765 13271 24823 13277
rect 24857 13311 24915 13317
rect 24857 13277 24869 13311
rect 24903 13308 24915 13311
rect 24946 13308 24952 13320
rect 24903 13280 24952 13308
rect 24903 13277 24915 13280
rect 24857 13271 24915 13277
rect 24946 13268 24952 13280
rect 25004 13268 25010 13320
rect 25130 13308 25136 13320
rect 25091 13280 25136 13308
rect 25130 13268 25136 13280
rect 25188 13268 25194 13320
rect 24581 13243 24639 13249
rect 24581 13209 24593 13243
rect 24627 13240 24639 13243
rect 25976 13240 26004 13348
rect 31570 13336 31576 13348
rect 31628 13336 31634 13388
rect 41598 13376 41604 13388
rect 31864 13348 33180 13376
rect 28258 13308 28264 13320
rect 28219 13280 28264 13308
rect 28258 13268 28264 13280
rect 28316 13268 28322 13320
rect 28445 13311 28503 13317
rect 28445 13277 28457 13311
rect 28491 13308 28503 13311
rect 29086 13308 29092 13320
rect 28491 13280 29092 13308
rect 28491 13277 28503 13280
rect 28445 13271 28503 13277
rect 29086 13268 29092 13280
rect 29144 13268 29150 13320
rect 31864 13317 31892 13348
rect 31849 13311 31907 13317
rect 31849 13277 31861 13311
rect 31895 13277 31907 13311
rect 32217 13311 32275 13317
rect 32217 13308 32229 13311
rect 31849 13271 31907 13277
rect 31956 13280 32229 13308
rect 24627 13212 26004 13240
rect 26053 13243 26111 13249
rect 24627 13209 24639 13212
rect 24581 13203 24639 13209
rect 26053 13209 26065 13243
rect 26099 13240 26111 13243
rect 28626 13240 28632 13252
rect 26099 13212 28632 13240
rect 26099 13209 26111 13212
rect 26053 13203 26111 13209
rect 28626 13200 28632 13212
rect 28684 13200 28690 13252
rect 31570 13200 31576 13252
rect 31628 13240 31634 13252
rect 31956 13240 31984 13280
rect 32217 13277 32229 13280
rect 32263 13308 32275 13311
rect 32490 13308 32496 13320
rect 32263 13280 32496 13308
rect 32263 13277 32275 13280
rect 32217 13271 32275 13277
rect 32490 13268 32496 13280
rect 32548 13268 32554 13320
rect 33152 13308 33180 13348
rect 35912 13348 41604 13376
rect 35912 13308 35940 13348
rect 41598 13336 41604 13348
rect 41656 13336 41662 13388
rect 42628 13320 42656 13416
rect 42797 13413 42809 13447
rect 42843 13413 42855 13447
rect 43180 13444 43208 13484
rect 43254 13472 43260 13524
rect 43312 13512 43318 13524
rect 43625 13515 43683 13521
rect 43625 13512 43637 13515
rect 43312 13484 43637 13512
rect 43312 13472 43318 13484
rect 43625 13481 43637 13484
rect 43671 13481 43683 13515
rect 43625 13475 43683 13481
rect 48406 13444 48412 13456
rect 43180 13416 48412 13444
rect 42797 13407 42855 13413
rect 42812 13376 42840 13407
rect 48406 13404 48412 13416
rect 48464 13404 48470 13456
rect 58158 13376 58164 13388
rect 42812 13348 43484 13376
rect 58119 13348 58164 13376
rect 36262 13308 36268 13320
rect 33152 13280 35940 13308
rect 36223 13280 36268 13308
rect 36262 13268 36268 13280
rect 36320 13268 36326 13320
rect 36354 13268 36360 13320
rect 36412 13308 36418 13320
rect 36449 13311 36507 13317
rect 36449 13308 36461 13311
rect 36412 13280 36461 13308
rect 36412 13268 36418 13280
rect 36449 13277 36461 13280
rect 36495 13277 36507 13311
rect 36449 13271 36507 13277
rect 37108 13280 37504 13308
rect 31628 13212 31984 13240
rect 32033 13243 32091 13249
rect 31628 13200 31634 13212
rect 32033 13209 32045 13243
rect 32079 13209 32091 13243
rect 32033 13203 32091 13209
rect 22060 13144 24256 13172
rect 22060 13132 22066 13144
rect 24946 13132 24952 13184
rect 25004 13172 25010 13184
rect 29546 13172 29552 13184
rect 25004 13144 29552 13172
rect 25004 13132 25010 13144
rect 29546 13132 29552 13144
rect 29604 13132 29610 13184
rect 32048 13172 32076 13203
rect 32122 13200 32128 13252
rect 32180 13240 32186 13252
rect 32582 13240 32588 13252
rect 32180 13212 32225 13240
rect 32324 13212 32588 13240
rect 32180 13200 32186 13212
rect 32324 13172 32352 13212
rect 32582 13200 32588 13212
rect 32640 13200 32646 13252
rect 35986 13200 35992 13252
rect 36044 13240 36050 13252
rect 37108 13240 37136 13280
rect 36044 13212 37136 13240
rect 37185 13243 37243 13249
rect 36044 13200 36050 13212
rect 37185 13209 37197 13243
rect 37231 13209 37243 13243
rect 37185 13203 37243 13209
rect 32048 13144 32352 13172
rect 32401 13175 32459 13181
rect 32401 13141 32413 13175
rect 32447 13172 32459 13175
rect 32490 13172 32496 13184
rect 32447 13144 32496 13172
rect 32447 13141 32459 13144
rect 32401 13135 32459 13141
rect 32490 13132 32496 13144
rect 32548 13132 32554 13184
rect 32858 13132 32864 13184
rect 32916 13172 32922 13184
rect 34698 13172 34704 13184
rect 32916 13144 34704 13172
rect 32916 13132 32922 13144
rect 34698 13132 34704 13144
rect 34756 13132 34762 13184
rect 36630 13172 36636 13184
rect 36591 13144 36636 13172
rect 36630 13132 36636 13144
rect 36688 13132 36694 13184
rect 37090 13132 37096 13184
rect 37148 13172 37154 13184
rect 37200 13172 37228 13203
rect 37148 13144 37228 13172
rect 37148 13132 37154 13144
rect 37274 13132 37280 13184
rect 37332 13172 37338 13184
rect 37476 13172 37504 13280
rect 37826 13268 37832 13320
rect 37884 13308 37890 13320
rect 38105 13311 38163 13317
rect 38105 13308 38117 13311
rect 37884 13280 38117 13308
rect 37884 13268 37890 13280
rect 38105 13277 38117 13280
rect 38151 13277 38163 13311
rect 38654 13308 38660 13320
rect 38615 13280 38660 13308
rect 38105 13271 38163 13277
rect 38654 13268 38660 13280
rect 38712 13268 38718 13320
rect 41414 13268 41420 13320
rect 41472 13308 41478 13320
rect 42245 13311 42303 13317
rect 42245 13308 42257 13311
rect 41472 13280 42257 13308
rect 41472 13268 41478 13280
rect 42245 13277 42257 13280
rect 42291 13277 42303 13311
rect 42610 13308 42616 13320
rect 42571 13280 42616 13308
rect 42245 13271 42303 13277
rect 42610 13268 42616 13280
rect 42668 13268 42674 13320
rect 43162 13268 43168 13320
rect 43220 13308 43226 13320
rect 43456 13317 43484 13348
rect 58158 13336 58164 13348
rect 58216 13336 58222 13388
rect 43257 13311 43315 13317
rect 43257 13308 43269 13311
rect 43220 13280 43269 13308
rect 43220 13268 43226 13280
rect 43257 13277 43269 13280
rect 43303 13277 43315 13311
rect 43257 13271 43315 13277
rect 43441 13311 43499 13317
rect 43441 13277 43453 13311
rect 43487 13277 43499 13311
rect 56962 13308 56968 13320
rect 56923 13280 56968 13308
rect 43441 13271 43499 13277
rect 56962 13268 56968 13280
rect 57020 13268 57026 13320
rect 57882 13308 57888 13320
rect 57843 13280 57888 13308
rect 57882 13268 57888 13280
rect 57940 13268 57946 13320
rect 38470 13200 38476 13252
rect 38528 13240 38534 13252
rect 39298 13240 39304 13252
rect 38528 13212 39304 13240
rect 38528 13200 38534 13212
rect 39298 13200 39304 13212
rect 39356 13200 39362 13252
rect 42429 13243 42487 13249
rect 42429 13209 42441 13243
rect 42475 13209 42487 13243
rect 42429 13203 42487 13209
rect 42521 13243 42579 13249
rect 42521 13209 42533 13243
rect 42567 13240 42579 13243
rect 44542 13240 44548 13252
rect 42567 13212 44548 13240
rect 42567 13209 42579 13212
rect 42521 13203 42579 13209
rect 38197 13175 38255 13181
rect 38197 13172 38209 13175
rect 37332 13144 37377 13172
rect 37476 13144 38209 13172
rect 37332 13132 37338 13144
rect 38197 13141 38209 13144
rect 38243 13172 38255 13175
rect 41690 13172 41696 13184
rect 38243 13144 41696 13172
rect 38243 13141 38255 13144
rect 38197 13135 38255 13141
rect 41690 13132 41696 13144
rect 41748 13172 41754 13184
rect 42444 13172 42472 13203
rect 44542 13200 44548 13212
rect 44600 13200 44606 13252
rect 55858 13200 55864 13252
rect 55916 13240 55922 13252
rect 57241 13243 57299 13249
rect 57241 13240 57253 13243
rect 55916 13212 57253 13240
rect 55916 13200 55922 13212
rect 57241 13209 57253 13212
rect 57287 13209 57299 13243
rect 57241 13203 57299 13209
rect 41748 13144 42472 13172
rect 41748 13132 41754 13144
rect 42610 13132 42616 13184
rect 42668 13172 42674 13184
rect 43714 13172 43720 13184
rect 42668 13144 43720 13172
rect 42668 13132 42674 13144
rect 43714 13132 43720 13144
rect 43772 13172 43778 13184
rect 44450 13172 44456 13184
rect 43772 13144 44456 13172
rect 43772 13132 43778 13144
rect 44450 13132 44456 13144
rect 44508 13132 44514 13184
rect 1104 13082 58880 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 58880 13082
rect 1104 13008 58880 13030
rect 9766 12928 9772 12980
rect 9824 12968 9830 12980
rect 9953 12971 10011 12977
rect 9953 12968 9965 12971
rect 9824 12940 9965 12968
rect 9824 12928 9830 12940
rect 9953 12937 9965 12940
rect 9999 12937 10011 12971
rect 11146 12968 11152 12980
rect 11107 12940 11152 12968
rect 9953 12931 10011 12937
rect 11146 12928 11152 12940
rect 11204 12928 11210 12980
rect 13538 12968 13544 12980
rect 13499 12940 13544 12968
rect 13538 12928 13544 12940
rect 13596 12928 13602 12980
rect 15378 12968 15384 12980
rect 15339 12940 15384 12968
rect 15378 12928 15384 12940
rect 15436 12928 15442 12980
rect 17218 12928 17224 12980
rect 17276 12968 17282 12980
rect 17276 12940 17321 12968
rect 17276 12928 17282 12940
rect 17770 12928 17776 12980
rect 17828 12968 17834 12980
rect 18138 12968 18144 12980
rect 17828 12940 18144 12968
rect 17828 12928 17834 12940
rect 18138 12928 18144 12940
rect 18196 12928 18202 12980
rect 23014 12968 23020 12980
rect 21008 12940 23020 12968
rect 11882 12900 11888 12912
rect 11843 12872 11888 12900
rect 11882 12860 11888 12872
rect 11940 12860 11946 12912
rect 11974 12860 11980 12912
rect 12032 12900 12038 12912
rect 12161 12903 12219 12909
rect 12161 12900 12173 12903
rect 12032 12872 12173 12900
rect 12032 12860 12038 12872
rect 12161 12869 12173 12872
rect 12207 12869 12219 12903
rect 12161 12863 12219 12869
rect 12253 12903 12311 12909
rect 12253 12869 12265 12903
rect 12299 12900 12311 12903
rect 12299 12872 13124 12900
rect 12299 12869 12311 12872
rect 12253 12863 12311 12869
rect 9585 12835 9643 12841
rect 9585 12801 9597 12835
rect 9631 12832 9643 12835
rect 12066 12832 12072 12844
rect 9631 12804 12072 12832
rect 9631 12801 9643 12804
rect 9585 12795 9643 12801
rect 12066 12792 12072 12804
rect 12124 12792 12130 12844
rect 12618 12832 12624 12844
rect 12579 12804 12624 12832
rect 12618 12792 12624 12804
rect 12676 12792 12682 12844
rect 8846 12724 8852 12776
rect 8904 12764 8910 12776
rect 9490 12764 9496 12776
rect 8904 12736 9496 12764
rect 8904 12724 8910 12736
rect 9490 12724 9496 12736
rect 9548 12724 9554 12776
rect 10689 12767 10747 12773
rect 10689 12733 10701 12767
rect 10735 12764 10747 12767
rect 12636 12764 12664 12792
rect 13096 12776 13124 12872
rect 15194 12860 15200 12912
rect 15252 12900 15258 12912
rect 15930 12900 15936 12912
rect 15252 12872 15936 12900
rect 15252 12860 15258 12872
rect 15930 12860 15936 12872
rect 15988 12860 15994 12912
rect 16853 12903 16911 12909
rect 16853 12869 16865 12903
rect 16899 12900 16911 12903
rect 16899 12872 17816 12900
rect 16899 12869 16911 12872
rect 16853 12863 16911 12869
rect 13998 12832 14004 12844
rect 13959 12804 14004 12832
rect 13998 12792 14004 12804
rect 14056 12792 14062 12844
rect 17037 12835 17095 12841
rect 17037 12801 17049 12835
rect 17083 12801 17095 12835
rect 17310 12832 17316 12844
rect 17271 12804 17316 12832
rect 17037 12795 17095 12801
rect 13078 12764 13084 12776
rect 10735 12736 12664 12764
rect 13039 12736 13084 12764
rect 10735 12733 10747 12736
rect 10689 12727 10747 12733
rect 13078 12724 13084 12736
rect 13136 12724 13142 12776
rect 10965 12699 11023 12705
rect 10965 12665 10977 12699
rect 11011 12696 11023 12699
rect 11238 12696 11244 12708
rect 11011 12668 11244 12696
rect 11011 12665 11023 12668
rect 10965 12659 11023 12665
rect 11238 12656 11244 12668
rect 11296 12656 11302 12708
rect 13449 12699 13507 12705
rect 13449 12665 13461 12699
rect 13495 12696 13507 12699
rect 16666 12696 16672 12708
rect 13495 12668 16672 12696
rect 13495 12665 13507 12668
rect 13449 12659 13507 12665
rect 16666 12656 16672 12668
rect 16724 12656 16730 12708
rect 17052 12696 17080 12795
rect 17310 12792 17316 12804
rect 17368 12792 17374 12844
rect 17788 12841 17816 12872
rect 17862 12860 17868 12912
rect 17920 12900 17926 12912
rect 19610 12900 19616 12912
rect 17920 12872 19616 12900
rect 17920 12860 17926 12872
rect 19610 12860 19616 12872
rect 19668 12860 19674 12912
rect 21008 12841 21036 12940
rect 23014 12928 23020 12940
rect 23072 12928 23078 12980
rect 23474 12928 23480 12980
rect 23532 12968 23538 12980
rect 25130 12968 25136 12980
rect 23532 12940 25136 12968
rect 23532 12928 23538 12940
rect 25130 12928 25136 12940
rect 25188 12968 25194 12980
rect 26142 12968 26148 12980
rect 25188 12940 26148 12968
rect 25188 12928 25194 12940
rect 26142 12928 26148 12940
rect 26200 12928 26206 12980
rect 26234 12928 26240 12980
rect 26292 12968 26298 12980
rect 28534 12968 28540 12980
rect 26292 12940 28540 12968
rect 26292 12928 26298 12940
rect 28534 12928 28540 12940
rect 28592 12928 28598 12980
rect 37182 12968 37188 12980
rect 28644 12940 37188 12968
rect 28644 12912 28672 12940
rect 37182 12928 37188 12940
rect 37240 12928 37246 12980
rect 40862 12928 40868 12980
rect 40920 12968 40926 12980
rect 42794 12968 42800 12980
rect 40920 12940 42800 12968
rect 40920 12928 40926 12940
rect 42794 12928 42800 12940
rect 42852 12928 42858 12980
rect 43165 12971 43223 12977
rect 43165 12937 43177 12971
rect 43211 12968 43223 12971
rect 43346 12968 43352 12980
rect 43211 12940 43352 12968
rect 43211 12937 43223 12940
rect 43165 12931 43223 12937
rect 43346 12928 43352 12940
rect 43404 12928 43410 12980
rect 46658 12928 46664 12980
rect 46716 12968 46722 12980
rect 57882 12968 57888 12980
rect 46716 12940 57888 12968
rect 46716 12928 46722 12940
rect 57882 12928 57888 12940
rect 57940 12928 57946 12980
rect 27798 12900 27804 12912
rect 22020 12872 27804 12900
rect 22020 12841 22048 12872
rect 27798 12860 27804 12872
rect 27856 12860 27862 12912
rect 28626 12900 28632 12912
rect 28587 12872 28632 12900
rect 28626 12860 28632 12872
rect 28684 12860 28690 12912
rect 29730 12860 29736 12912
rect 29788 12900 29794 12912
rect 30285 12903 30343 12909
rect 30285 12900 30297 12903
rect 29788 12872 30297 12900
rect 29788 12860 29794 12872
rect 30285 12869 30297 12872
rect 30331 12900 30343 12903
rect 33226 12900 33232 12912
rect 30331 12872 33232 12900
rect 30331 12869 30343 12872
rect 30285 12863 30343 12869
rect 33226 12860 33232 12872
rect 33284 12900 33290 12912
rect 35986 12900 35992 12912
rect 33284 12872 33916 12900
rect 35947 12872 35992 12900
rect 33284 12860 33290 12872
rect 17773 12835 17831 12841
rect 17773 12801 17785 12835
rect 17819 12801 17831 12835
rect 17773 12795 17831 12801
rect 20993 12835 21051 12841
rect 20993 12801 21005 12835
rect 21039 12801 21051 12835
rect 20993 12795 21051 12801
rect 22005 12835 22063 12841
rect 22005 12801 22017 12835
rect 22051 12801 22063 12835
rect 22005 12795 22063 12801
rect 22554 12792 22560 12844
rect 22612 12832 22618 12844
rect 23014 12832 23020 12844
rect 22612 12804 23020 12832
rect 22612 12792 22618 12804
rect 23014 12792 23020 12804
rect 23072 12792 23078 12844
rect 24762 12832 24768 12844
rect 24723 12804 24768 12832
rect 24762 12792 24768 12804
rect 24820 12792 24826 12844
rect 25032 12835 25090 12841
rect 25032 12801 25044 12835
rect 25078 12832 25090 12835
rect 25406 12832 25412 12844
rect 25078 12804 25412 12832
rect 25078 12801 25090 12804
rect 25032 12795 25090 12801
rect 25406 12792 25412 12804
rect 25464 12792 25470 12844
rect 26142 12792 26148 12844
rect 26200 12832 26206 12844
rect 27341 12835 27399 12841
rect 27341 12832 27353 12835
rect 26200 12804 27353 12832
rect 26200 12792 26206 12804
rect 27341 12801 27353 12804
rect 27387 12801 27399 12835
rect 27341 12795 27399 12801
rect 17402 12724 17408 12776
rect 17460 12764 17466 12776
rect 20806 12764 20812 12776
rect 17460 12736 20812 12764
rect 17460 12724 17466 12736
rect 20806 12724 20812 12736
rect 20864 12724 20870 12776
rect 20898 12724 20904 12776
rect 20956 12764 20962 12776
rect 21177 12767 21235 12773
rect 21177 12764 21189 12767
rect 20956 12736 21189 12764
rect 20956 12724 20962 12736
rect 21177 12733 21189 12736
rect 21223 12733 21235 12767
rect 27356 12764 27384 12795
rect 27430 12792 27436 12844
rect 27488 12832 27494 12844
rect 27488 12804 27533 12832
rect 27488 12792 27494 12804
rect 27614 12792 27620 12844
rect 27672 12832 27678 12844
rect 30374 12832 30380 12844
rect 27672 12804 30380 12832
rect 27672 12792 27678 12804
rect 30374 12792 30380 12804
rect 30432 12792 30438 12844
rect 30926 12832 30932 12844
rect 30887 12804 30932 12832
rect 30926 12792 30932 12804
rect 30984 12792 30990 12844
rect 31110 12832 31116 12844
rect 31071 12804 31116 12832
rect 31110 12792 31116 12804
rect 31168 12792 31174 12844
rect 31205 12835 31263 12841
rect 31205 12801 31217 12835
rect 31251 12832 31263 12835
rect 31386 12832 31392 12844
rect 31251 12804 31392 12832
rect 31251 12801 31263 12804
rect 31205 12795 31263 12801
rect 31386 12792 31392 12804
rect 31444 12792 31450 12844
rect 32674 12832 32680 12844
rect 32635 12804 32680 12832
rect 32674 12792 32680 12804
rect 32732 12792 32738 12844
rect 32950 12832 32956 12844
rect 32911 12804 32956 12832
rect 32950 12792 32956 12804
rect 33008 12792 33014 12844
rect 33888 12841 33916 12872
rect 35986 12860 35992 12872
rect 36044 12860 36050 12912
rect 36081 12903 36139 12909
rect 36081 12869 36093 12903
rect 36127 12900 36139 12903
rect 38010 12900 38016 12912
rect 36127 12872 38016 12900
rect 36127 12869 36139 12872
rect 36081 12863 36139 12869
rect 38010 12860 38016 12872
rect 38068 12860 38074 12912
rect 38194 12860 38200 12912
rect 38252 12900 38258 12912
rect 43530 12900 43536 12912
rect 38252 12872 43536 12900
rect 38252 12860 38258 12872
rect 43530 12860 43536 12872
rect 43588 12860 43594 12912
rect 33873 12835 33931 12841
rect 33873 12801 33885 12835
rect 33919 12832 33931 12835
rect 33962 12832 33968 12844
rect 33919 12804 33968 12832
rect 33919 12801 33931 12804
rect 33873 12795 33931 12801
rect 33962 12792 33968 12804
rect 34020 12792 34026 12844
rect 34140 12835 34198 12841
rect 34140 12801 34152 12835
rect 34186 12832 34198 12835
rect 34514 12832 34520 12844
rect 34186 12804 34520 12832
rect 34186 12801 34198 12804
rect 34140 12795 34198 12801
rect 34514 12792 34520 12804
rect 34572 12792 34578 12844
rect 34698 12792 34704 12844
rect 34756 12832 34762 12844
rect 35802 12832 35808 12844
rect 34756 12804 34928 12832
rect 35763 12804 35808 12832
rect 34756 12792 34762 12804
rect 28077 12767 28135 12773
rect 28077 12764 28089 12767
rect 27356 12736 28089 12764
rect 21177 12727 21235 12733
rect 28077 12733 28089 12736
rect 28123 12764 28135 12767
rect 32769 12767 32827 12773
rect 28123 12736 31248 12764
rect 28123 12733 28135 12736
rect 28077 12727 28135 12733
rect 19426 12696 19432 12708
rect 17052 12668 19432 12696
rect 19426 12656 19432 12668
rect 19484 12656 19490 12708
rect 19518 12656 19524 12708
rect 19576 12696 19582 12708
rect 19576 12668 23796 12696
rect 19576 12656 19582 12668
rect 15010 12588 15016 12640
rect 15068 12628 15074 12640
rect 18969 12631 19027 12637
rect 18969 12628 18981 12631
rect 15068 12600 18981 12628
rect 15068 12588 15074 12600
rect 18969 12597 18981 12600
rect 19015 12597 19027 12631
rect 18969 12591 19027 12597
rect 21450 12588 21456 12640
rect 21508 12628 21514 12640
rect 23201 12631 23259 12637
rect 23201 12628 23213 12631
rect 21508 12600 23213 12628
rect 21508 12588 21514 12600
rect 23201 12597 23213 12600
rect 23247 12597 23259 12631
rect 23768 12628 23796 12668
rect 27062 12656 27068 12708
rect 27120 12696 27126 12708
rect 28258 12696 28264 12708
rect 27120 12668 28264 12696
rect 27120 12656 27126 12668
rect 28258 12656 28264 12668
rect 28316 12696 28322 12708
rect 31220 12696 31248 12736
rect 32769 12733 32781 12767
rect 32815 12764 32827 12767
rect 32858 12764 32864 12776
rect 32815 12736 32864 12764
rect 32815 12733 32827 12736
rect 32769 12727 32827 12733
rect 32858 12724 32864 12736
rect 32916 12724 32922 12776
rect 33410 12764 33416 12776
rect 33371 12736 33416 12764
rect 33410 12724 33416 12736
rect 33468 12724 33474 12776
rect 34900 12764 34928 12804
rect 35802 12792 35808 12804
rect 35860 12792 35866 12844
rect 36173 12835 36231 12841
rect 36173 12801 36185 12835
rect 36219 12832 36231 12835
rect 36262 12832 36268 12844
rect 36219 12804 36268 12832
rect 36219 12801 36231 12804
rect 36173 12795 36231 12801
rect 36262 12792 36268 12804
rect 36320 12792 36326 12844
rect 36446 12792 36452 12844
rect 36504 12832 36510 12844
rect 37826 12832 37832 12844
rect 36504 12804 37832 12832
rect 36504 12792 36510 12804
rect 37826 12792 37832 12804
rect 37884 12792 37890 12844
rect 41782 12832 41788 12844
rect 41743 12804 41788 12832
rect 41782 12792 41788 12804
rect 41840 12792 41846 12844
rect 42058 12792 42064 12844
rect 42116 12832 42122 12844
rect 42981 12835 43039 12841
rect 42981 12832 42993 12835
rect 42116 12804 42993 12832
rect 42116 12792 42122 12804
rect 42981 12801 42993 12804
rect 43027 12801 43039 12835
rect 42981 12795 43039 12801
rect 37090 12764 37096 12776
rect 34900 12736 37096 12764
rect 37090 12724 37096 12736
rect 37148 12724 37154 12776
rect 41138 12724 41144 12776
rect 41196 12764 41202 12776
rect 42797 12767 42855 12773
rect 42797 12764 42809 12767
rect 41196 12736 42809 12764
rect 41196 12724 41202 12736
rect 42797 12733 42809 12736
rect 42843 12764 42855 12767
rect 43162 12764 43168 12776
rect 42843 12736 43168 12764
rect 42843 12733 42855 12736
rect 42797 12727 42855 12733
rect 43162 12724 43168 12736
rect 43220 12724 43226 12776
rect 31938 12696 31944 12708
rect 28316 12668 31156 12696
rect 31220 12668 31944 12696
rect 28316 12656 28322 12668
rect 25498 12628 25504 12640
rect 23768 12600 25504 12628
rect 23201 12591 23259 12597
rect 25498 12588 25504 12600
rect 25556 12588 25562 12640
rect 25866 12588 25872 12640
rect 25924 12628 25930 12640
rect 26145 12631 26203 12637
rect 26145 12628 26157 12631
rect 25924 12600 26157 12628
rect 25924 12588 25930 12600
rect 26145 12597 26157 12600
rect 26191 12597 26203 12631
rect 26145 12591 26203 12597
rect 26602 12588 26608 12640
rect 26660 12628 26666 12640
rect 27341 12631 27399 12637
rect 27341 12628 27353 12631
rect 26660 12600 27353 12628
rect 26660 12588 26666 12600
rect 27341 12597 27353 12600
rect 27387 12597 27399 12631
rect 27706 12628 27712 12640
rect 27667 12600 27712 12628
rect 27341 12591 27399 12597
rect 27706 12588 27712 12600
rect 27764 12588 27770 12640
rect 28166 12588 28172 12640
rect 28224 12628 28230 12640
rect 28534 12628 28540 12640
rect 28224 12600 28540 12628
rect 28224 12588 28230 12600
rect 28534 12588 28540 12600
rect 28592 12588 28598 12640
rect 30929 12631 30987 12637
rect 30929 12597 30941 12631
rect 30975 12628 30987 12631
rect 31018 12628 31024 12640
rect 30975 12600 31024 12628
rect 30975 12597 30987 12600
rect 30929 12591 30987 12597
rect 31018 12588 31024 12600
rect 31076 12588 31082 12640
rect 31128 12628 31156 12668
rect 31938 12656 31944 12668
rect 31996 12656 32002 12708
rect 36354 12696 36360 12708
rect 36315 12668 36360 12696
rect 36354 12656 36360 12668
rect 36412 12656 36418 12708
rect 41969 12699 42027 12705
rect 41969 12665 41981 12699
rect 42015 12696 42027 12699
rect 43438 12696 43444 12708
rect 42015 12668 43444 12696
rect 42015 12665 42027 12668
rect 41969 12659 42027 12665
rect 31846 12628 31852 12640
rect 31128 12600 31852 12628
rect 31846 12588 31852 12600
rect 31904 12588 31910 12640
rect 33226 12588 33232 12640
rect 33284 12628 33290 12640
rect 33502 12628 33508 12640
rect 33284 12600 33508 12628
rect 33284 12588 33290 12600
rect 33502 12588 33508 12600
rect 33560 12588 33566 12640
rect 34514 12588 34520 12640
rect 34572 12628 34578 12640
rect 35253 12631 35311 12637
rect 35253 12628 35265 12631
rect 34572 12600 35265 12628
rect 34572 12588 34578 12600
rect 35253 12597 35265 12600
rect 35299 12597 35311 12631
rect 35253 12591 35311 12597
rect 37090 12588 37096 12640
rect 37148 12628 37154 12640
rect 41984 12628 42012 12659
rect 43438 12656 43444 12668
rect 43496 12656 43502 12708
rect 37148 12600 42012 12628
rect 37148 12588 37154 12600
rect 1104 12538 58880 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 58880 12538
rect 1104 12464 58880 12486
rect 2222 12424 2228 12436
rect 2183 12396 2228 12424
rect 2222 12384 2228 12396
rect 2280 12384 2286 12436
rect 10134 12384 10140 12436
rect 10192 12424 10198 12436
rect 10873 12427 10931 12433
rect 10873 12424 10885 12427
rect 10192 12396 10885 12424
rect 10192 12384 10198 12396
rect 10873 12393 10885 12396
rect 10919 12393 10931 12427
rect 10873 12387 10931 12393
rect 11422 12384 11428 12436
rect 11480 12424 11486 12436
rect 11701 12427 11759 12433
rect 11701 12424 11713 12427
rect 11480 12396 11713 12424
rect 11480 12384 11486 12396
rect 11701 12393 11713 12396
rect 11747 12393 11759 12427
rect 11701 12387 11759 12393
rect 11974 12384 11980 12436
rect 12032 12424 12038 12436
rect 12250 12424 12256 12436
rect 12032 12396 12256 12424
rect 12032 12384 12038 12396
rect 12250 12384 12256 12396
rect 12308 12384 12314 12436
rect 13078 12424 13084 12436
rect 12406 12396 13084 12424
rect 12406 12356 12434 12396
rect 13078 12384 13084 12396
rect 13136 12424 13142 12436
rect 15197 12427 15255 12433
rect 15197 12424 15209 12427
rect 13136 12396 15209 12424
rect 13136 12384 13142 12396
rect 15197 12393 15209 12396
rect 15243 12393 15255 12427
rect 15197 12387 15255 12393
rect 16114 12384 16120 12436
rect 16172 12424 16178 12436
rect 16390 12424 16396 12436
rect 16172 12396 16396 12424
rect 16172 12384 16178 12396
rect 16390 12384 16396 12396
rect 16448 12384 16454 12436
rect 16666 12384 16672 12436
rect 16724 12424 16730 12436
rect 17129 12427 17187 12433
rect 17129 12424 17141 12427
rect 16724 12396 17141 12424
rect 16724 12384 16730 12396
rect 17129 12393 17141 12396
rect 17175 12393 17187 12427
rect 17129 12387 17187 12393
rect 19150 12384 19156 12436
rect 19208 12424 19214 12436
rect 19797 12427 19855 12433
rect 19797 12424 19809 12427
rect 19208 12396 19809 12424
rect 19208 12384 19214 12396
rect 19797 12393 19809 12396
rect 19843 12393 19855 12427
rect 19797 12387 19855 12393
rect 23474 12384 23480 12436
rect 23532 12424 23538 12436
rect 25038 12424 25044 12436
rect 23532 12396 25044 12424
rect 23532 12384 23538 12396
rect 25038 12384 25044 12396
rect 25096 12384 25102 12436
rect 25406 12424 25412 12436
rect 25367 12396 25412 12424
rect 25406 12384 25412 12396
rect 25464 12384 25470 12436
rect 25498 12384 25504 12436
rect 25556 12424 25562 12436
rect 25556 12396 28028 12424
rect 25556 12384 25562 12396
rect 13722 12356 13728 12368
rect 11900 12328 12434 12356
rect 13683 12328 13728 12356
rect 10318 12288 10324 12300
rect 2148 12260 10324 12288
rect 2148 12229 2176 12260
rect 10318 12248 10324 12260
rect 10376 12248 10382 12300
rect 11900 12297 11928 12328
rect 13722 12316 13728 12328
rect 13780 12316 13786 12368
rect 18506 12356 18512 12368
rect 14936 12328 18512 12356
rect 14936 12300 14964 12328
rect 18506 12316 18512 12328
rect 18564 12316 18570 12368
rect 18690 12316 18696 12368
rect 18748 12356 18754 12368
rect 19168 12356 19196 12384
rect 18748 12328 19196 12356
rect 18748 12316 18754 12328
rect 19426 12316 19432 12368
rect 19484 12356 19490 12368
rect 21269 12359 21327 12365
rect 21269 12356 21281 12359
rect 19484 12328 21281 12356
rect 19484 12316 19490 12328
rect 21269 12325 21281 12328
rect 21315 12325 21327 12359
rect 21269 12319 21327 12325
rect 23014 12316 23020 12368
rect 23072 12356 23078 12368
rect 23382 12356 23388 12368
rect 23072 12328 23388 12356
rect 23072 12316 23078 12328
rect 23382 12316 23388 12328
rect 23440 12316 23446 12368
rect 24762 12316 24768 12368
rect 24820 12356 24826 12368
rect 26510 12356 26516 12368
rect 24820 12328 26516 12356
rect 24820 12316 24826 12328
rect 26510 12316 26516 12328
rect 26568 12316 26574 12368
rect 28000 12356 28028 12396
rect 28350 12384 28356 12436
rect 28408 12424 28414 12436
rect 28408 12396 32260 12424
rect 28408 12384 28414 12396
rect 29822 12356 29828 12368
rect 28000 12328 29828 12356
rect 29822 12316 29828 12328
rect 29880 12316 29886 12368
rect 32232 12356 32260 12396
rect 32306 12384 32312 12436
rect 32364 12424 32370 12436
rect 32401 12427 32459 12433
rect 32401 12424 32413 12427
rect 32364 12396 32413 12424
rect 32364 12384 32370 12396
rect 32401 12393 32413 12396
rect 32447 12393 32459 12427
rect 32401 12387 32459 12393
rect 32674 12384 32680 12436
rect 32732 12424 32738 12436
rect 32861 12427 32919 12433
rect 32861 12424 32873 12427
rect 32732 12396 32873 12424
rect 32732 12384 32738 12396
rect 32861 12393 32873 12396
rect 32907 12393 32919 12427
rect 32861 12387 32919 12393
rect 32950 12384 32956 12436
rect 33008 12424 33014 12436
rect 40770 12424 40776 12436
rect 33008 12396 40776 12424
rect 33008 12384 33014 12396
rect 40770 12384 40776 12396
rect 40828 12384 40834 12436
rect 42334 12424 42340 12436
rect 41892 12396 42340 12424
rect 41230 12356 41236 12368
rect 32232 12328 36032 12356
rect 11885 12291 11943 12297
rect 11885 12288 11897 12291
rect 10520 12260 11897 12288
rect 10520 12232 10548 12260
rect 11885 12257 11897 12260
rect 11931 12257 11943 12291
rect 11885 12251 11943 12257
rect 11977 12291 12035 12297
rect 11977 12257 11989 12291
rect 12023 12288 12035 12291
rect 13449 12291 13507 12297
rect 12023 12260 12434 12288
rect 12023 12257 12035 12260
rect 11977 12251 12035 12257
rect 2133 12223 2191 12229
rect 2133 12189 2145 12223
rect 2179 12189 2191 12223
rect 2133 12183 2191 12189
rect 2593 12223 2651 12229
rect 2593 12189 2605 12223
rect 2639 12220 2651 12223
rect 10502 12220 10508 12232
rect 2639 12192 2774 12220
rect 10415 12192 10508 12220
rect 2639 12189 2651 12192
rect 2593 12183 2651 12189
rect 2746 12084 2774 12192
rect 10502 12180 10508 12192
rect 10560 12180 10566 12232
rect 12066 12220 12072 12232
rect 12027 12192 12072 12220
rect 12066 12180 12072 12192
rect 12124 12180 12130 12232
rect 12161 12223 12219 12229
rect 12161 12189 12173 12223
rect 12207 12189 12219 12223
rect 12406 12220 12434 12260
rect 13449 12257 13461 12291
rect 13495 12288 13507 12291
rect 14553 12291 14611 12297
rect 14553 12288 14565 12291
rect 13495 12260 14565 12288
rect 13495 12257 13507 12260
rect 13449 12251 13507 12257
rect 14553 12257 14565 12260
rect 14599 12288 14611 12291
rect 14599 12260 14872 12288
rect 14599 12257 14611 12260
rect 14553 12251 14611 12257
rect 12526 12220 12532 12232
rect 12406 12192 12532 12220
rect 12161 12183 12219 12189
rect 10689 12155 10747 12161
rect 10689 12121 10701 12155
rect 10735 12152 10747 12155
rect 11054 12152 11060 12164
rect 10735 12124 11060 12152
rect 10735 12121 10747 12124
rect 10689 12115 10747 12121
rect 11054 12112 11060 12124
rect 11112 12112 11118 12164
rect 11882 12112 11888 12164
rect 11940 12152 11946 12164
rect 12176 12152 12204 12183
rect 12526 12180 12532 12192
rect 12584 12180 12590 12232
rect 13357 12223 13415 12229
rect 13357 12189 13369 12223
rect 13403 12220 13415 12223
rect 14844 12220 14872 12260
rect 14918 12248 14924 12300
rect 14976 12288 14982 12300
rect 14976 12260 15069 12288
rect 15304 12260 20392 12288
rect 14976 12248 14982 12260
rect 15304 12220 15332 12260
rect 13403 12192 14780 12220
rect 14844 12192 15332 12220
rect 13403 12189 13415 12192
rect 13357 12183 13415 12189
rect 11940 12124 12204 12152
rect 11940 12112 11946 12124
rect 14752 12096 14780 12192
rect 15378 12180 15384 12232
rect 15436 12220 15442 12232
rect 15654 12220 15660 12232
rect 15436 12192 15660 12220
rect 15436 12180 15442 12192
rect 15654 12180 15660 12192
rect 15712 12180 15718 12232
rect 15930 12220 15936 12232
rect 15891 12192 15936 12220
rect 15930 12180 15936 12192
rect 15988 12180 15994 12232
rect 18138 12220 18144 12232
rect 16040 12192 18144 12220
rect 15013 12155 15071 12161
rect 15013 12121 15025 12155
rect 15059 12152 15071 12155
rect 16040 12152 16068 12192
rect 18138 12180 18144 12192
rect 18196 12180 18202 12232
rect 18690 12220 18696 12232
rect 18651 12192 18696 12220
rect 18690 12180 18696 12192
rect 18748 12180 18754 12232
rect 18874 12220 18880 12232
rect 18835 12192 18880 12220
rect 18874 12180 18880 12192
rect 18932 12180 18938 12232
rect 19426 12220 19432 12232
rect 19387 12192 19432 12220
rect 19426 12180 19432 12192
rect 19484 12180 19490 12232
rect 19610 12220 19616 12232
rect 19571 12192 19616 12220
rect 19610 12180 19616 12192
rect 19668 12180 19674 12232
rect 20073 12223 20131 12229
rect 20073 12189 20085 12223
rect 20119 12189 20131 12223
rect 20073 12183 20131 12189
rect 15059 12124 16068 12152
rect 15059 12121 15071 12124
rect 15013 12115 15071 12121
rect 15672 12096 15700 12124
rect 16114 12112 16120 12164
rect 16172 12152 16178 12164
rect 19978 12152 19984 12164
rect 16172 12124 19984 12152
rect 16172 12112 16178 12124
rect 19978 12112 19984 12124
rect 20036 12112 20042 12164
rect 11238 12084 11244 12096
rect 2746 12056 11244 12084
rect 11238 12044 11244 12056
rect 11296 12044 11302 12096
rect 14734 12044 14740 12096
rect 14792 12084 14798 12096
rect 14829 12087 14887 12093
rect 14829 12084 14841 12087
rect 14792 12056 14841 12084
rect 14792 12044 14798 12056
rect 14829 12053 14841 12056
rect 14875 12053 14887 12087
rect 14829 12047 14887 12053
rect 15654 12044 15660 12096
rect 15712 12044 15718 12096
rect 17862 12044 17868 12096
rect 17920 12084 17926 12096
rect 18785 12087 18843 12093
rect 18785 12084 18797 12087
rect 17920 12056 18797 12084
rect 17920 12044 17926 12056
rect 18785 12053 18797 12056
rect 18831 12053 18843 12087
rect 18785 12047 18843 12053
rect 18966 12044 18972 12096
rect 19024 12084 19030 12096
rect 20088 12084 20116 12183
rect 20364 12152 20392 12260
rect 20530 12248 20536 12300
rect 20588 12288 20594 12300
rect 22741 12291 22799 12297
rect 22741 12288 22753 12291
rect 20588 12260 22753 12288
rect 20588 12248 20594 12260
rect 22741 12257 22753 12260
rect 22787 12288 22799 12291
rect 23290 12288 23296 12300
rect 22787 12260 23296 12288
rect 22787 12257 22799 12260
rect 22741 12251 22799 12257
rect 23290 12248 23296 12260
rect 23348 12248 23354 12300
rect 23661 12291 23719 12297
rect 23661 12257 23673 12291
rect 23707 12288 23719 12291
rect 24854 12288 24860 12300
rect 23707 12260 24860 12288
rect 23707 12257 23719 12260
rect 23661 12251 23719 12257
rect 24854 12248 24860 12260
rect 24912 12248 24918 12300
rect 24949 12291 25007 12297
rect 24949 12257 24961 12291
rect 24995 12288 25007 12291
rect 25222 12288 25228 12300
rect 24995 12260 25228 12288
rect 24995 12257 25007 12260
rect 24949 12251 25007 12257
rect 25222 12248 25228 12260
rect 25280 12248 25286 12300
rect 26053 12291 26111 12297
rect 26053 12257 26065 12291
rect 26099 12257 26111 12291
rect 26053 12251 26111 12257
rect 20898 12180 20904 12232
rect 20956 12220 20962 12232
rect 23198 12220 23204 12232
rect 20956 12192 23204 12220
rect 20956 12180 20962 12192
rect 23198 12180 23204 12192
rect 23256 12220 23262 12232
rect 23385 12223 23443 12229
rect 23385 12220 23397 12223
rect 23256 12192 23397 12220
rect 23256 12180 23262 12192
rect 23385 12189 23397 12192
rect 23431 12189 23443 12223
rect 23385 12183 23443 12189
rect 23750 12180 23756 12232
rect 23808 12220 23814 12232
rect 24578 12220 24584 12232
rect 23808 12192 24584 12220
rect 23808 12180 23814 12192
rect 24578 12180 24584 12192
rect 24636 12180 24642 12232
rect 24762 12220 24768 12232
rect 24723 12192 24768 12220
rect 24762 12180 24768 12192
rect 24820 12180 24826 12232
rect 25038 12180 25044 12232
rect 25096 12220 25102 12232
rect 25866 12220 25872 12232
rect 25096 12192 25872 12220
rect 25096 12180 25102 12192
rect 25866 12180 25872 12192
rect 25924 12180 25930 12232
rect 26068 12220 26096 12251
rect 26970 12248 26976 12300
rect 27028 12288 27034 12300
rect 27065 12291 27123 12297
rect 27065 12288 27077 12291
rect 27028 12260 27077 12288
rect 27028 12248 27034 12260
rect 27065 12257 27077 12260
rect 27111 12257 27123 12291
rect 27065 12251 27123 12257
rect 29086 12248 29092 12300
rect 29144 12288 29150 12300
rect 31478 12288 31484 12300
rect 29144 12260 31484 12288
rect 29144 12248 29150 12260
rect 28902 12220 28908 12232
rect 26068 12192 28908 12220
rect 28902 12180 28908 12192
rect 28960 12180 28966 12232
rect 30116 12229 30144 12260
rect 31036 12229 31064 12260
rect 31478 12248 31484 12260
rect 31536 12248 31542 12300
rect 31846 12288 31852 12300
rect 31772 12260 31852 12288
rect 30101 12223 30159 12229
rect 30101 12189 30113 12223
rect 30147 12189 30159 12223
rect 30101 12183 30159 12189
rect 30377 12223 30435 12229
rect 30377 12189 30389 12223
rect 30423 12189 30435 12223
rect 30377 12183 30435 12189
rect 31021 12223 31079 12229
rect 31021 12189 31033 12223
rect 31067 12189 31079 12223
rect 31294 12220 31300 12232
rect 31255 12192 31300 12220
rect 31021 12183 31079 12189
rect 25406 12152 25412 12164
rect 20364 12124 25412 12152
rect 25406 12112 25412 12124
rect 25464 12112 25470 12164
rect 26786 12112 26792 12164
rect 26844 12152 26850 12164
rect 27310 12155 27368 12161
rect 27310 12152 27322 12155
rect 26844 12124 27322 12152
rect 26844 12112 26850 12124
rect 27310 12121 27322 12124
rect 27356 12121 27368 12155
rect 27310 12115 27368 12121
rect 29178 12112 29184 12164
rect 29236 12152 29242 12164
rect 30285 12155 30343 12161
rect 30285 12152 30297 12155
rect 29236 12124 30297 12152
rect 29236 12112 29242 12124
rect 30285 12121 30297 12124
rect 30331 12121 30343 12155
rect 30392 12152 30420 12183
rect 31294 12180 31300 12192
rect 31352 12180 31358 12232
rect 31772 12229 31800 12260
rect 31846 12248 31852 12260
rect 31904 12248 31910 12300
rect 32490 12248 32496 12300
rect 32548 12288 32554 12300
rect 32548 12260 32593 12288
rect 32548 12248 32554 12260
rect 35526 12248 35532 12300
rect 35584 12288 35590 12300
rect 36004 12288 36032 12328
rect 40328 12328 41236 12356
rect 36630 12288 36636 12300
rect 35584 12260 35664 12288
rect 36004 12260 36492 12288
rect 36591 12260 36636 12288
rect 35584 12248 35590 12260
rect 31757 12223 31815 12229
rect 31757 12189 31769 12223
rect 31803 12189 31815 12223
rect 31938 12220 31944 12232
rect 31899 12192 31944 12220
rect 31757 12183 31815 12189
rect 31938 12180 31944 12192
rect 31996 12180 32002 12232
rect 32582 12220 32588 12232
rect 32232 12192 32588 12220
rect 30466 12152 30472 12164
rect 30379 12124 30472 12152
rect 30285 12115 30343 12121
rect 30466 12112 30472 12124
rect 30524 12152 30530 12164
rect 31849 12155 31907 12161
rect 31849 12152 31861 12155
rect 30524 12124 31861 12152
rect 30524 12112 30530 12124
rect 31849 12121 31861 12124
rect 31895 12121 31907 12155
rect 31849 12115 31907 12121
rect 20898 12084 20904 12096
rect 19024 12056 20904 12084
rect 19024 12044 19030 12056
rect 20898 12044 20904 12056
rect 20956 12044 20962 12096
rect 23014 12084 23020 12096
rect 22975 12056 23020 12084
rect 23014 12044 23020 12056
rect 23072 12044 23078 12096
rect 23290 12044 23296 12096
rect 23348 12084 23354 12096
rect 23477 12087 23535 12093
rect 23477 12084 23489 12087
rect 23348 12056 23489 12084
rect 23348 12044 23354 12056
rect 23477 12053 23489 12056
rect 23523 12084 23535 12087
rect 24302 12084 24308 12096
rect 23523 12056 24308 12084
rect 23523 12053 23535 12056
rect 23477 12047 23535 12053
rect 24302 12044 24308 12056
rect 24360 12044 24366 12096
rect 24854 12044 24860 12096
rect 24912 12084 24918 12096
rect 25498 12084 25504 12096
rect 24912 12056 25504 12084
rect 24912 12044 24918 12056
rect 25498 12044 25504 12056
rect 25556 12044 25562 12096
rect 25777 12087 25835 12093
rect 25777 12053 25789 12087
rect 25823 12084 25835 12087
rect 26878 12084 26884 12096
rect 25823 12056 26884 12084
rect 25823 12053 25835 12056
rect 25777 12047 25835 12053
rect 26878 12044 26884 12056
rect 26936 12044 26942 12096
rect 28442 12044 28448 12096
rect 28500 12084 28506 12096
rect 29914 12084 29920 12096
rect 28500 12056 28545 12084
rect 29875 12056 29920 12084
rect 28500 12044 28506 12056
rect 29914 12044 29920 12056
rect 29972 12044 29978 12096
rect 30834 12084 30840 12096
rect 30795 12056 30840 12084
rect 30834 12044 30840 12056
rect 30892 12044 30898 12096
rect 31202 12084 31208 12096
rect 31163 12056 31208 12084
rect 31202 12044 31208 12056
rect 31260 12044 31266 12096
rect 31386 12044 31392 12096
rect 31444 12084 31450 12096
rect 32232 12084 32260 12192
rect 32582 12180 32588 12192
rect 32640 12220 32646 12232
rect 32677 12223 32735 12229
rect 32677 12220 32689 12223
rect 32640 12192 32689 12220
rect 32640 12180 32646 12192
rect 32677 12189 32689 12192
rect 32723 12189 32735 12223
rect 32677 12183 32735 12189
rect 32950 12180 32956 12232
rect 33008 12220 33014 12232
rect 34238 12220 34244 12232
rect 33008 12192 34244 12220
rect 33008 12180 33014 12192
rect 34238 12180 34244 12192
rect 34296 12180 34302 12232
rect 35342 12220 35348 12232
rect 35303 12192 35348 12220
rect 35342 12180 35348 12192
rect 35400 12180 35406 12232
rect 35636 12229 35664 12260
rect 35621 12223 35679 12229
rect 35621 12189 35633 12223
rect 35667 12189 35679 12223
rect 35621 12183 35679 12189
rect 35713 12223 35771 12229
rect 35713 12189 35725 12223
rect 35759 12220 35771 12223
rect 35802 12220 35808 12232
rect 35759 12192 35808 12220
rect 35759 12189 35771 12192
rect 35713 12183 35771 12189
rect 35802 12180 35808 12192
rect 35860 12180 35866 12232
rect 35894 12180 35900 12232
rect 35952 12220 35958 12232
rect 36357 12223 36415 12229
rect 36357 12220 36369 12223
rect 35952 12192 36369 12220
rect 35952 12180 35958 12192
rect 36357 12189 36369 12192
rect 36403 12189 36415 12223
rect 36464 12220 36492 12260
rect 36630 12248 36636 12260
rect 36688 12248 36694 12300
rect 40328 12288 40356 12328
rect 41230 12316 41236 12328
rect 41288 12316 41294 12368
rect 41892 12297 41920 12396
rect 42334 12384 42340 12396
rect 42392 12384 42398 12436
rect 44634 12356 44640 12368
rect 42168 12328 44640 12356
rect 38626 12260 40356 12288
rect 38626 12220 38654 12260
rect 40034 12220 40040 12232
rect 36464 12192 38654 12220
rect 39995 12192 40040 12220
rect 36357 12183 36415 12189
rect 40034 12180 40040 12192
rect 40092 12180 40098 12232
rect 40126 12180 40132 12232
rect 40184 12220 40190 12232
rect 40184 12192 40229 12220
rect 40184 12180 40190 12192
rect 32401 12155 32459 12161
rect 32401 12121 32413 12155
rect 32447 12121 32459 12155
rect 32401 12115 32459 12121
rect 31444 12056 32260 12084
rect 32416 12084 32444 12115
rect 33870 12112 33876 12164
rect 33928 12152 33934 12164
rect 35529 12155 35587 12161
rect 35529 12152 35541 12155
rect 33928 12124 35541 12152
rect 33928 12112 33934 12124
rect 35529 12121 35541 12124
rect 35575 12121 35587 12155
rect 38010 12152 38016 12164
rect 37971 12124 38016 12152
rect 35529 12115 35587 12121
rect 38010 12112 38016 12124
rect 38068 12112 38074 12164
rect 40328 12161 40356 12260
rect 41877 12291 41935 12297
rect 41877 12257 41889 12291
rect 41923 12257 41935 12291
rect 41877 12251 41935 12257
rect 40586 12229 40592 12232
rect 40543 12223 40592 12229
rect 40543 12189 40555 12223
rect 40589 12189 40592 12223
rect 40543 12183 40592 12189
rect 40586 12180 40592 12183
rect 40644 12180 40650 12232
rect 41230 12180 41236 12232
rect 41288 12220 41294 12232
rect 41785 12223 41843 12229
rect 41288 12192 41736 12220
rect 41288 12180 41294 12192
rect 40313 12155 40371 12161
rect 40313 12121 40325 12155
rect 40359 12121 40371 12155
rect 40313 12115 40371 12121
rect 40405 12155 40463 12161
rect 40405 12121 40417 12155
rect 40451 12121 40463 12155
rect 40405 12115 40463 12121
rect 41141 12155 41199 12161
rect 41141 12121 41153 12155
rect 41187 12152 41199 12155
rect 41414 12152 41420 12164
rect 41187 12124 41420 12152
rect 41187 12121 41199 12124
rect 41141 12115 41199 12121
rect 35897 12087 35955 12093
rect 35897 12084 35909 12087
rect 32416 12056 35909 12084
rect 31444 12044 31450 12056
rect 35897 12053 35909 12056
rect 35943 12053 35955 12087
rect 35897 12047 35955 12053
rect 37918 12044 37924 12096
rect 37976 12084 37982 12096
rect 40420 12084 40448 12115
rect 41414 12112 41420 12124
rect 41472 12112 41478 12164
rect 41708 12152 41736 12192
rect 41785 12189 41797 12223
rect 41831 12220 41843 12223
rect 42058 12220 42064 12232
rect 41831 12192 42064 12220
rect 41831 12189 41843 12192
rect 41785 12183 41843 12189
rect 42058 12180 42064 12192
rect 42116 12180 42122 12232
rect 42168 12229 42196 12328
rect 44634 12316 44640 12328
rect 44692 12316 44698 12368
rect 42153 12223 42211 12229
rect 42153 12189 42165 12223
rect 42199 12189 42211 12223
rect 42153 12183 42211 12189
rect 42337 12223 42395 12229
rect 42337 12189 42349 12223
rect 42383 12189 42395 12223
rect 57882 12220 57888 12232
rect 57843 12192 57888 12220
rect 42337 12183 42395 12189
rect 42242 12152 42248 12164
rect 41708 12124 42248 12152
rect 42242 12112 42248 12124
rect 42300 12112 42306 12164
rect 42352 12152 42380 12183
rect 57882 12180 57888 12192
rect 57940 12180 57946 12232
rect 43346 12152 43352 12164
rect 42352 12124 43352 12152
rect 43346 12112 43352 12124
rect 43404 12152 43410 12164
rect 43714 12152 43720 12164
rect 43404 12124 43720 12152
rect 43404 12112 43410 12124
rect 43714 12112 43720 12124
rect 43772 12112 43778 12164
rect 58158 12152 58164 12164
rect 58119 12124 58164 12152
rect 58158 12112 58164 12124
rect 58216 12112 58222 12164
rect 37976 12056 40448 12084
rect 40681 12087 40739 12093
rect 37976 12044 37982 12056
rect 40681 12053 40693 12087
rect 40727 12084 40739 12087
rect 43254 12084 43260 12096
rect 40727 12056 43260 12084
rect 40727 12053 40739 12056
rect 40681 12047 40739 12053
rect 43254 12044 43260 12056
rect 43312 12044 43318 12096
rect 1104 11994 58880 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 58880 11994
rect 1104 11920 58880 11942
rect 9490 11840 9496 11892
rect 9548 11880 9554 11892
rect 10597 11883 10655 11889
rect 10597 11880 10609 11883
rect 9548 11852 10609 11880
rect 9548 11840 9554 11852
rect 10597 11849 10609 11852
rect 10643 11849 10655 11883
rect 10597 11843 10655 11849
rect 13998 11840 14004 11892
rect 14056 11880 14062 11892
rect 14553 11883 14611 11889
rect 14553 11880 14565 11883
rect 14056 11852 14565 11880
rect 14056 11840 14062 11852
rect 14553 11849 14565 11852
rect 14599 11849 14611 11883
rect 14553 11843 14611 11849
rect 15013 11883 15071 11889
rect 15013 11849 15025 11883
rect 15059 11880 15071 11883
rect 15930 11880 15936 11892
rect 15059 11852 15936 11880
rect 15059 11849 15071 11852
rect 15013 11843 15071 11849
rect 15930 11840 15936 11852
rect 15988 11840 15994 11892
rect 17402 11880 17408 11892
rect 16040 11852 17408 11880
rect 1854 11812 1860 11824
rect 1815 11784 1860 11812
rect 1854 11772 1860 11784
rect 1912 11772 1918 11824
rect 11054 11812 11060 11824
rect 10704 11784 11060 11812
rect 1581 11747 1639 11753
rect 1581 11713 1593 11747
rect 1627 11744 1639 11747
rect 10502 11744 10508 11756
rect 1627 11716 2774 11744
rect 10463 11716 10508 11744
rect 1627 11713 1639 11716
rect 1581 11707 1639 11713
rect 2746 11676 2774 11716
rect 10502 11704 10508 11716
rect 10560 11704 10566 11756
rect 10704 11753 10732 11784
rect 11054 11772 11060 11784
rect 11112 11812 11118 11824
rect 12250 11812 12256 11824
rect 11112 11784 12256 11812
rect 11112 11772 11118 11784
rect 12250 11772 12256 11784
rect 12308 11772 12314 11824
rect 13173 11815 13231 11821
rect 13173 11781 13185 11815
rect 13219 11812 13231 11815
rect 13262 11812 13268 11824
rect 13219 11784 13268 11812
rect 13219 11781 13231 11784
rect 13173 11775 13231 11781
rect 13262 11772 13268 11784
rect 13320 11772 13326 11824
rect 13389 11815 13447 11821
rect 13389 11781 13401 11815
rect 13435 11812 13447 11815
rect 13630 11812 13636 11824
rect 13435 11784 13636 11812
rect 13435 11781 13447 11784
rect 13389 11775 13447 11781
rect 13630 11772 13636 11784
rect 13688 11772 13694 11824
rect 14936 11784 15542 11812
rect 14936 11756 14964 11784
rect 10689 11747 10747 11753
rect 10689 11713 10701 11747
rect 10735 11713 10747 11747
rect 11882 11744 11888 11756
rect 11843 11716 11888 11744
rect 10689 11707 10747 11713
rect 11882 11704 11888 11716
rect 11940 11704 11946 11756
rect 11977 11747 12035 11753
rect 11977 11713 11989 11747
rect 12023 11744 12035 11747
rect 12342 11744 12348 11756
rect 12023 11716 12348 11744
rect 12023 11713 12035 11716
rect 11977 11707 12035 11713
rect 12342 11704 12348 11716
rect 12400 11704 12406 11756
rect 14185 11747 14243 11753
rect 14185 11713 14197 11747
rect 14231 11744 14243 11747
rect 14918 11744 14924 11756
rect 14231 11716 14924 11744
rect 14231 11713 14243 11716
rect 14185 11707 14243 11713
rect 14918 11704 14924 11716
rect 14976 11704 14982 11756
rect 15197 11747 15255 11753
rect 15197 11742 15209 11747
rect 15120 11714 15209 11742
rect 11701 11679 11759 11685
rect 11701 11676 11713 11679
rect 2746 11648 11713 11676
rect 11701 11645 11713 11648
rect 11747 11645 11759 11679
rect 11701 11639 11759 11645
rect 12069 11679 12127 11685
rect 12069 11645 12081 11679
rect 12115 11645 12127 11679
rect 12069 11639 12127 11645
rect 11790 11568 11796 11620
rect 11848 11608 11854 11620
rect 12084 11608 12112 11639
rect 12158 11636 12164 11688
rect 12216 11676 12222 11688
rect 14277 11679 14335 11685
rect 12216 11648 12261 11676
rect 12216 11636 12222 11648
rect 14277 11645 14289 11679
rect 14323 11645 14335 11679
rect 14277 11639 14335 11645
rect 11848 11580 12112 11608
rect 14292 11608 14320 11639
rect 14826 11636 14832 11688
rect 14884 11676 14890 11688
rect 15120 11676 15148 11714
rect 15197 11713 15209 11714
rect 15243 11713 15255 11747
rect 15197 11707 15255 11713
rect 15372 11747 15430 11753
rect 15372 11713 15384 11747
rect 15418 11742 15430 11747
rect 15514 11742 15542 11784
rect 16040 11753 16068 11852
rect 17402 11840 17408 11852
rect 17460 11840 17466 11892
rect 18995 11883 19053 11889
rect 18995 11849 19007 11883
rect 19041 11880 19053 11883
rect 19426 11880 19432 11892
rect 19041 11852 19432 11880
rect 19041 11849 19053 11852
rect 18995 11843 19053 11849
rect 19426 11840 19432 11852
rect 19484 11840 19490 11892
rect 19886 11840 19892 11892
rect 19944 11880 19950 11892
rect 19981 11883 20039 11889
rect 19981 11880 19993 11883
rect 19944 11852 19993 11880
rect 19944 11840 19950 11852
rect 19981 11849 19993 11852
rect 20027 11849 20039 11883
rect 19981 11843 20039 11849
rect 20070 11840 20076 11892
rect 20128 11880 20134 11892
rect 20349 11883 20407 11889
rect 20349 11880 20361 11883
rect 20128 11852 20361 11880
rect 20128 11840 20134 11852
rect 20349 11849 20361 11852
rect 20395 11849 20407 11883
rect 20349 11843 20407 11849
rect 20441 11883 20499 11889
rect 20441 11849 20453 11883
rect 20487 11880 20499 11883
rect 20898 11880 20904 11892
rect 20487 11852 20904 11880
rect 20487 11849 20499 11852
rect 20441 11843 20499 11849
rect 20898 11840 20904 11852
rect 20956 11840 20962 11892
rect 22370 11880 22376 11892
rect 22331 11852 22376 11880
rect 22370 11840 22376 11852
rect 22428 11840 22434 11892
rect 22738 11840 22744 11892
rect 22796 11880 22802 11892
rect 23474 11880 23480 11892
rect 22796 11852 23480 11880
rect 22796 11840 22802 11852
rect 23474 11840 23480 11852
rect 23532 11840 23538 11892
rect 25222 11840 25228 11892
rect 25280 11840 25286 11892
rect 26605 11883 26663 11889
rect 26605 11849 26617 11883
rect 26651 11880 26663 11883
rect 26786 11880 26792 11892
rect 26651 11852 26792 11880
rect 26651 11849 26663 11852
rect 26605 11843 26663 11849
rect 26786 11840 26792 11852
rect 26844 11840 26850 11892
rect 29914 11840 29920 11892
rect 29972 11880 29978 11892
rect 29972 11852 36584 11880
rect 29972 11840 29978 11852
rect 17120 11815 17178 11821
rect 17120 11781 17132 11815
rect 17166 11812 17178 11815
rect 17770 11812 17776 11824
rect 17166 11784 17776 11812
rect 17166 11781 17178 11784
rect 17120 11775 17178 11781
rect 17770 11772 17776 11784
rect 17828 11772 17834 11824
rect 18785 11815 18843 11821
rect 18785 11781 18797 11815
rect 18831 11812 18843 11815
rect 18874 11812 18880 11824
rect 18831 11784 18880 11812
rect 18831 11781 18843 11784
rect 18785 11775 18843 11781
rect 18874 11772 18880 11784
rect 18932 11772 18938 11824
rect 21082 11812 21088 11824
rect 20640 11784 21088 11812
rect 15418 11714 15542 11742
rect 16025 11747 16083 11753
rect 15418 11713 15430 11714
rect 15372 11707 15430 11713
rect 16025 11713 16037 11747
rect 16071 11713 16083 11747
rect 16025 11707 16083 11713
rect 16209 11747 16267 11753
rect 16209 11713 16221 11747
rect 16255 11744 16267 11747
rect 16666 11744 16672 11756
rect 16255 11716 16672 11744
rect 16255 11713 16267 11716
rect 16209 11707 16267 11713
rect 16666 11704 16672 11716
rect 16724 11704 16730 11756
rect 16850 11744 16856 11756
rect 16811 11716 16856 11744
rect 16850 11704 16856 11716
rect 16908 11704 16914 11756
rect 17402 11704 17408 11756
rect 17460 11744 17466 11756
rect 19794 11744 19800 11756
rect 17460 11716 19800 11744
rect 17460 11704 17466 11716
rect 19794 11704 19800 11716
rect 19852 11704 19858 11756
rect 20530 11744 20536 11756
rect 19904 11716 20536 11744
rect 14884 11648 15148 11676
rect 14884 11636 14890 11648
rect 15286 11636 15292 11688
rect 15344 11676 15350 11688
rect 15474 11679 15532 11685
rect 15344 11648 15389 11676
rect 15344 11636 15350 11648
rect 15474 11645 15486 11679
rect 15520 11676 15532 11679
rect 15654 11676 15660 11688
rect 15520 11648 15660 11676
rect 15520 11645 15532 11648
rect 15474 11639 15532 11645
rect 15654 11636 15660 11648
rect 15712 11636 15718 11688
rect 18156 11648 19012 11676
rect 16117 11611 16175 11617
rect 16117 11608 16129 11611
rect 14292 11580 16129 11608
rect 11848 11568 11854 11580
rect 16117 11577 16129 11580
rect 16163 11577 16175 11611
rect 16117 11571 16175 11577
rect 10318 11500 10324 11552
rect 10376 11540 10382 11552
rect 13170 11540 13176 11552
rect 10376 11512 13176 11540
rect 10376 11500 10382 11512
rect 13170 11500 13176 11512
rect 13228 11500 13234 11552
rect 13354 11540 13360 11552
rect 13315 11512 13360 11540
rect 13354 11500 13360 11512
rect 13412 11500 13418 11552
rect 13541 11543 13599 11549
rect 13541 11509 13553 11543
rect 13587 11540 13599 11543
rect 15654 11540 15660 11552
rect 13587 11512 15660 11540
rect 13587 11509 13599 11512
rect 13541 11503 13599 11509
rect 15654 11500 15660 11512
rect 15712 11500 15718 11552
rect 16390 11500 16396 11552
rect 16448 11540 16454 11552
rect 18156 11540 18184 11648
rect 18233 11611 18291 11617
rect 18233 11577 18245 11611
rect 18279 11608 18291 11611
rect 18874 11608 18880 11620
rect 18279 11580 18880 11608
rect 18279 11577 18291 11580
rect 18233 11571 18291 11577
rect 18874 11568 18880 11580
rect 18932 11568 18938 11620
rect 18984 11608 19012 11648
rect 19150 11636 19156 11688
rect 19208 11676 19214 11688
rect 19904 11676 19932 11716
rect 20530 11704 20536 11716
rect 20588 11704 20594 11756
rect 20640 11685 20668 11784
rect 21082 11772 21088 11784
rect 21140 11772 21146 11824
rect 25240 11812 25268 11840
rect 23860 11784 25268 11812
rect 22189 11747 22247 11753
rect 22189 11713 22201 11747
rect 22235 11744 22247 11747
rect 23014 11744 23020 11756
rect 22235 11716 23020 11744
rect 22235 11713 22247 11716
rect 22189 11707 22247 11713
rect 23014 11704 23020 11716
rect 23072 11704 23078 11756
rect 23860 11753 23888 11784
rect 25406 11772 25412 11824
rect 25464 11812 25470 11824
rect 30282 11812 30288 11824
rect 25464 11784 30288 11812
rect 25464 11772 25470 11784
rect 30282 11772 30288 11784
rect 30340 11772 30346 11824
rect 30834 11772 30840 11824
rect 30892 11812 30898 11824
rect 32858 11812 32864 11824
rect 30892 11784 32864 11812
rect 30892 11772 30898 11784
rect 32858 11772 32864 11784
rect 32916 11772 32922 11824
rect 34146 11812 34152 11824
rect 33060 11784 34152 11812
rect 23845 11747 23903 11753
rect 23845 11713 23857 11747
rect 23891 11713 23903 11747
rect 23845 11707 23903 11713
rect 25041 11747 25099 11753
rect 25041 11713 25053 11747
rect 25087 11713 25099 11747
rect 25222 11744 25228 11756
rect 25183 11716 25228 11744
rect 25041 11707 25099 11713
rect 19208 11648 19932 11676
rect 20625 11679 20683 11685
rect 19208 11636 19214 11648
rect 20625 11645 20637 11679
rect 20671 11645 20683 11679
rect 20625 11639 20683 11645
rect 22005 11679 22063 11685
rect 22005 11645 22017 11679
rect 22051 11645 22063 11679
rect 22005 11639 22063 11645
rect 18984 11580 19196 11608
rect 16448 11512 18184 11540
rect 16448 11500 16454 11512
rect 18690 11500 18696 11552
rect 18748 11540 18754 11552
rect 19168 11549 19196 11580
rect 19242 11568 19248 11620
rect 19300 11608 19306 11620
rect 19702 11608 19708 11620
rect 19300 11580 19708 11608
rect 19300 11568 19306 11580
rect 19702 11568 19708 11580
rect 19760 11568 19766 11620
rect 20070 11568 20076 11620
rect 20128 11608 20134 11620
rect 20346 11608 20352 11620
rect 20128 11580 20352 11608
rect 20128 11568 20134 11580
rect 20346 11568 20352 11580
rect 20404 11568 20410 11620
rect 20806 11568 20812 11620
rect 20864 11608 20870 11620
rect 22020 11608 22048 11639
rect 22278 11636 22284 11688
rect 22336 11676 22342 11688
rect 24670 11676 24676 11688
rect 22336 11648 24676 11676
rect 22336 11636 22342 11648
rect 24670 11636 24676 11648
rect 24728 11636 24734 11688
rect 25056 11676 25084 11707
rect 25222 11704 25228 11716
rect 25280 11704 25286 11756
rect 25498 11744 25504 11756
rect 25332 11716 25504 11744
rect 25332 11676 25360 11716
rect 25498 11704 25504 11716
rect 25556 11704 25562 11756
rect 26234 11744 26240 11756
rect 26195 11716 26240 11744
rect 26234 11704 26240 11716
rect 26292 11704 26298 11756
rect 26418 11744 26424 11756
rect 26379 11716 26424 11744
rect 26418 11704 26424 11716
rect 26476 11704 26482 11756
rect 27525 11747 27583 11753
rect 27525 11744 27537 11747
rect 27356 11716 27537 11744
rect 27356 11688 27384 11716
rect 27525 11713 27537 11716
rect 27571 11713 27583 11747
rect 30466 11744 30472 11756
rect 30427 11716 30472 11744
rect 27525 11707 27583 11713
rect 30466 11704 30472 11716
rect 30524 11704 30530 11756
rect 30561 11747 30619 11753
rect 30561 11713 30573 11747
rect 30607 11744 30619 11747
rect 30926 11744 30932 11756
rect 30607 11716 30932 11744
rect 30607 11713 30619 11716
rect 30561 11707 30619 11713
rect 30926 11704 30932 11716
rect 30984 11744 30990 11756
rect 31113 11747 31171 11753
rect 31113 11744 31125 11747
rect 30984 11716 31125 11744
rect 30984 11704 30990 11716
rect 31113 11713 31125 11716
rect 31159 11713 31171 11747
rect 31113 11707 31171 11713
rect 31297 11747 31355 11753
rect 31297 11713 31309 11747
rect 31343 11744 31355 11747
rect 32306 11744 32312 11756
rect 31343 11716 32312 11744
rect 31343 11713 31355 11716
rect 31297 11707 31355 11713
rect 25056 11648 25360 11676
rect 25406 11636 25412 11688
rect 25464 11676 25470 11688
rect 25464 11648 25509 11676
rect 25464 11636 25470 11648
rect 25590 11636 25596 11688
rect 25648 11676 25654 11688
rect 25648 11648 25693 11676
rect 25648 11636 25654 11648
rect 27338 11636 27344 11688
rect 27396 11636 27402 11688
rect 27430 11636 27436 11688
rect 27488 11676 27494 11688
rect 27985 11679 28043 11685
rect 27985 11676 27997 11679
rect 27488 11648 27997 11676
rect 27488 11636 27494 11648
rect 27985 11645 27997 11648
rect 28031 11676 28043 11679
rect 31312 11676 31340 11707
rect 32306 11704 32312 11716
rect 32364 11704 32370 11756
rect 32953 11747 33011 11753
rect 32953 11713 32965 11747
rect 32999 11744 33011 11747
rect 33060 11744 33088 11784
rect 34146 11772 34152 11784
rect 34204 11772 34210 11824
rect 35894 11812 35900 11824
rect 34716 11784 35900 11812
rect 32999 11716 33088 11744
rect 32999 11713 33011 11716
rect 32953 11707 33011 11713
rect 33134 11704 33140 11756
rect 33192 11744 33198 11756
rect 33229 11747 33287 11753
rect 33229 11744 33241 11747
rect 33192 11716 33241 11744
rect 33192 11704 33198 11716
rect 33229 11713 33241 11716
rect 33275 11713 33287 11747
rect 33229 11707 33287 11713
rect 33962 11704 33968 11756
rect 34020 11744 34026 11756
rect 34716 11753 34744 11784
rect 35894 11772 35900 11784
rect 35952 11772 35958 11824
rect 36556 11812 36584 11852
rect 37182 11840 37188 11892
rect 37240 11880 37246 11892
rect 44174 11880 44180 11892
rect 37240 11852 44180 11880
rect 37240 11840 37246 11852
rect 39114 11812 39120 11824
rect 36556 11784 39120 11812
rect 39114 11772 39120 11784
rect 39172 11772 39178 11824
rect 40512 11821 40540 11852
rect 44174 11840 44180 11852
rect 44232 11840 44238 11892
rect 46290 11840 46296 11892
rect 46348 11880 46354 11892
rect 59078 11880 59084 11892
rect 46348 11852 59084 11880
rect 46348 11840 46354 11852
rect 59078 11840 59084 11852
rect 59136 11840 59142 11892
rect 40497 11815 40555 11821
rect 40497 11781 40509 11815
rect 40543 11781 40555 11815
rect 40497 11775 40555 11781
rect 40586 11772 40592 11824
rect 40644 11812 40650 11824
rect 42886 11812 42892 11824
rect 40644 11784 42892 11812
rect 40644 11772 40650 11784
rect 42886 11772 42892 11784
rect 42944 11772 42950 11824
rect 43990 11812 43996 11824
rect 43364 11784 43996 11812
rect 34701 11747 34759 11753
rect 34701 11744 34713 11747
rect 34020 11716 34713 11744
rect 34020 11704 34026 11716
rect 34701 11713 34713 11716
rect 34747 11713 34759 11747
rect 34701 11707 34759 11713
rect 34968 11747 35026 11753
rect 34968 11713 34980 11747
rect 35014 11744 35026 11747
rect 35342 11744 35348 11756
rect 35014 11716 35348 11744
rect 35014 11713 35026 11716
rect 34968 11707 35026 11713
rect 35342 11704 35348 11716
rect 35400 11704 35406 11756
rect 38746 11744 38752 11756
rect 38707 11716 38752 11744
rect 38746 11704 38752 11716
rect 38804 11704 38810 11756
rect 38930 11704 38936 11756
rect 38988 11744 38994 11756
rect 38988 11716 41368 11744
rect 38988 11704 38994 11716
rect 28031 11648 31340 11676
rect 28031 11645 28043 11648
rect 27985 11639 28043 11645
rect 31478 11636 31484 11688
rect 31536 11676 31542 11688
rect 31846 11676 31852 11688
rect 31536 11648 31852 11676
rect 31536 11636 31542 11648
rect 31846 11636 31852 11648
rect 31904 11636 31910 11688
rect 32766 11636 32772 11688
rect 32824 11676 32830 11688
rect 33413 11679 33471 11685
rect 32824 11648 32996 11676
rect 32824 11636 32830 11648
rect 23750 11608 23756 11620
rect 20864 11580 23756 11608
rect 20864 11568 20870 11580
rect 23750 11568 23756 11580
rect 23808 11568 23814 11620
rect 31202 11608 31208 11620
rect 23860 11580 31208 11608
rect 18969 11543 19027 11549
rect 18969 11540 18981 11543
rect 18748 11512 18981 11540
rect 18748 11500 18754 11512
rect 18969 11509 18981 11512
rect 19015 11509 19027 11543
rect 18969 11503 19027 11509
rect 19153 11543 19211 11549
rect 19153 11509 19165 11543
rect 19199 11509 19211 11543
rect 19153 11503 19211 11509
rect 19518 11500 19524 11552
rect 19576 11540 19582 11552
rect 23860 11540 23888 11580
rect 31202 11568 31208 11580
rect 31260 11568 31266 11620
rect 31938 11568 31944 11620
rect 31996 11608 32002 11620
rect 32398 11608 32404 11620
rect 31996 11580 32404 11608
rect 31996 11568 32002 11580
rect 32398 11568 32404 11580
rect 32456 11568 32462 11620
rect 32968 11608 32996 11648
rect 33413 11645 33425 11679
rect 33459 11645 33471 11679
rect 41230 11676 41236 11688
rect 33413 11639 33471 11645
rect 35820 11648 41236 11676
rect 33045 11611 33103 11617
rect 33045 11608 33057 11611
rect 32968 11580 33057 11608
rect 33045 11577 33057 11580
rect 33091 11577 33103 11611
rect 33045 11571 33103 11577
rect 33134 11568 33140 11620
rect 33192 11608 33198 11620
rect 33428 11608 33456 11639
rect 35820 11608 35848 11648
rect 41230 11636 41236 11648
rect 41288 11636 41294 11688
rect 41340 11676 41368 11716
rect 42058 11704 42064 11756
rect 42116 11744 42122 11756
rect 43070 11744 43076 11756
rect 42116 11716 43076 11744
rect 42116 11704 42122 11716
rect 43070 11704 43076 11716
rect 43128 11704 43134 11756
rect 43254 11744 43260 11756
rect 43215 11716 43260 11744
rect 43254 11704 43260 11716
rect 43312 11704 43318 11756
rect 43364 11753 43392 11784
rect 43990 11772 43996 11784
rect 44048 11772 44054 11824
rect 44266 11772 44272 11824
rect 44324 11812 44330 11824
rect 50706 11812 50712 11824
rect 44324 11784 50712 11812
rect 44324 11772 44330 11784
rect 50706 11772 50712 11784
rect 50764 11772 50770 11824
rect 43349 11747 43407 11753
rect 43349 11713 43361 11747
rect 43395 11713 43407 11747
rect 43349 11707 43407 11713
rect 43625 11747 43683 11753
rect 43625 11713 43637 11747
rect 43671 11744 43683 11747
rect 43671 11716 45140 11744
rect 43671 11713 43683 11716
rect 43625 11707 43683 11713
rect 41414 11676 41420 11688
rect 41340 11648 41420 11676
rect 41414 11636 41420 11648
rect 41472 11636 41478 11688
rect 41506 11636 41512 11688
rect 41564 11676 41570 11688
rect 42702 11676 42708 11688
rect 41564 11648 42708 11676
rect 41564 11636 41570 11648
rect 42702 11636 42708 11648
rect 42760 11636 42766 11688
rect 43714 11676 43720 11688
rect 43675 11648 43720 11676
rect 43714 11636 43720 11648
rect 43772 11636 43778 11688
rect 45112 11676 45140 11716
rect 45186 11704 45192 11756
rect 45244 11744 45250 11756
rect 45462 11744 45468 11756
rect 45244 11716 45468 11744
rect 45244 11704 45250 11716
rect 45462 11704 45468 11716
rect 45520 11704 45526 11756
rect 45554 11704 45560 11756
rect 45612 11704 45618 11756
rect 45732 11747 45790 11753
rect 45732 11713 45744 11747
rect 45778 11744 45790 11747
rect 46106 11744 46112 11756
rect 45778 11716 46112 11744
rect 45778 11713 45790 11716
rect 45732 11707 45790 11713
rect 46106 11704 46112 11716
rect 46164 11704 46170 11756
rect 57146 11744 57152 11756
rect 57107 11716 57152 11744
rect 57146 11704 57152 11716
rect 57204 11704 57210 11756
rect 45572 11676 45600 11704
rect 45112 11648 45600 11676
rect 33192 11580 33456 11608
rect 35636 11580 35848 11608
rect 33192 11568 33198 11580
rect 19576 11512 23888 11540
rect 23937 11543 23995 11549
rect 19576 11500 19582 11512
rect 23937 11509 23949 11543
rect 23983 11540 23995 11543
rect 24026 11540 24032 11552
rect 23983 11512 24032 11540
rect 23983 11509 23995 11512
rect 23937 11503 23995 11509
rect 24026 11500 24032 11512
rect 24084 11500 24090 11552
rect 24762 11500 24768 11552
rect 24820 11540 24826 11552
rect 26694 11540 26700 11552
rect 24820 11512 26700 11540
rect 24820 11500 24826 11512
rect 26694 11500 26700 11512
rect 26752 11500 26758 11552
rect 31113 11543 31171 11549
rect 31113 11509 31125 11543
rect 31159 11540 31171 11543
rect 31294 11540 31300 11552
rect 31159 11512 31300 11540
rect 31159 11509 31171 11512
rect 31113 11503 31171 11509
rect 31294 11500 31300 11512
rect 31352 11540 31358 11552
rect 32122 11540 32128 11552
rect 31352 11512 32128 11540
rect 31352 11500 31358 11512
rect 32122 11500 32128 11512
rect 32180 11500 32186 11552
rect 32214 11500 32220 11552
rect 32272 11540 32278 11552
rect 35636 11540 35664 11580
rect 38010 11568 38016 11620
rect 38068 11608 38074 11620
rect 57422 11608 57428 11620
rect 38068 11580 45508 11608
rect 38068 11568 38074 11580
rect 32272 11512 35664 11540
rect 32272 11500 32278 11512
rect 35802 11500 35808 11552
rect 35860 11540 35866 11552
rect 36081 11543 36139 11549
rect 36081 11540 36093 11543
rect 35860 11512 36093 11540
rect 35860 11500 35866 11512
rect 36081 11509 36093 11512
rect 36127 11509 36139 11543
rect 36081 11503 36139 11509
rect 39850 11500 39856 11552
rect 39908 11540 39914 11552
rect 42058 11540 42064 11552
rect 39908 11512 42064 11540
rect 39908 11500 39914 11512
rect 42058 11500 42064 11512
rect 42116 11500 42122 11552
rect 42702 11540 42708 11552
rect 42615 11512 42708 11540
rect 42702 11500 42708 11512
rect 42760 11540 42766 11552
rect 43162 11540 43168 11552
rect 42760 11512 43168 11540
rect 42760 11500 42766 11512
rect 43162 11500 43168 11512
rect 43220 11500 43226 11552
rect 45480 11540 45508 11580
rect 46400 11580 57428 11608
rect 46400 11540 46428 11580
rect 57422 11568 57428 11580
rect 57480 11568 57486 11620
rect 46842 11540 46848 11552
rect 45480 11512 46428 11540
rect 46803 11512 46848 11540
rect 46842 11500 46848 11512
rect 46900 11500 46906 11552
rect 48314 11500 48320 11552
rect 48372 11540 48378 11552
rect 57241 11543 57299 11549
rect 57241 11540 57253 11543
rect 48372 11512 57253 11540
rect 48372 11500 48378 11512
rect 57241 11509 57253 11512
rect 57287 11509 57299 11543
rect 57241 11503 57299 11509
rect 1104 11450 58880 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 58880 11450
rect 1104 11376 58880 11398
rect 11882 11336 11888 11348
rect 11164 11308 11888 11336
rect 1762 11200 1768 11212
rect 1723 11172 1768 11200
rect 1762 11160 1768 11172
rect 1820 11160 1826 11212
rect 11164 11209 11192 11308
rect 11882 11296 11888 11308
rect 11940 11296 11946 11348
rect 15197 11339 15255 11345
rect 15197 11305 15209 11339
rect 15243 11336 15255 11339
rect 16758 11336 16764 11348
rect 15243 11308 16764 11336
rect 15243 11305 15255 11308
rect 15197 11299 15255 11305
rect 16758 11296 16764 11308
rect 16816 11296 16822 11348
rect 18046 11336 18052 11348
rect 18007 11308 18052 11336
rect 18046 11296 18052 11308
rect 18104 11296 18110 11348
rect 19334 11296 19340 11348
rect 19392 11336 19398 11348
rect 20254 11336 20260 11348
rect 19392 11308 20260 11336
rect 19392 11296 19398 11308
rect 20254 11296 20260 11308
rect 20312 11296 20318 11348
rect 20346 11296 20352 11348
rect 20404 11336 20410 11348
rect 20993 11339 21051 11345
rect 20993 11336 21005 11339
rect 20404 11308 21005 11336
rect 20404 11296 20410 11308
rect 20993 11305 21005 11308
rect 21039 11305 21051 11339
rect 20993 11299 21051 11305
rect 21082 11296 21088 11348
rect 21140 11336 21146 11348
rect 24029 11339 24087 11345
rect 24029 11336 24041 11339
rect 21140 11308 24041 11336
rect 21140 11296 21146 11308
rect 24029 11305 24041 11308
rect 24075 11305 24087 11339
rect 25222 11336 25228 11348
rect 24029 11299 24087 11305
rect 24136 11308 25228 11336
rect 11256 11240 16896 11268
rect 11256 11209 11284 11240
rect 10965 11203 11023 11209
rect 10965 11200 10977 11203
rect 2746 11172 10977 11200
rect 1581 11135 1639 11141
rect 1581 11101 1593 11135
rect 1627 11132 1639 11135
rect 2746 11132 2774 11172
rect 10965 11169 10977 11172
rect 11011 11169 11023 11203
rect 10965 11163 11023 11169
rect 11149 11203 11207 11209
rect 11149 11169 11161 11203
rect 11195 11169 11207 11203
rect 11149 11163 11207 11169
rect 11241 11203 11299 11209
rect 11241 11169 11253 11203
rect 11287 11169 11299 11203
rect 11241 11163 11299 11169
rect 11333 11203 11391 11209
rect 11333 11169 11345 11203
rect 11379 11200 11391 11203
rect 11698 11200 11704 11212
rect 11379 11172 11704 11200
rect 11379 11169 11391 11172
rect 11333 11163 11391 11169
rect 11698 11160 11704 11172
rect 11756 11160 11762 11212
rect 13170 11200 13176 11212
rect 13131 11172 13176 11200
rect 13170 11160 13176 11172
rect 13228 11160 13234 11212
rect 14826 11200 14832 11212
rect 14787 11172 14832 11200
rect 14826 11160 14832 11172
rect 14884 11160 14890 11212
rect 16868 11200 16896 11240
rect 20622 11228 20628 11280
rect 20680 11268 20686 11280
rect 21100 11268 21128 11296
rect 20680 11240 21128 11268
rect 23109 11271 23167 11277
rect 20680 11228 20686 11240
rect 23109 11237 23121 11271
rect 23155 11237 23167 11271
rect 23109 11231 23167 11237
rect 17862 11200 17868 11212
rect 16868 11172 17080 11200
rect 17823 11172 17868 11200
rect 1627 11104 2774 11132
rect 8588 11104 11284 11132
rect 1627 11101 1639 11104
rect 1581 11095 1639 11101
rect 8588 11076 8616 11104
rect 2866 11024 2872 11076
rect 2924 11064 2930 11076
rect 8570 11064 8576 11076
rect 2924 11036 8576 11064
rect 2924 11024 2930 11036
rect 8570 11024 8576 11036
rect 8628 11024 8634 11076
rect 11256 11064 11284 11104
rect 11422 11092 11428 11144
rect 11480 11132 11486 11144
rect 12989 11135 13047 11141
rect 12989 11132 13001 11135
rect 11480 11104 11525 11132
rect 12406 11104 13001 11132
rect 11480 11092 11486 11104
rect 12406 11064 12434 11104
rect 12989 11101 13001 11104
rect 13035 11101 13047 11135
rect 15010 11132 15016 11144
rect 14971 11104 15016 11132
rect 12989 11095 13047 11101
rect 15010 11092 15016 11104
rect 15068 11092 15074 11144
rect 15933 11135 15991 11141
rect 15933 11101 15945 11135
rect 15979 11101 15991 11135
rect 16390 11132 16396 11144
rect 16351 11104 16396 11132
rect 15933 11095 15991 11101
rect 15948 11064 15976 11095
rect 16390 11092 16396 11104
rect 16448 11092 16454 11144
rect 16574 11132 16580 11144
rect 16535 11104 16580 11132
rect 16574 11092 16580 11104
rect 16632 11092 16638 11144
rect 16666 11092 16672 11144
rect 16724 11132 16730 11144
rect 16853 11135 16911 11141
rect 16853 11132 16865 11135
rect 16724 11104 16865 11132
rect 16724 11092 16730 11104
rect 16853 11101 16865 11104
rect 16899 11101 16911 11135
rect 17052 11132 17080 11172
rect 17862 11160 17868 11172
rect 17920 11160 17926 11212
rect 17954 11160 17960 11212
rect 18012 11200 18018 11212
rect 19518 11200 19524 11212
rect 18012 11172 19524 11200
rect 18012 11160 18018 11172
rect 19518 11160 19524 11172
rect 19576 11160 19582 11212
rect 23124 11200 23152 11231
rect 23842 11228 23848 11280
rect 23900 11268 23906 11280
rect 24136 11268 24164 11308
rect 25222 11296 25228 11308
rect 25280 11296 25286 11348
rect 26142 11336 26148 11348
rect 25976 11308 26148 11336
rect 23900 11240 24164 11268
rect 23900 11228 23906 11240
rect 24302 11228 24308 11280
rect 24360 11268 24366 11280
rect 24578 11268 24584 11280
rect 24360 11240 24584 11268
rect 24360 11228 24366 11240
rect 24578 11228 24584 11240
rect 24636 11268 24642 11280
rect 25682 11268 25688 11280
rect 24636 11240 25688 11268
rect 24636 11228 24642 11240
rect 25682 11228 25688 11240
rect 25740 11268 25746 11280
rect 25976 11268 26004 11308
rect 26142 11296 26148 11308
rect 26200 11296 26206 11348
rect 27798 11296 27804 11348
rect 27856 11336 27862 11348
rect 28261 11339 28319 11345
rect 28261 11336 28273 11339
rect 27856 11308 28273 11336
rect 27856 11296 27862 11308
rect 28261 11305 28273 11308
rect 28307 11305 28319 11339
rect 28261 11299 28319 11305
rect 28994 11296 29000 11348
rect 29052 11336 29058 11348
rect 30466 11336 30472 11348
rect 29052 11308 30472 11336
rect 29052 11296 29058 11308
rect 30466 11296 30472 11308
rect 30524 11296 30530 11348
rect 35342 11336 35348 11348
rect 35303 11308 35348 11336
rect 35342 11296 35348 11308
rect 35400 11296 35406 11348
rect 36538 11296 36544 11348
rect 36596 11336 36602 11348
rect 36596 11308 40632 11336
rect 36596 11296 36602 11308
rect 25740 11240 26004 11268
rect 25740 11228 25746 11240
rect 26050 11228 26056 11280
rect 26108 11268 26114 11280
rect 29730 11268 29736 11280
rect 26108 11240 29736 11268
rect 26108 11228 26114 11240
rect 29730 11228 29736 11240
rect 29788 11228 29794 11280
rect 29822 11228 29828 11280
rect 29880 11268 29886 11280
rect 31389 11271 31447 11277
rect 29880 11240 30880 11268
rect 29880 11228 29886 11240
rect 30282 11200 30288 11212
rect 23124 11172 30288 11200
rect 30282 11160 30288 11172
rect 30340 11160 30346 11212
rect 30742 11200 30748 11212
rect 30703 11172 30748 11200
rect 30742 11160 30748 11172
rect 30800 11160 30806 11212
rect 30852 11200 30880 11240
rect 31389 11237 31401 11271
rect 31435 11268 31447 11271
rect 32398 11268 32404 11280
rect 31435 11240 32404 11268
rect 31435 11237 31447 11240
rect 31389 11231 31447 11237
rect 32398 11228 32404 11240
rect 32456 11228 32462 11280
rect 36078 11228 36084 11280
rect 36136 11268 36142 11280
rect 39850 11268 39856 11280
rect 36136 11240 39856 11268
rect 36136 11228 36142 11240
rect 39850 11228 39856 11240
rect 39908 11228 39914 11280
rect 30852 11172 31616 11200
rect 17052 11104 17264 11132
rect 16853 11095 16911 11101
rect 17126 11064 17132 11076
rect 10888 11036 11100 11064
rect 11256 11036 12434 11064
rect 15120 11036 15884 11064
rect 15948 11036 17132 11064
rect 1578 10956 1584 11008
rect 1636 10996 1642 11008
rect 10888 10996 10916 11036
rect 1636 10968 10916 10996
rect 11072 10996 11100 11036
rect 15120 10996 15148 11036
rect 15746 10996 15752 11008
rect 11072 10968 15148 10996
rect 15707 10968 15752 10996
rect 1636 10956 1642 10968
rect 15746 10956 15752 10968
rect 15804 10956 15810 11008
rect 15856 10996 15884 11036
rect 17126 11024 17132 11036
rect 17184 11024 17190 11076
rect 17236 11064 17264 11104
rect 17586 11092 17592 11144
rect 17644 11132 17650 11144
rect 17773 11135 17831 11141
rect 17773 11132 17785 11135
rect 17644 11104 17785 11132
rect 17644 11092 17650 11104
rect 17773 11101 17785 11104
rect 17819 11101 17831 11135
rect 17773 11095 17831 11101
rect 19426 11092 19432 11144
rect 19484 11132 19490 11144
rect 19886 11141 19892 11144
rect 19613 11135 19671 11141
rect 19613 11132 19625 11135
rect 19484 11104 19625 11132
rect 19484 11092 19490 11104
rect 19613 11101 19625 11104
rect 19659 11101 19671 11135
rect 19613 11095 19671 11101
rect 19869 11135 19892 11141
rect 19869 11101 19881 11135
rect 19869 11095 19892 11101
rect 19886 11092 19892 11095
rect 19944 11092 19950 11144
rect 23014 11132 23020 11144
rect 19996 11104 21220 11132
rect 22975 11104 23020 11132
rect 19996 11064 20024 11104
rect 21192 11064 21220 11104
rect 23014 11092 23020 11104
rect 23072 11092 23078 11144
rect 23106 11092 23112 11144
rect 23164 11132 23170 11144
rect 23201 11135 23259 11141
rect 23201 11132 23213 11135
rect 23164 11104 23213 11132
rect 23164 11092 23170 11104
rect 23201 11101 23213 11104
rect 23247 11101 23259 11135
rect 23750 11132 23756 11144
rect 23711 11104 23756 11132
rect 23201 11095 23259 11101
rect 23750 11092 23756 11104
rect 23808 11092 23814 11144
rect 23845 11135 23903 11141
rect 23845 11101 23857 11135
rect 23891 11132 23903 11135
rect 24486 11132 24492 11144
rect 23891 11104 24492 11132
rect 23891 11101 23903 11104
rect 23845 11095 23903 11101
rect 24486 11092 24492 11104
rect 24544 11092 24550 11144
rect 24581 11135 24639 11141
rect 24581 11101 24593 11135
rect 24627 11101 24639 11135
rect 24581 11095 24639 11101
rect 22738 11064 22744 11076
rect 17236 11036 20024 11064
rect 20916 11036 21128 11064
rect 21192 11036 22744 11064
rect 20916 10996 20944 11036
rect 15856 10968 20944 10996
rect 21100 10996 21128 11036
rect 22738 11024 22744 11036
rect 22796 11024 22802 11076
rect 23934 11024 23940 11076
rect 23992 11064 23998 11076
rect 24596 11064 24624 11095
rect 24670 11092 24676 11144
rect 24728 11132 24734 11144
rect 26050 11132 26056 11144
rect 24728 11104 26056 11132
rect 24728 11092 24734 11104
rect 26050 11092 26056 11104
rect 26108 11092 26114 11144
rect 26142 11092 26148 11144
rect 26200 11132 26206 11144
rect 28902 11132 28908 11144
rect 26200 11104 28908 11132
rect 26200 11092 26206 11104
rect 28902 11092 28908 11104
rect 28960 11092 28966 11144
rect 28994 11092 29000 11144
rect 29052 11132 29058 11144
rect 29917 11135 29975 11141
rect 29917 11132 29929 11135
rect 29052 11104 29929 11132
rect 29052 11092 29058 11104
rect 29917 11101 29929 11104
rect 29963 11101 29975 11135
rect 29917 11095 29975 11101
rect 31110 11092 31116 11144
rect 31168 11132 31174 11144
rect 31389 11135 31447 11141
rect 31389 11132 31401 11135
rect 31168 11104 31401 11132
rect 31168 11092 31174 11104
rect 31389 11101 31401 11104
rect 31435 11132 31447 11135
rect 31478 11132 31484 11144
rect 31435 11104 31484 11132
rect 31435 11101 31447 11104
rect 31389 11095 31447 11101
rect 31478 11092 31484 11104
rect 31536 11092 31542 11144
rect 31588 11141 31616 11172
rect 31846 11160 31852 11212
rect 31904 11200 31910 11212
rect 32490 11200 32496 11212
rect 31904 11172 32496 11200
rect 31904 11160 31910 11172
rect 32490 11160 32496 11172
rect 32548 11160 32554 11212
rect 35802 11200 35808 11212
rect 33612 11172 35808 11200
rect 31573 11135 31631 11141
rect 31573 11101 31585 11135
rect 31619 11101 31631 11135
rect 31573 11095 31631 11101
rect 31665 11135 31723 11141
rect 31665 11101 31677 11135
rect 31711 11132 31723 11135
rect 31864 11132 31892 11160
rect 32122 11132 32128 11144
rect 31711 11104 31892 11132
rect 32083 11104 32128 11132
rect 31711 11101 31723 11104
rect 31665 11095 31723 11101
rect 32122 11092 32128 11104
rect 32180 11092 32186 11144
rect 32217 11135 32275 11141
rect 32217 11101 32229 11135
rect 32263 11132 32275 11135
rect 32306 11132 32312 11144
rect 32263 11104 32312 11132
rect 32263 11101 32275 11104
rect 32217 11095 32275 11101
rect 32306 11092 32312 11104
rect 32364 11092 32370 11144
rect 23992 11036 24624 11064
rect 25409 11067 25467 11073
rect 23992 11024 23998 11036
rect 25409 11033 25421 11067
rect 25455 11064 25467 11067
rect 25682 11064 25688 11076
rect 25455 11036 25688 11064
rect 25455 11033 25467 11036
rect 25409 11027 25467 11033
rect 25682 11024 25688 11036
rect 25740 11024 25746 11076
rect 27706 11024 27712 11076
rect 27764 11064 27770 11076
rect 33612 11064 33640 11172
rect 35802 11160 35808 11172
rect 35860 11160 35866 11212
rect 35986 11160 35992 11212
rect 36044 11200 36050 11212
rect 38930 11200 38936 11212
rect 36044 11172 36089 11200
rect 36188 11172 38936 11200
rect 36044 11160 36050 11172
rect 33778 11132 33784 11144
rect 33739 11104 33784 11132
rect 33778 11092 33784 11104
rect 33836 11092 33842 11144
rect 34054 11132 34060 11144
rect 34015 11104 34060 11132
rect 34054 11092 34060 11104
rect 34112 11092 34118 11144
rect 34149 11135 34207 11141
rect 34149 11101 34161 11135
rect 34195 11132 34207 11135
rect 34422 11132 34428 11144
rect 34195 11104 34428 11132
rect 34195 11101 34207 11104
rect 34149 11095 34207 11101
rect 34422 11092 34428 11104
rect 34480 11092 34486 11144
rect 35710 11132 35716 11144
rect 35671 11104 35716 11132
rect 35710 11092 35716 11104
rect 35768 11092 35774 11144
rect 27764 11036 33640 11064
rect 27764 11024 27770 11036
rect 33870 11024 33876 11076
rect 33928 11064 33934 11076
rect 33965 11067 34023 11073
rect 33965 11064 33977 11067
rect 33928 11036 33977 11064
rect 33928 11024 33934 11036
rect 33965 11033 33977 11036
rect 34011 11033 34023 11067
rect 36188 11064 36216 11172
rect 38930 11160 38936 11172
rect 38988 11160 38994 11212
rect 40604 11200 40632 11308
rect 41322 11296 41328 11348
rect 41380 11336 41386 11348
rect 46106 11336 46112 11348
rect 41380 11308 45968 11336
rect 46067 11308 46112 11336
rect 41380 11296 41386 11308
rect 42058 11228 42064 11280
rect 42116 11268 42122 11280
rect 43070 11268 43076 11280
rect 42116 11240 42840 11268
rect 43031 11240 43076 11268
rect 42116 11228 42122 11240
rect 40604 11172 40724 11200
rect 38378 11092 38384 11144
rect 38436 11132 38442 11144
rect 38473 11135 38531 11141
rect 38473 11132 38485 11135
rect 38436 11104 38485 11132
rect 38436 11092 38442 11104
rect 38473 11101 38485 11104
rect 38519 11101 38531 11135
rect 38473 11095 38531 11101
rect 39942 11092 39948 11144
rect 40000 11132 40006 11144
rect 40589 11135 40647 11141
rect 40589 11132 40601 11135
rect 40000 11104 40601 11132
rect 40000 11092 40006 11104
rect 40589 11101 40601 11104
rect 40635 11101 40647 11135
rect 40696 11132 40724 11172
rect 42242 11160 42248 11212
rect 42300 11200 42306 11212
rect 42300 11172 42748 11200
rect 42300 11160 42306 11172
rect 42426 11132 42432 11144
rect 40696 11104 42288 11132
rect 42387 11104 42432 11132
rect 40589 11095 40647 11101
rect 33965 11027 34023 11033
rect 34072 11036 36216 11064
rect 34072 11008 34100 11036
rect 36354 11024 36360 11076
rect 36412 11064 36418 11076
rect 37090 11064 37096 11076
rect 36412 11036 37096 11064
rect 36412 11024 36418 11036
rect 37090 11024 37096 11036
rect 37148 11064 37154 11076
rect 38289 11067 38347 11073
rect 38289 11064 38301 11067
rect 37148 11036 38301 11064
rect 37148 11024 37154 11036
rect 38289 11033 38301 11036
rect 38335 11033 38347 11067
rect 38289 11027 38347 11033
rect 38654 11024 38660 11076
rect 38712 11064 38718 11076
rect 38841 11067 38899 11073
rect 38841 11064 38853 11067
rect 38712 11036 38853 11064
rect 38712 11024 38718 11036
rect 38841 11033 38853 11036
rect 38887 11033 38899 11067
rect 38841 11027 38899 11033
rect 40856 11067 40914 11073
rect 40856 11033 40868 11067
rect 40902 11064 40914 11067
rect 41138 11064 41144 11076
rect 40902 11036 41144 11064
rect 40902 11033 40914 11036
rect 40856 11027 40914 11033
rect 41138 11024 41144 11036
rect 41196 11024 41202 11076
rect 42260 11064 42288 11104
rect 42426 11092 42432 11104
rect 42484 11092 42490 11144
rect 42610 11141 42616 11144
rect 42577 11135 42616 11141
rect 42577 11101 42589 11135
rect 42577 11095 42616 11101
rect 42610 11092 42616 11095
rect 42668 11092 42674 11144
rect 42720 11141 42748 11172
rect 42812 11141 42840 11240
rect 43070 11228 43076 11240
rect 43128 11228 43134 11280
rect 45940 11268 45968 11308
rect 46106 11296 46112 11308
rect 46164 11296 46170 11348
rect 46216 11308 51074 11336
rect 46216 11268 46244 11308
rect 44192 11240 45232 11268
rect 45940 11240 46244 11268
rect 42705 11135 42763 11141
rect 42705 11101 42717 11135
rect 42751 11101 42763 11135
rect 42705 11095 42763 11101
rect 42797 11135 42855 11141
rect 42797 11101 42809 11135
rect 42843 11101 42855 11135
rect 42797 11095 42855 11101
rect 42886 11092 42892 11144
rect 42944 11141 42950 11144
rect 44192 11141 44220 11240
rect 45204 11200 45232 11240
rect 46566 11228 46572 11280
rect 46624 11268 46630 11280
rect 51046 11268 51074 11308
rect 56137 11271 56195 11277
rect 46624 11240 46704 11268
rect 51046 11240 55214 11268
rect 46624 11228 46630 11240
rect 46676 11209 46704 11240
rect 46661 11203 46719 11209
rect 45204 11172 46612 11200
rect 42944 11132 42952 11141
rect 44177 11135 44235 11141
rect 42944 11104 42989 11132
rect 42944 11095 42952 11104
rect 44177 11101 44189 11135
rect 44223 11101 44235 11135
rect 44450 11132 44456 11144
rect 44363 11104 44456 11132
rect 44177 11095 44235 11101
rect 42944 11092 42950 11095
rect 44450 11092 44456 11104
rect 44508 11132 44514 11144
rect 45094 11132 45100 11144
rect 44508 11104 45100 11132
rect 44508 11092 44514 11104
rect 45094 11092 45100 11104
rect 45152 11092 45158 11144
rect 46290 11092 46296 11144
rect 46348 11132 46354 11144
rect 46477 11135 46535 11141
rect 46477 11132 46489 11135
rect 46348 11104 46489 11132
rect 46348 11092 46354 11104
rect 46477 11101 46489 11104
rect 46523 11101 46535 11135
rect 46584 11132 46612 11172
rect 46661 11169 46673 11203
rect 46707 11169 46719 11203
rect 46661 11163 46719 11169
rect 46750 11132 46756 11144
rect 46584 11104 46756 11132
rect 46477 11095 46535 11101
rect 46750 11092 46756 11104
rect 46808 11092 46814 11144
rect 55186 11132 55214 11240
rect 56137 11237 56149 11271
rect 56183 11237 56195 11271
rect 56137 11231 56195 11237
rect 56152 11200 56180 11231
rect 57882 11228 57888 11280
rect 57940 11268 57946 11280
rect 58253 11271 58311 11277
rect 58253 11268 58265 11271
rect 57940 11240 58265 11268
rect 57940 11228 57946 11240
rect 58253 11237 58265 11240
rect 58299 11237 58311 11271
rect 58253 11231 58311 11237
rect 56152 11172 57008 11200
rect 56413 11135 56471 11141
rect 56413 11132 56425 11135
rect 55186 11104 56425 11132
rect 56413 11101 56425 11104
rect 56459 11101 56471 11135
rect 56870 11132 56876 11144
rect 56831 11104 56876 11132
rect 56413 11095 56471 11101
rect 56870 11092 56876 11104
rect 56928 11092 56934 11144
rect 56980 11132 57008 11172
rect 57129 11135 57187 11141
rect 57129 11132 57141 11135
rect 56980 11104 57141 11132
rect 57129 11101 57141 11104
rect 57175 11101 57187 11135
rect 57129 11095 57187 11101
rect 46569 11067 46627 11073
rect 46569 11064 46581 11067
rect 42260 11036 46581 11064
rect 46569 11033 46581 11036
rect 46615 11064 46627 11067
rect 46842 11064 46848 11076
rect 46615 11036 46848 11064
rect 46615 11033 46627 11036
rect 46569 11027 46627 11033
rect 46842 11024 46848 11036
rect 46900 11024 46906 11076
rect 56134 11064 56140 11076
rect 56095 11036 56140 11064
rect 56134 11024 56140 11036
rect 56192 11024 56198 11076
rect 56321 11067 56379 11073
rect 56321 11033 56333 11067
rect 56367 11064 56379 11067
rect 56962 11064 56968 11076
rect 56367 11036 56968 11064
rect 56367 11033 56379 11036
rect 56321 11027 56379 11033
rect 56962 11024 56968 11036
rect 57020 11024 57026 11076
rect 24578 10996 24584 11008
rect 21100 10968 24584 10996
rect 24578 10956 24584 10968
rect 24636 10956 24642 11008
rect 24670 10956 24676 11008
rect 24728 10996 24734 11008
rect 31294 10996 31300 11008
rect 24728 10968 31300 10996
rect 24728 10956 24734 10968
rect 31294 10956 31300 10968
rect 31352 10956 31358 11008
rect 31478 10956 31484 11008
rect 31536 10996 31542 11008
rect 32766 10996 32772 11008
rect 31536 10968 32772 10996
rect 31536 10956 31542 10968
rect 32766 10956 32772 10968
rect 32824 10956 32830 11008
rect 34054 10956 34060 11008
rect 34112 10956 34118 11008
rect 34330 10996 34336 11008
rect 34291 10968 34336 10996
rect 34330 10956 34336 10968
rect 34388 10956 34394 11008
rect 36078 10956 36084 11008
rect 36136 10996 36142 11008
rect 40954 10996 40960 11008
rect 36136 10968 40960 10996
rect 36136 10956 36142 10968
rect 40954 10956 40960 10968
rect 41012 10956 41018 11008
rect 41969 10999 42027 11005
rect 41969 10965 41981 10999
rect 42015 10996 42027 10999
rect 42058 10996 42064 11008
rect 42015 10968 42064 10996
rect 42015 10965 42027 10968
rect 41969 10959 42027 10965
rect 42058 10956 42064 10968
rect 42116 10956 42122 11008
rect 1104 10906 58880 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 58880 10906
rect 1104 10832 58880 10854
rect 1670 10752 1676 10804
rect 1728 10792 1734 10804
rect 1728 10764 2774 10792
rect 1728 10752 1734 10764
rect 1854 10724 1860 10736
rect 1815 10696 1860 10724
rect 1854 10684 1860 10696
rect 1912 10684 1918 10736
rect 2746 10724 2774 10764
rect 7374 10752 7380 10804
rect 7432 10792 7438 10804
rect 9217 10795 9275 10801
rect 9217 10792 9229 10795
rect 7432 10764 9229 10792
rect 7432 10752 7438 10764
rect 9217 10761 9229 10764
rect 9263 10761 9275 10795
rect 12158 10792 12164 10804
rect 12119 10764 12164 10792
rect 9217 10755 9275 10761
rect 12158 10752 12164 10764
rect 12216 10752 12222 10804
rect 13357 10795 13415 10801
rect 13357 10792 13369 10795
rect 12406 10764 13369 10792
rect 12406 10724 12434 10764
rect 13357 10761 13369 10764
rect 13403 10761 13415 10795
rect 25038 10792 25044 10804
rect 13357 10755 13415 10761
rect 15580 10764 25044 10792
rect 2746 10696 12434 10724
rect 1578 10656 1584 10668
rect 1539 10628 1584 10656
rect 1578 10616 1584 10628
rect 1636 10616 1642 10668
rect 9401 10659 9459 10665
rect 9401 10625 9413 10659
rect 9447 10656 9459 10659
rect 12710 10656 12716 10668
rect 9447 10628 12716 10656
rect 9447 10625 9459 10628
rect 9401 10619 9459 10625
rect 12710 10616 12716 10628
rect 12768 10616 12774 10668
rect 12894 10656 12900 10668
rect 12855 10628 12900 10656
rect 12894 10616 12900 10628
rect 12952 10616 12958 10668
rect 13173 10659 13231 10665
rect 13173 10625 13185 10659
rect 13219 10656 13231 10659
rect 13354 10656 13360 10668
rect 13219 10628 13360 10656
rect 13219 10625 13231 10628
rect 13173 10619 13231 10625
rect 13354 10616 13360 10628
rect 13412 10656 13418 10668
rect 15286 10656 15292 10668
rect 13412 10628 15292 10656
rect 13412 10616 13418 10628
rect 15286 10616 15292 10628
rect 15344 10616 15350 10668
rect 8941 10591 8999 10597
rect 8941 10557 8953 10591
rect 8987 10588 8999 10591
rect 9490 10588 9496 10600
rect 8987 10560 9496 10588
rect 8987 10557 8999 10560
rect 8941 10551 8999 10557
rect 9490 10548 9496 10560
rect 9548 10548 9554 10600
rect 9585 10591 9643 10597
rect 9585 10557 9597 10591
rect 9631 10557 9643 10591
rect 9585 10551 9643 10557
rect 9600 10520 9628 10551
rect 9674 10548 9680 10600
rect 9732 10588 9738 10600
rect 11698 10588 11704 10600
rect 9732 10560 9777 10588
rect 9876 10560 11704 10588
rect 9732 10548 9738 10560
rect 9876 10520 9904 10560
rect 11698 10548 11704 10560
rect 11756 10548 11762 10600
rect 12250 10548 12256 10600
rect 12308 10588 12314 10600
rect 15580 10588 15608 10764
rect 25038 10752 25044 10764
rect 25096 10752 25102 10804
rect 25332 10764 25728 10792
rect 15838 10684 15844 10736
rect 15896 10684 15902 10736
rect 16206 10684 16212 10736
rect 16264 10724 16270 10736
rect 16482 10724 16488 10736
rect 16264 10696 16488 10724
rect 16264 10684 16270 10696
rect 16482 10684 16488 10696
rect 16540 10684 16546 10736
rect 17034 10724 17040 10736
rect 16995 10696 17040 10724
rect 17034 10684 17040 10696
rect 17092 10684 17098 10736
rect 17497 10727 17555 10733
rect 17497 10693 17509 10727
rect 17543 10724 17555 10727
rect 17954 10724 17960 10736
rect 17543 10696 17960 10724
rect 17543 10693 17555 10696
rect 17497 10687 17555 10693
rect 17954 10684 17960 10696
rect 18012 10684 18018 10736
rect 19950 10727 20008 10733
rect 19950 10724 19962 10727
rect 18524 10696 19962 10724
rect 15654 10616 15660 10668
rect 15712 10656 15718 10668
rect 15749 10659 15807 10665
rect 15749 10656 15761 10659
rect 15712 10628 15761 10656
rect 15712 10616 15718 10628
rect 15749 10625 15761 10628
rect 15795 10625 15807 10659
rect 15856 10656 15884 10684
rect 16117 10659 16175 10665
rect 16117 10656 16129 10659
rect 15856 10628 16129 10656
rect 15749 10619 15807 10625
rect 16117 10625 16129 10628
rect 16163 10625 16175 10659
rect 16117 10619 16175 10625
rect 17310 10616 17316 10668
rect 17368 10656 17374 10668
rect 17405 10659 17463 10665
rect 17405 10656 17417 10659
rect 17368 10628 17417 10656
rect 17368 10616 17374 10628
rect 17405 10625 17417 10628
rect 17451 10625 17463 10659
rect 17405 10619 17463 10625
rect 12308 10560 15608 10588
rect 15841 10591 15899 10597
rect 12308 10548 12314 10560
rect 15841 10557 15853 10591
rect 15887 10557 15899 10591
rect 16206 10588 16212 10600
rect 16167 10560 16212 10588
rect 15841 10551 15899 10557
rect 9600 10492 9904 10520
rect 11146 10480 11152 10532
rect 11204 10520 11210 10532
rect 11977 10523 12035 10529
rect 11977 10520 11989 10523
rect 11204 10492 11989 10520
rect 11204 10480 11210 10492
rect 11977 10489 11989 10492
rect 12023 10489 12035 10523
rect 11977 10483 12035 10489
rect 12989 10523 13047 10529
rect 12989 10489 13001 10523
rect 13035 10520 13047 10523
rect 13170 10520 13176 10532
rect 13035 10492 13176 10520
rect 13035 10489 13047 10492
rect 12989 10483 13047 10489
rect 13170 10480 13176 10492
rect 13228 10480 13234 10532
rect 15194 10520 15200 10532
rect 15155 10492 15200 10520
rect 15194 10480 15200 10492
rect 15252 10480 15258 10532
rect 12158 10412 12164 10464
rect 12216 10452 12222 10464
rect 15212 10452 15240 10480
rect 12216 10424 15240 10452
rect 15856 10452 15884 10551
rect 16206 10548 16212 10560
rect 16264 10548 16270 10600
rect 16482 10548 16488 10600
rect 16540 10588 16546 10600
rect 16945 10591 17003 10597
rect 16945 10588 16957 10591
rect 16540 10560 16957 10588
rect 16540 10548 16546 10560
rect 16945 10557 16957 10560
rect 16991 10557 17003 10591
rect 16945 10551 17003 10557
rect 17126 10548 17132 10600
rect 17184 10588 17190 10600
rect 17957 10591 18015 10597
rect 17957 10588 17969 10591
rect 17184 10560 17969 10588
rect 17184 10548 17190 10560
rect 17957 10557 17969 10560
rect 18003 10557 18015 10591
rect 17957 10551 18015 10557
rect 18524 10529 18552 10696
rect 19950 10693 19962 10696
rect 19996 10693 20008 10727
rect 19950 10687 20008 10693
rect 20622 10684 20628 10736
rect 20680 10724 20686 10736
rect 20680 10696 20760 10724
rect 20680 10684 20686 10696
rect 18877 10659 18935 10665
rect 18877 10625 18889 10659
rect 18923 10625 18935 10659
rect 20530 10656 20536 10668
rect 18877 10619 18935 10625
rect 19168 10628 20536 10656
rect 18509 10523 18567 10529
rect 18509 10489 18521 10523
rect 18555 10489 18567 10523
rect 18892 10520 18920 10619
rect 18966 10548 18972 10600
rect 19024 10588 19030 10600
rect 19168 10597 19196 10628
rect 20530 10616 20536 10628
rect 20588 10616 20594 10668
rect 19153 10591 19211 10597
rect 19024 10560 19069 10588
rect 19024 10548 19030 10560
rect 19153 10557 19165 10591
rect 19199 10557 19211 10591
rect 19153 10551 19211 10557
rect 19426 10548 19432 10600
rect 19484 10588 19490 10600
rect 19705 10591 19763 10597
rect 19705 10588 19717 10591
rect 19484 10560 19717 10588
rect 19484 10548 19490 10560
rect 19705 10557 19717 10560
rect 19751 10557 19763 10591
rect 20732 10588 20760 10696
rect 23382 10684 23388 10736
rect 23440 10724 23446 10736
rect 23845 10727 23903 10733
rect 23440 10696 23796 10724
rect 23440 10684 23446 10696
rect 23768 10656 23796 10696
rect 23845 10693 23857 10727
rect 23891 10724 23903 10727
rect 25332 10724 25360 10764
rect 23891 10696 25360 10724
rect 25700 10724 25728 10764
rect 26418 10752 26424 10804
rect 26476 10792 26482 10804
rect 27157 10795 27215 10801
rect 27157 10792 27169 10795
rect 26476 10764 27169 10792
rect 26476 10752 26482 10764
rect 27157 10761 27169 10764
rect 27203 10761 27215 10795
rect 27157 10755 27215 10761
rect 28442 10752 28448 10804
rect 28500 10792 28506 10804
rect 29086 10792 29092 10804
rect 28500 10764 29092 10792
rect 28500 10752 28506 10764
rect 29086 10752 29092 10764
rect 29144 10752 29150 10804
rect 30282 10752 30288 10804
rect 30340 10792 30346 10804
rect 31297 10795 31355 10801
rect 31297 10792 31309 10795
rect 30340 10764 31309 10792
rect 30340 10752 30346 10764
rect 31297 10761 31309 10764
rect 31343 10761 31355 10795
rect 31297 10755 31355 10761
rect 32122 10752 32128 10804
rect 32180 10792 32186 10804
rect 32180 10764 34928 10792
rect 32180 10752 32186 10764
rect 27614 10724 27620 10736
rect 25700 10696 27620 10724
rect 23891 10693 23903 10696
rect 23845 10687 23903 10693
rect 27614 10684 27620 10696
rect 27672 10684 27678 10736
rect 29822 10684 29828 10736
rect 29880 10724 29886 10736
rect 29880 10696 33456 10724
rect 29880 10684 29886 10696
rect 24184 10659 24242 10665
rect 24184 10656 24196 10659
rect 23768 10628 24196 10656
rect 24184 10625 24196 10628
rect 24230 10625 24242 10659
rect 24184 10619 24242 10625
rect 25501 10659 25559 10665
rect 25501 10625 25513 10659
rect 25547 10625 25559 10659
rect 25866 10656 25872 10668
rect 25827 10628 25872 10656
rect 25501 10619 25559 10625
rect 23474 10588 23480 10600
rect 20732 10560 23480 10588
rect 19705 10551 19763 10557
rect 23474 10548 23480 10560
rect 23532 10548 23538 10600
rect 19518 10520 19524 10532
rect 18892 10492 19524 10520
rect 18509 10483 18567 10489
rect 19518 10480 19524 10492
rect 19576 10480 19582 10532
rect 21910 10520 21916 10532
rect 21008 10492 21916 10520
rect 21008 10452 21036 10492
rect 21910 10480 21916 10492
rect 21968 10480 21974 10532
rect 24121 10523 24179 10529
rect 24121 10489 24133 10523
rect 24167 10520 24179 10523
rect 24946 10520 24952 10532
rect 24167 10492 24952 10520
rect 24167 10489 24179 10492
rect 24121 10483 24179 10489
rect 24946 10480 24952 10492
rect 25004 10480 25010 10532
rect 25314 10520 25320 10532
rect 25275 10492 25320 10520
rect 25314 10480 25320 10492
rect 25372 10480 25378 10532
rect 25516 10520 25544 10619
rect 25866 10616 25872 10628
rect 25924 10616 25930 10668
rect 27525 10659 27583 10665
rect 27525 10656 27537 10659
rect 27356 10628 27537 10656
rect 25958 10588 25964 10600
rect 25919 10560 25964 10588
rect 25958 10548 25964 10560
rect 26016 10548 26022 10600
rect 26050 10520 26056 10532
rect 25516 10492 26056 10520
rect 26050 10480 26056 10492
rect 26108 10520 26114 10532
rect 27246 10520 27252 10532
rect 26108 10492 27252 10520
rect 26108 10480 26114 10492
rect 27246 10480 27252 10492
rect 27304 10480 27310 10532
rect 15856 10424 21036 10452
rect 21085 10455 21143 10461
rect 12216 10412 12222 10424
rect 21085 10421 21097 10455
rect 21131 10452 21143 10455
rect 21174 10452 21180 10464
rect 21131 10424 21180 10452
rect 21131 10421 21143 10424
rect 21085 10415 21143 10421
rect 21174 10412 21180 10424
rect 21232 10412 21238 10464
rect 22094 10412 22100 10464
rect 22152 10452 22158 10464
rect 23658 10452 23664 10464
rect 22152 10424 23664 10452
rect 22152 10412 22158 10424
rect 23658 10412 23664 10424
rect 23716 10412 23722 10464
rect 24010 10455 24068 10461
rect 24010 10421 24022 10455
rect 24056 10452 24068 10455
rect 24302 10452 24308 10464
rect 24056 10424 24308 10452
rect 24056 10421 24068 10424
rect 24010 10415 24068 10421
rect 24302 10412 24308 10424
rect 24360 10412 24366 10464
rect 24486 10452 24492 10464
rect 24447 10424 24492 10452
rect 24486 10412 24492 10424
rect 24544 10412 24550 10464
rect 24670 10412 24676 10464
rect 24728 10452 24734 10464
rect 27356 10452 27384 10628
rect 27525 10625 27537 10628
rect 27571 10656 27583 10659
rect 28442 10656 28448 10668
rect 27571 10628 28448 10656
rect 27571 10625 27583 10628
rect 27525 10619 27583 10625
rect 28442 10616 28448 10628
rect 28500 10616 28506 10668
rect 28721 10659 28779 10665
rect 28721 10625 28733 10659
rect 28767 10656 28779 10659
rect 29914 10656 29920 10668
rect 28767 10628 29920 10656
rect 28767 10625 28779 10628
rect 28721 10619 28779 10625
rect 29914 10616 29920 10628
rect 29972 10616 29978 10668
rect 31018 10616 31024 10668
rect 31076 10656 31082 10668
rect 31238 10659 31296 10665
rect 31238 10656 31250 10659
rect 31076 10628 31250 10656
rect 31076 10616 31082 10628
rect 31238 10625 31250 10628
rect 31284 10625 31296 10659
rect 31238 10619 31296 10625
rect 31478 10616 31484 10668
rect 31536 10656 31542 10668
rect 33321 10659 33379 10665
rect 33321 10656 33333 10659
rect 31536 10628 33333 10656
rect 31536 10616 31542 10628
rect 33321 10625 33333 10628
rect 33367 10625 33379 10659
rect 33428 10656 33456 10696
rect 34330 10684 34336 10736
rect 34388 10724 34394 10736
rect 34793 10727 34851 10733
rect 34793 10724 34805 10727
rect 34388 10696 34805 10724
rect 34388 10684 34394 10696
rect 34793 10693 34805 10696
rect 34839 10693 34851 10727
rect 34900 10724 34928 10764
rect 34974 10752 34980 10804
rect 35032 10792 35038 10804
rect 39390 10792 39396 10804
rect 35032 10764 39396 10792
rect 35032 10752 35038 10764
rect 39390 10752 39396 10764
rect 39448 10752 39454 10804
rect 41138 10792 41144 10804
rect 41099 10764 41144 10792
rect 41138 10752 41144 10764
rect 41196 10752 41202 10804
rect 49418 10792 49424 10804
rect 41248 10764 49424 10792
rect 41248 10724 41276 10764
rect 49418 10752 49424 10764
rect 49476 10752 49482 10804
rect 54018 10792 54024 10804
rect 53208 10764 54024 10792
rect 42058 10724 42064 10736
rect 34900 10696 41276 10724
rect 41432 10696 42064 10724
rect 34793 10687 34851 10693
rect 35109 10659 35167 10665
rect 33428 10628 35011 10656
rect 33321 10619 33379 10625
rect 27617 10591 27675 10597
rect 27617 10557 27629 10591
rect 27663 10557 27675 10591
rect 27798 10588 27804 10600
rect 27759 10560 27804 10588
rect 27617 10551 27675 10557
rect 27632 10520 27660 10551
rect 27798 10548 27804 10560
rect 27856 10548 27862 10600
rect 28166 10548 28172 10600
rect 28224 10588 28230 10600
rect 28997 10591 29055 10597
rect 28997 10588 29009 10591
rect 28224 10560 29009 10588
rect 28224 10548 28230 10560
rect 28997 10557 29009 10560
rect 29043 10557 29055 10591
rect 28997 10551 29055 10557
rect 29086 10548 29092 10600
rect 29144 10588 29150 10600
rect 31665 10591 31723 10597
rect 31665 10588 31677 10591
rect 29144 10560 31677 10588
rect 29144 10548 29150 10560
rect 31665 10557 31677 10560
rect 31711 10557 31723 10591
rect 31665 10551 31723 10557
rect 31754 10548 31760 10600
rect 31812 10588 31818 10600
rect 31812 10560 31857 10588
rect 31812 10548 31818 10560
rect 32582 10548 32588 10600
rect 32640 10588 32646 10600
rect 33689 10591 33747 10597
rect 33689 10588 33701 10591
rect 32640 10560 33701 10588
rect 32640 10548 32646 10560
rect 33336 10532 33364 10560
rect 33689 10557 33701 10560
rect 33735 10557 33747 10591
rect 33689 10551 33747 10557
rect 34790 10548 34796 10600
rect 34848 10588 34854 10600
rect 34885 10591 34943 10597
rect 34885 10588 34897 10591
rect 34848 10560 34897 10588
rect 34848 10548 34854 10560
rect 34885 10557 34897 10560
rect 34931 10557 34943 10591
rect 34983 10588 35011 10628
rect 35109 10625 35121 10659
rect 35155 10656 35167 10659
rect 35250 10656 35256 10668
rect 35155 10628 35256 10656
rect 35155 10625 35167 10628
rect 35109 10619 35167 10625
rect 35250 10616 35256 10628
rect 35308 10616 35314 10668
rect 35526 10616 35532 10668
rect 35584 10656 35590 10668
rect 37461 10659 37519 10665
rect 37461 10656 37473 10659
rect 35584 10628 37473 10656
rect 35584 10616 35590 10628
rect 37461 10625 37473 10628
rect 37507 10625 37519 10659
rect 41432 10656 41460 10696
rect 42058 10684 42064 10696
rect 42116 10684 42122 10736
rect 42886 10684 42892 10736
rect 42944 10724 42950 10736
rect 53208 10724 53236 10764
rect 54018 10752 54024 10764
rect 54076 10752 54082 10804
rect 56962 10752 56968 10804
rect 57020 10792 57026 10804
rect 57241 10795 57299 10801
rect 57241 10792 57253 10795
rect 57020 10764 57253 10792
rect 57020 10752 57026 10764
rect 57241 10761 57253 10764
rect 57287 10761 57299 10795
rect 57241 10755 57299 10761
rect 53374 10724 53380 10736
rect 42944 10696 53236 10724
rect 53335 10696 53380 10724
rect 42944 10684 42950 10696
rect 37461 10619 37519 10625
rect 37568 10628 41460 10656
rect 37568 10588 37596 10628
rect 37734 10588 37740 10600
rect 34983 10560 37596 10588
rect 37695 10560 37740 10588
rect 34885 10551 34943 10557
rect 37734 10548 37740 10560
rect 37792 10548 37798 10600
rect 38010 10548 38016 10600
rect 38068 10588 38074 10600
rect 38654 10588 38660 10600
rect 38068 10560 38660 10588
rect 38068 10548 38074 10560
rect 38654 10548 38660 10560
rect 38712 10548 38718 10600
rect 38746 10548 38752 10600
rect 38804 10588 38810 10600
rect 39114 10588 39120 10600
rect 38804 10560 39120 10588
rect 38804 10548 38810 10560
rect 39114 10548 39120 10560
rect 39172 10548 39178 10600
rect 41432 10588 41460 10628
rect 41509 10659 41567 10665
rect 41509 10625 41521 10659
rect 41555 10656 41567 10659
rect 41966 10656 41972 10668
rect 41555 10628 41972 10656
rect 41555 10625 41567 10628
rect 41509 10619 41567 10625
rect 41966 10616 41972 10628
rect 42024 10616 42030 10668
rect 44174 10656 44180 10668
rect 44135 10628 44180 10656
rect 44174 10616 44180 10628
rect 44232 10656 44238 10668
rect 46842 10656 46848 10668
rect 44232 10628 46848 10656
rect 44232 10616 44238 10628
rect 46842 10616 46848 10628
rect 46900 10616 46906 10668
rect 53101 10659 53159 10665
rect 53101 10625 53113 10659
rect 53147 10625 53159 10659
rect 53208 10656 53236 10696
rect 53374 10684 53380 10696
rect 53432 10684 53438 10736
rect 53285 10659 53343 10665
rect 53285 10656 53297 10659
rect 53208 10628 53297 10656
rect 53101 10619 53159 10625
rect 53285 10625 53297 10628
rect 53331 10625 53343 10659
rect 53466 10656 53472 10668
rect 53427 10628 53472 10656
rect 53285 10619 53343 10625
rect 41601 10591 41659 10597
rect 41601 10588 41613 10591
rect 41432 10560 41613 10588
rect 41601 10557 41613 10560
rect 41647 10557 41659 10591
rect 41601 10551 41659 10557
rect 41785 10591 41843 10597
rect 41785 10557 41797 10591
rect 41831 10588 41843 10591
rect 46566 10588 46572 10600
rect 41831 10560 46572 10588
rect 41831 10557 41843 10560
rect 41785 10551 41843 10557
rect 46566 10548 46572 10560
rect 46624 10548 46630 10600
rect 53116 10588 53144 10619
rect 53466 10616 53472 10628
rect 53524 10656 53530 10668
rect 54294 10656 54300 10668
rect 53524 10628 54300 10656
rect 53524 10616 53530 10628
rect 54294 10616 54300 10628
rect 54352 10616 54358 10668
rect 57054 10616 57060 10668
rect 57112 10656 57118 10668
rect 57149 10659 57207 10665
rect 57149 10656 57161 10659
rect 57112 10628 57161 10656
rect 57112 10616 57118 10628
rect 57149 10625 57161 10628
rect 57195 10625 57207 10659
rect 57149 10619 57207 10625
rect 57333 10659 57391 10665
rect 57333 10625 57345 10659
rect 57379 10656 57391 10659
rect 57882 10656 57888 10668
rect 57379 10628 57888 10656
rect 57379 10625 57391 10628
rect 57333 10619 57391 10625
rect 57882 10616 57888 10628
rect 57940 10616 57946 10668
rect 54202 10588 54208 10600
rect 53116 10560 54208 10588
rect 54202 10548 54208 10560
rect 54260 10548 54266 10600
rect 28350 10520 28356 10532
rect 27632 10492 28356 10520
rect 28350 10480 28356 10492
rect 28408 10480 28414 10532
rect 31113 10523 31171 10529
rect 31113 10489 31125 10523
rect 31159 10520 31171 10523
rect 31159 10492 33272 10520
rect 31159 10489 31171 10492
rect 31113 10483 31171 10489
rect 24728 10424 27384 10452
rect 24728 10412 24734 10424
rect 27798 10412 27804 10464
rect 27856 10452 27862 10464
rect 29178 10452 29184 10464
rect 27856 10424 29184 10452
rect 27856 10412 27862 10424
rect 29178 10412 29184 10424
rect 29236 10412 29242 10464
rect 29730 10412 29736 10464
rect 29788 10452 29794 10464
rect 30282 10452 30288 10464
rect 29788 10424 30288 10452
rect 29788 10412 29794 10424
rect 30282 10412 30288 10424
rect 30340 10412 30346 10464
rect 33244 10452 33272 10492
rect 33318 10480 33324 10532
rect 33376 10480 33382 10532
rect 53653 10523 53711 10529
rect 53653 10520 53665 10523
rect 35176 10492 44956 10520
rect 34974 10452 34980 10464
rect 33244 10424 34980 10452
rect 34974 10412 34980 10424
rect 35032 10412 35038 10464
rect 35069 10455 35127 10461
rect 35069 10421 35081 10455
rect 35115 10452 35127 10455
rect 35176 10452 35204 10492
rect 35115 10424 35204 10452
rect 35253 10455 35311 10461
rect 35115 10421 35127 10424
rect 35069 10415 35127 10421
rect 35253 10421 35265 10455
rect 35299 10452 35311 10455
rect 35342 10452 35348 10464
rect 35299 10424 35348 10452
rect 35299 10421 35311 10424
rect 35253 10415 35311 10421
rect 35342 10412 35348 10424
rect 35400 10412 35406 10464
rect 38102 10412 38108 10464
rect 38160 10452 38166 10464
rect 44818 10452 44824 10464
rect 38160 10424 44824 10452
rect 38160 10412 38166 10424
rect 44818 10412 44824 10424
rect 44876 10412 44882 10464
rect 44928 10452 44956 10492
rect 45112 10492 53665 10520
rect 45112 10452 45140 10492
rect 53653 10489 53665 10492
rect 53699 10489 53711 10523
rect 53653 10483 53711 10489
rect 44928 10424 45140 10452
rect 45186 10412 45192 10464
rect 45244 10452 45250 10464
rect 45465 10455 45523 10461
rect 45465 10452 45477 10455
rect 45244 10424 45477 10452
rect 45244 10412 45250 10424
rect 45465 10421 45477 10424
rect 45511 10421 45523 10455
rect 45465 10415 45523 10421
rect 45646 10412 45652 10464
rect 45704 10452 45710 10464
rect 53466 10452 53472 10464
rect 45704 10424 53472 10452
rect 45704 10412 45710 10424
rect 53466 10412 53472 10424
rect 53524 10412 53530 10464
rect 1104 10362 58880 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 58880 10362
rect 1104 10288 58880 10310
rect 11422 10208 11428 10260
rect 11480 10248 11486 10260
rect 11517 10251 11575 10257
rect 11517 10248 11529 10251
rect 11480 10220 11529 10248
rect 11480 10208 11486 10220
rect 11517 10217 11529 10220
rect 11563 10217 11575 10251
rect 11517 10211 11575 10217
rect 12268 10220 13768 10248
rect 11330 10180 11336 10192
rect 11291 10152 11336 10180
rect 11330 10140 11336 10152
rect 11388 10140 11394 10192
rect 1762 10112 1768 10124
rect 1723 10084 1768 10112
rect 1762 10072 1768 10084
rect 1820 10072 1826 10124
rect 2590 10072 2596 10124
rect 2648 10112 2654 10124
rect 12268 10112 12296 10220
rect 12897 10183 12955 10189
rect 12897 10149 12909 10183
rect 12943 10180 12955 10183
rect 13170 10180 13176 10192
rect 12943 10152 13176 10180
rect 12943 10149 12955 10152
rect 12897 10143 12955 10149
rect 13170 10140 13176 10152
rect 13228 10140 13234 10192
rect 13740 10180 13768 10220
rect 13814 10208 13820 10260
rect 13872 10248 13878 10260
rect 13872 10220 19472 10248
rect 13872 10208 13878 10220
rect 16206 10180 16212 10192
rect 13740 10152 16212 10180
rect 16206 10140 16212 10152
rect 16264 10140 16270 10192
rect 17678 10140 17684 10192
rect 17736 10180 17742 10192
rect 17862 10180 17868 10192
rect 17736 10152 17868 10180
rect 17736 10140 17742 10152
rect 17862 10140 17868 10152
rect 17920 10140 17926 10192
rect 18141 10183 18199 10189
rect 18141 10149 18153 10183
rect 18187 10180 18199 10183
rect 19334 10180 19340 10192
rect 18187 10152 19340 10180
rect 18187 10149 18199 10152
rect 18141 10143 18199 10149
rect 19334 10140 19340 10152
rect 19392 10140 19398 10192
rect 19444 10180 19472 10220
rect 19518 10208 19524 10260
rect 19576 10248 19582 10260
rect 21082 10248 21088 10260
rect 19576 10220 21088 10248
rect 19576 10208 19582 10220
rect 21082 10208 21088 10220
rect 21140 10208 21146 10260
rect 23658 10208 23664 10260
rect 23716 10248 23722 10260
rect 24486 10248 24492 10260
rect 23716 10220 24492 10248
rect 23716 10208 23722 10220
rect 24486 10208 24492 10220
rect 24544 10208 24550 10260
rect 25130 10248 25136 10260
rect 24596 10220 25136 10248
rect 19794 10180 19800 10192
rect 19444 10152 19800 10180
rect 19794 10140 19800 10152
rect 19852 10140 19858 10192
rect 21634 10180 21640 10192
rect 21595 10152 21640 10180
rect 21634 10140 21640 10152
rect 21692 10140 21698 10192
rect 23474 10180 23480 10192
rect 23435 10152 23480 10180
rect 23474 10140 23480 10152
rect 23532 10140 23538 10192
rect 14921 10115 14979 10121
rect 2648 10084 12296 10112
rect 12406 10084 14872 10112
rect 2648 10072 2654 10084
rect 1581 10047 1639 10053
rect 1581 10013 1593 10047
rect 1627 10044 1639 10047
rect 12406 10044 12434 10084
rect 1627 10016 12434 10044
rect 12805 10047 12863 10053
rect 1627 10013 1639 10016
rect 1581 10007 1639 10013
rect 12805 10013 12817 10047
rect 12851 10013 12863 10047
rect 12805 10007 12863 10013
rect 13081 10047 13139 10053
rect 13081 10013 13093 10047
rect 13127 10044 13139 10047
rect 13446 10044 13452 10056
rect 13127 10016 13452 10044
rect 13127 10013 13139 10016
rect 13081 10007 13139 10013
rect 11057 9979 11115 9985
rect 11057 9945 11069 9979
rect 11103 9976 11115 9979
rect 11698 9976 11704 9988
rect 11103 9948 11704 9976
rect 11103 9945 11115 9948
rect 11057 9939 11115 9945
rect 11698 9936 11704 9948
rect 11756 9936 11762 9988
rect 12820 9976 12848 10007
rect 13446 10004 13452 10016
rect 13504 10004 13510 10056
rect 14369 10047 14427 10053
rect 14369 10013 14381 10047
rect 14415 10013 14427 10047
rect 14844 10044 14872 10084
rect 14921 10081 14933 10115
rect 14967 10112 14979 10115
rect 15102 10112 15108 10124
rect 14967 10084 15108 10112
rect 14967 10081 14979 10084
rect 14921 10075 14979 10081
rect 15102 10072 15108 10084
rect 15160 10072 15166 10124
rect 15286 10072 15292 10124
rect 15344 10112 15350 10124
rect 18601 10115 18659 10121
rect 15344 10084 16344 10112
rect 15344 10072 15350 10084
rect 15654 10044 15660 10056
rect 14844 10016 15660 10044
rect 14369 10007 14427 10013
rect 12894 9976 12900 9988
rect 12807 9948 12900 9976
rect 12894 9936 12900 9948
rect 12952 9976 12958 9988
rect 13354 9976 13360 9988
rect 12952 9948 13360 9976
rect 12952 9936 12958 9948
rect 13354 9936 13360 9948
rect 13412 9936 13418 9988
rect 14384 9976 14412 10007
rect 15654 10004 15660 10016
rect 15712 10004 15718 10056
rect 16316 10053 16344 10084
rect 18601 10081 18613 10115
rect 18647 10112 18659 10115
rect 18690 10112 18696 10124
rect 18647 10084 18696 10112
rect 18647 10081 18659 10084
rect 18601 10075 18659 10081
rect 18690 10072 18696 10084
rect 18748 10072 18754 10124
rect 18782 10072 18788 10124
rect 18840 10112 18846 10124
rect 18840 10084 18885 10112
rect 18840 10072 18846 10084
rect 21818 10072 21824 10124
rect 21876 10112 21882 10124
rect 22189 10115 22247 10121
rect 22189 10112 22201 10115
rect 21876 10084 22201 10112
rect 21876 10072 21882 10084
rect 22189 10081 22201 10084
rect 22235 10081 22247 10115
rect 22189 10075 22247 10081
rect 22278 10072 22284 10124
rect 22336 10112 22342 10124
rect 24596 10112 24624 10220
rect 25130 10208 25136 10220
rect 25188 10208 25194 10260
rect 26510 10248 26516 10260
rect 25240 10220 26516 10248
rect 24762 10180 24768 10192
rect 22336 10084 24624 10112
rect 24688 10152 24768 10180
rect 22336 10072 22342 10084
rect 15933 10047 15991 10053
rect 15933 10013 15945 10047
rect 15979 10013 15991 10047
rect 15933 10007 15991 10013
rect 16301 10047 16359 10053
rect 16301 10013 16313 10047
rect 16347 10044 16359 10047
rect 16482 10044 16488 10056
rect 16347 10016 16488 10044
rect 16347 10013 16359 10016
rect 16301 10007 16359 10013
rect 15286 9976 15292 9988
rect 14384 9948 15292 9976
rect 15286 9936 15292 9948
rect 15344 9936 15350 9988
rect 1946 9868 1952 9920
rect 2004 9908 2010 9920
rect 13265 9911 13323 9917
rect 13265 9908 13277 9911
rect 2004 9880 13277 9908
rect 2004 9868 2010 9880
rect 13265 9877 13277 9880
rect 13311 9877 13323 9911
rect 13265 9871 13323 9877
rect 14182 9868 14188 9920
rect 14240 9908 14246 9920
rect 15948 9908 15976 10007
rect 16482 10004 16488 10016
rect 16540 10004 16546 10056
rect 16666 10044 16672 10056
rect 16627 10016 16672 10044
rect 16666 10004 16672 10016
rect 16724 10004 16730 10056
rect 17313 10047 17371 10053
rect 17313 10013 17325 10047
rect 17359 10044 17371 10047
rect 17402 10044 17408 10056
rect 17359 10016 17408 10044
rect 17359 10013 17371 10016
rect 17313 10007 17371 10013
rect 17402 10004 17408 10016
rect 17460 10004 17466 10056
rect 18509 10047 18567 10053
rect 18509 10013 18521 10047
rect 18555 10044 18567 10047
rect 19150 10044 19156 10056
rect 18555 10016 19156 10044
rect 18555 10013 18567 10016
rect 18509 10007 18567 10013
rect 19150 10004 19156 10016
rect 19208 10004 19214 10056
rect 19426 10004 19432 10056
rect 19484 10044 19490 10056
rect 19797 10047 19855 10053
rect 19797 10044 19809 10047
rect 19484 10016 19809 10044
rect 19484 10004 19490 10016
rect 19797 10013 19809 10016
rect 19843 10013 19855 10047
rect 19797 10007 19855 10013
rect 20990 10004 20996 10056
rect 21048 10044 21054 10056
rect 22005 10047 22063 10053
rect 22005 10044 22017 10047
rect 21048 10016 22017 10044
rect 21048 10004 21054 10016
rect 22005 10013 22017 10016
rect 22051 10013 22063 10047
rect 24029 10047 24087 10053
rect 24029 10044 24041 10047
rect 22005 10007 22063 10013
rect 23032 10016 24041 10044
rect 16853 9979 16911 9985
rect 16853 9945 16865 9979
rect 16899 9976 16911 9979
rect 19610 9976 19616 9988
rect 16899 9948 19616 9976
rect 16899 9945 16911 9948
rect 16853 9939 16911 9945
rect 19610 9936 19616 9948
rect 19668 9936 19674 9988
rect 20064 9979 20122 9985
rect 20064 9945 20076 9979
rect 20110 9976 20122 9979
rect 21634 9976 21640 9988
rect 20110 9948 21640 9976
rect 20110 9945 20122 9948
rect 20064 9939 20122 9945
rect 21634 9936 21640 9948
rect 21692 9936 21698 9988
rect 21818 9936 21824 9988
rect 21876 9976 21882 9988
rect 23032 9976 23060 10016
rect 24029 10013 24041 10016
rect 24075 10013 24087 10047
rect 24578 10044 24584 10056
rect 24539 10016 24584 10044
rect 24029 10007 24087 10013
rect 24578 10004 24584 10016
rect 24636 10004 24642 10056
rect 23658 9976 23664 9988
rect 21876 9948 23060 9976
rect 23619 9948 23664 9976
rect 21876 9936 21882 9948
rect 23658 9936 23664 9948
rect 23716 9936 23722 9988
rect 24688 9976 24716 10152
rect 24762 10140 24768 10152
rect 24820 10140 24826 10192
rect 25240 10180 25268 10220
rect 26510 10208 26516 10220
rect 26568 10208 26574 10260
rect 28166 10248 28172 10260
rect 28127 10220 28172 10248
rect 28166 10208 28172 10220
rect 28224 10208 28230 10260
rect 31478 10248 31484 10260
rect 28276 10220 31484 10248
rect 24872 10152 25268 10180
rect 24872 10112 24900 10152
rect 25314 10140 25320 10192
rect 25372 10180 25378 10192
rect 28276 10180 28304 10220
rect 31478 10208 31484 10220
rect 31536 10208 31542 10260
rect 31941 10251 31999 10257
rect 31941 10217 31953 10251
rect 31987 10248 31999 10251
rect 32214 10248 32220 10260
rect 31987 10220 32220 10248
rect 31987 10217 31999 10220
rect 31941 10211 31999 10217
rect 32214 10208 32220 10220
rect 32272 10208 32278 10260
rect 34422 10208 34428 10260
rect 34480 10248 34486 10260
rect 35526 10248 35532 10260
rect 34480 10220 35532 10248
rect 34480 10208 34486 10220
rect 35526 10208 35532 10220
rect 35584 10208 35590 10260
rect 36906 10208 36912 10260
rect 36964 10248 36970 10260
rect 38746 10248 38752 10260
rect 36964 10220 38752 10248
rect 36964 10208 36970 10220
rect 38746 10208 38752 10220
rect 38804 10208 38810 10260
rect 45462 10208 45468 10260
rect 45520 10248 45526 10260
rect 48133 10251 48191 10257
rect 48133 10248 48145 10251
rect 45520 10220 48145 10248
rect 45520 10208 45526 10220
rect 48133 10217 48145 10220
rect 48179 10248 48191 10251
rect 48774 10248 48780 10260
rect 48179 10220 48780 10248
rect 48179 10217 48191 10220
rect 48133 10211 48191 10217
rect 48774 10208 48780 10220
rect 48832 10208 48838 10260
rect 25372 10152 28304 10180
rect 25372 10140 25378 10152
rect 28810 10140 28816 10192
rect 28868 10180 28874 10192
rect 30650 10180 30656 10192
rect 28868 10152 30656 10180
rect 28868 10140 28874 10152
rect 30650 10140 30656 10152
rect 30708 10140 30714 10192
rect 30742 10140 30748 10192
rect 30800 10140 30806 10192
rect 33870 10140 33876 10192
rect 33928 10140 33934 10192
rect 37734 10140 37740 10192
rect 37792 10180 37798 10192
rect 38608 10180 38614 10192
rect 37792 10152 38614 10180
rect 37792 10140 37798 10152
rect 38608 10140 38614 10152
rect 38666 10140 38672 10192
rect 44192 10152 44490 10180
rect 24783 10084 24900 10112
rect 24783 10053 24811 10084
rect 26234 10072 26240 10124
rect 26292 10112 26298 10124
rect 26878 10112 26884 10124
rect 26292 10084 26884 10112
rect 26292 10072 26298 10084
rect 26878 10072 26884 10084
rect 26936 10112 26942 10124
rect 27801 10115 27859 10121
rect 27801 10112 27813 10115
rect 26936 10084 27813 10112
rect 26936 10072 26942 10084
rect 27801 10081 27813 10084
rect 27847 10081 27859 10115
rect 30760 10112 30788 10140
rect 32030 10112 32036 10124
rect 27801 10075 27859 10081
rect 29932 10084 30788 10112
rect 31726 10084 32036 10112
rect 24768 10047 24826 10053
rect 24768 10013 24780 10047
rect 24814 10013 24826 10047
rect 25130 10044 25136 10056
rect 25091 10016 25136 10044
rect 24768 10007 24826 10013
rect 25130 10004 25136 10016
rect 25188 10004 25194 10056
rect 27246 10044 27252 10056
rect 27207 10016 27252 10044
rect 27246 10004 27252 10016
rect 27304 10004 27310 10056
rect 27982 10044 27988 10056
rect 27943 10016 27988 10044
rect 27982 10004 27988 10016
rect 28040 10004 28046 10056
rect 28810 10044 28816 10056
rect 28771 10016 28816 10044
rect 28810 10004 28816 10016
rect 28868 10004 28874 10056
rect 28902 10004 28908 10056
rect 28960 10044 28966 10056
rect 29932 10053 29960 10084
rect 29181 10047 29239 10053
rect 29181 10044 29193 10047
rect 28960 10016 29193 10044
rect 28960 10004 28966 10016
rect 29181 10013 29193 10016
rect 29227 10013 29239 10047
rect 29181 10007 29239 10013
rect 29917 10047 29975 10053
rect 29917 10013 29929 10047
rect 29963 10013 29975 10047
rect 29917 10007 29975 10013
rect 30006 10004 30012 10056
rect 30064 10044 30070 10056
rect 30190 10044 30196 10056
rect 30064 10016 30109 10044
rect 30151 10016 30196 10044
rect 30064 10004 30070 10016
rect 30190 10004 30196 10016
rect 30248 10004 30254 10056
rect 30285 10047 30343 10053
rect 30285 10013 30297 10047
rect 30331 10044 30343 10047
rect 30466 10044 30472 10056
rect 30331 10016 30472 10044
rect 30331 10013 30343 10016
rect 30285 10007 30343 10013
rect 30466 10004 30472 10016
rect 30524 10004 30530 10056
rect 30745 10047 30803 10053
rect 30745 10013 30757 10047
rect 30791 10044 30803 10047
rect 31726 10044 31754 10084
rect 32030 10072 32036 10084
rect 32088 10112 32094 10124
rect 32950 10112 32956 10124
rect 32088 10084 32956 10112
rect 32088 10072 32094 10084
rect 32950 10072 32956 10084
rect 33008 10072 33014 10124
rect 33888 10112 33916 10140
rect 33612 10084 33916 10112
rect 32122 10044 32128 10056
rect 30791 10016 31754 10044
rect 32083 10016 32128 10044
rect 30791 10013 30803 10016
rect 30745 10007 30803 10013
rect 32122 10004 32128 10016
rect 32180 10004 32186 10056
rect 32398 10044 32404 10056
rect 32359 10016 32404 10044
rect 32398 10004 32404 10016
rect 32456 10004 32462 10056
rect 33318 10044 33324 10056
rect 33279 10016 33324 10044
rect 33318 10004 33324 10016
rect 33376 10004 33382 10056
rect 33410 10004 33416 10056
rect 33468 10044 33474 10056
rect 33612 10053 33640 10084
rect 34238 10072 34244 10124
rect 34296 10112 34302 10124
rect 34790 10112 34796 10124
rect 34296 10084 34796 10112
rect 34296 10072 34302 10084
rect 34790 10072 34796 10084
rect 34848 10072 34854 10124
rect 35342 10072 35348 10124
rect 35400 10072 35406 10124
rect 36630 10072 36636 10124
rect 36688 10112 36694 10124
rect 36688 10084 37780 10112
rect 36688 10072 36694 10084
rect 33597 10047 33655 10053
rect 33468 10016 33513 10044
rect 33468 10004 33474 10016
rect 33597 10013 33609 10047
rect 33643 10013 33655 10047
rect 33827 10047 33885 10053
rect 33827 10044 33839 10047
rect 33597 10007 33655 10013
rect 33820 10013 33839 10044
rect 33873 10044 33885 10047
rect 34977 10047 35035 10053
rect 33873 10016 34928 10044
rect 33873 10013 33885 10016
rect 33820 10007 33885 10013
rect 24946 9976 24952 9988
rect 25004 9985 25010 9988
rect 25004 9979 25025 9985
rect 23768 9948 24716 9976
rect 24783 9948 24952 9976
rect 18966 9908 18972 9920
rect 14240 9880 18972 9908
rect 14240 9868 14246 9880
rect 18966 9868 18972 9880
rect 19024 9868 19030 9920
rect 20530 9868 20536 9920
rect 20588 9908 20594 9920
rect 23768 9917 23796 9948
rect 21177 9911 21235 9917
rect 21177 9908 21189 9911
rect 20588 9880 21189 9908
rect 20588 9868 20594 9880
rect 21177 9877 21189 9880
rect 21223 9908 21235 9911
rect 22097 9911 22155 9917
rect 22097 9908 22109 9911
rect 21223 9880 22109 9908
rect 21223 9877 21235 9880
rect 21177 9871 21235 9877
rect 22097 9877 22109 9880
rect 22143 9877 22155 9911
rect 22097 9871 22155 9877
rect 23753 9911 23811 9917
rect 23753 9877 23765 9911
rect 23799 9877 23811 9911
rect 23753 9871 23811 9877
rect 23845 9911 23903 9917
rect 23845 9877 23857 9911
rect 23891 9908 23903 9911
rect 24783 9908 24811 9948
rect 24946 9936 24952 9948
rect 25013 9945 25025 9979
rect 25590 9976 25596 9988
rect 25551 9948 25596 9976
rect 25004 9939 25025 9945
rect 25004 9936 25010 9939
rect 25590 9936 25596 9948
rect 25648 9936 25654 9988
rect 25774 9976 25780 9988
rect 25700 9948 25780 9976
rect 23891 9880 24811 9908
rect 24857 9911 24915 9917
rect 23891 9877 23903 9880
rect 23845 9871 23903 9877
rect 24857 9877 24869 9911
rect 24903 9908 24915 9911
rect 25700 9908 25728 9948
rect 25774 9936 25780 9948
rect 25832 9936 25838 9988
rect 27614 9936 27620 9988
rect 27672 9976 27678 9988
rect 28629 9979 28687 9985
rect 28629 9976 28641 9979
rect 27672 9948 28641 9976
rect 27672 9936 27678 9948
rect 28629 9945 28641 9948
rect 28675 9945 28687 9979
rect 29822 9976 29828 9988
rect 28629 9939 28687 9945
rect 28920 9948 29828 9976
rect 28920 9917 28948 9948
rect 29822 9936 29828 9948
rect 29880 9936 29886 9988
rect 30098 9936 30104 9988
rect 30156 9976 30162 9988
rect 31021 9979 31079 9985
rect 31021 9976 31033 9979
rect 30156 9948 31033 9976
rect 30156 9936 30162 9948
rect 31021 9945 31033 9948
rect 31067 9945 31079 9979
rect 31021 9939 31079 9945
rect 31110 9936 31116 9988
rect 31168 9976 31174 9988
rect 32309 9979 32367 9985
rect 32309 9976 32321 9979
rect 31168 9948 32321 9976
rect 31168 9936 31174 9948
rect 32309 9945 32321 9948
rect 32355 9945 32367 9979
rect 33686 9976 33692 9988
rect 33647 9948 33692 9976
rect 32309 9939 32367 9945
rect 33686 9936 33692 9948
rect 33744 9936 33750 9988
rect 24903 9880 25728 9908
rect 28905 9911 28963 9917
rect 24903 9877 24915 9880
rect 24857 9871 24915 9877
rect 28905 9877 28917 9911
rect 28951 9877 28963 9911
rect 28905 9871 28963 9877
rect 28997 9911 29055 9917
rect 28997 9877 29009 9911
rect 29043 9908 29055 9911
rect 29546 9908 29552 9920
rect 29043 9880 29552 9908
rect 29043 9877 29055 9880
rect 28997 9871 29055 9877
rect 29546 9868 29552 9880
rect 29604 9868 29610 9920
rect 29733 9911 29791 9917
rect 29733 9877 29745 9911
rect 29779 9908 29791 9911
rect 31202 9908 31208 9920
rect 29779 9880 31208 9908
rect 29779 9877 29791 9880
rect 29733 9871 29791 9877
rect 31202 9868 31208 9880
rect 31260 9868 31266 9920
rect 32214 9868 32220 9920
rect 32272 9908 32278 9920
rect 33820 9908 33848 10007
rect 34146 9976 34152 9988
rect 33980 9948 34152 9976
rect 33980 9917 34008 9948
rect 34146 9936 34152 9948
rect 34204 9936 34210 9988
rect 32272 9880 33848 9908
rect 33965 9911 34023 9917
rect 32272 9868 32278 9880
rect 33965 9877 33977 9911
rect 34011 9877 34023 9911
rect 34900 9908 34928 10016
rect 34977 10013 34989 10047
rect 35023 10044 35035 10047
rect 35360 10044 35388 10072
rect 35023 10016 35388 10044
rect 35023 10013 35035 10016
rect 34977 10007 35035 10013
rect 36906 10004 36912 10056
rect 36964 10044 36970 10056
rect 37093 10047 37151 10053
rect 37093 10044 37105 10047
rect 36964 10016 37105 10044
rect 36964 10004 36970 10016
rect 37093 10013 37105 10016
rect 37139 10013 37151 10047
rect 37366 10044 37372 10056
rect 37327 10016 37372 10044
rect 37093 10007 37151 10013
rect 37366 10004 37372 10016
rect 37424 10004 37430 10056
rect 37458 10004 37464 10056
rect 37516 10044 37522 10056
rect 37752 10044 37780 10084
rect 38120 10084 41092 10112
rect 38120 10053 38148 10084
rect 41064 10056 41092 10084
rect 41230 10072 41236 10124
rect 41288 10112 41294 10124
rect 44192 10112 44220 10152
rect 41288 10084 44220 10112
rect 41288 10072 41294 10084
rect 38105 10047 38163 10053
rect 37516 10016 37561 10044
rect 37752 10016 37872 10044
rect 37516 10004 37522 10016
rect 35158 9976 35164 9988
rect 35119 9948 35164 9976
rect 35158 9936 35164 9948
rect 35216 9936 35222 9988
rect 35342 9976 35348 9988
rect 35303 9948 35348 9976
rect 35342 9936 35348 9948
rect 35400 9936 35406 9988
rect 37277 9979 37335 9985
rect 37277 9945 37289 9979
rect 37323 9976 37335 9979
rect 37734 9976 37740 9988
rect 37323 9948 37740 9976
rect 37323 9945 37335 9948
rect 37277 9939 37335 9945
rect 37734 9936 37740 9948
rect 37792 9936 37798 9988
rect 37844 9976 37872 10016
rect 38105 10013 38117 10047
rect 38151 10013 38163 10047
rect 38378 10044 38384 10056
rect 38339 10016 38384 10044
rect 38105 10007 38163 10013
rect 38378 10004 38384 10016
rect 38436 10004 38442 10056
rect 38562 10053 38568 10056
rect 38519 10047 38568 10053
rect 38519 10013 38531 10047
rect 38565 10013 38568 10047
rect 38519 10007 38568 10013
rect 38562 10004 38568 10007
rect 38620 10004 38626 10056
rect 41046 10004 41052 10056
rect 41104 10004 41110 10056
rect 44082 10044 44088 10056
rect 44043 10016 44088 10044
rect 44082 10004 44088 10016
rect 44140 10004 44146 10056
rect 44462 10053 44490 10152
rect 44542 10140 44548 10192
rect 44600 10180 44606 10192
rect 44600 10152 51074 10180
rect 44600 10140 44606 10152
rect 44818 10072 44824 10124
rect 44876 10112 44882 10124
rect 45646 10112 45652 10124
rect 44876 10084 45652 10112
rect 44876 10072 44882 10084
rect 45646 10072 45652 10084
rect 45704 10072 45710 10124
rect 46658 10112 46664 10124
rect 45940 10084 46664 10112
rect 45940 10053 45968 10084
rect 46658 10072 46664 10084
rect 46716 10072 46722 10124
rect 44177 10047 44235 10053
rect 44177 10013 44189 10047
rect 44223 10013 44235 10047
rect 44177 10007 44235 10013
rect 44269 10047 44327 10053
rect 44269 10013 44281 10047
rect 44315 10041 44327 10047
rect 44447 10047 44505 10053
rect 44315 10013 44404 10041
rect 44269 10007 44327 10013
rect 38289 9979 38347 9985
rect 38289 9976 38301 9979
rect 37844 9948 38301 9976
rect 38289 9945 38301 9948
rect 38335 9945 38347 9979
rect 38289 9939 38347 9945
rect 39390 9936 39396 9988
rect 39448 9976 39454 9988
rect 44192 9976 44220 10007
rect 39448 9948 44220 9976
rect 44376 9976 44404 10013
rect 44447 10013 44459 10047
rect 44493 10013 44505 10047
rect 44447 10007 44505 10013
rect 45925 10047 45983 10053
rect 45925 10013 45937 10047
rect 45971 10013 45983 10047
rect 45925 10007 45983 10013
rect 46106 10004 46112 10056
rect 46164 10044 46170 10056
rect 46201 10047 46259 10053
rect 46201 10044 46213 10047
rect 46164 10016 46213 10044
rect 46164 10004 46170 10016
rect 46201 10013 46213 10016
rect 46247 10013 46259 10047
rect 46842 10044 46848 10056
rect 46803 10016 46848 10044
rect 46201 10007 46259 10013
rect 46842 10004 46848 10016
rect 46900 10004 46906 10056
rect 44376 9948 45784 9976
rect 39448 9936 39454 9948
rect 36170 9908 36176 9920
rect 34900 9880 36176 9908
rect 33965 9871 34023 9877
rect 36170 9868 36176 9880
rect 36228 9868 36234 9920
rect 37458 9868 37464 9920
rect 37516 9908 37522 9920
rect 37645 9911 37703 9917
rect 37645 9908 37657 9911
rect 37516 9880 37657 9908
rect 37516 9868 37522 9880
rect 37645 9877 37657 9880
rect 37691 9877 37703 9911
rect 37645 9871 37703 9877
rect 38562 9868 38568 9920
rect 38620 9908 38626 9920
rect 38657 9911 38715 9917
rect 38657 9908 38669 9911
rect 38620 9880 38669 9908
rect 38620 9868 38626 9880
rect 38657 9877 38669 9880
rect 38703 9877 38715 9911
rect 38657 9871 38715 9877
rect 40310 9868 40316 9920
rect 40368 9908 40374 9920
rect 40770 9908 40776 9920
rect 40368 9880 40776 9908
rect 40368 9868 40374 9880
rect 40770 9868 40776 9880
rect 40828 9868 40834 9920
rect 43809 9911 43867 9917
rect 43809 9877 43821 9911
rect 43855 9908 43867 9911
rect 45462 9908 45468 9920
rect 43855 9880 45468 9908
rect 43855 9877 43867 9880
rect 43809 9871 43867 9877
rect 45462 9868 45468 9880
rect 45520 9868 45526 9920
rect 45756 9917 45784 9948
rect 45741 9911 45799 9917
rect 45741 9877 45753 9911
rect 45787 9877 45799 9911
rect 45741 9871 45799 9877
rect 46109 9911 46167 9917
rect 46109 9877 46121 9911
rect 46155 9908 46167 9911
rect 46290 9908 46296 9920
rect 46155 9880 46296 9908
rect 46155 9877 46167 9880
rect 46109 9871 46167 9877
rect 46290 9868 46296 9880
rect 46348 9868 46354 9920
rect 51046 9908 51074 10152
rect 58158 10112 58164 10124
rect 58119 10084 58164 10112
rect 58158 10072 58164 10084
rect 58216 10072 58222 10124
rect 56502 10004 56508 10056
rect 56560 10044 56566 10056
rect 57885 10047 57943 10053
rect 57885 10044 57897 10047
rect 56560 10016 57897 10044
rect 56560 10004 56566 10016
rect 57885 10013 57897 10016
rect 57931 10013 57943 10047
rect 57885 10007 57943 10013
rect 57054 9976 57060 9988
rect 57015 9948 57060 9976
rect 57054 9936 57060 9948
rect 57112 9936 57118 9988
rect 51718 9908 51724 9920
rect 51046 9880 51724 9908
rect 51718 9868 51724 9880
rect 51776 9868 51782 9920
rect 57146 9908 57152 9920
rect 57107 9880 57152 9908
rect 57146 9868 57152 9880
rect 57204 9868 57210 9920
rect 1104 9818 58880 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 58880 9818
rect 1104 9744 58880 9766
rect 16390 9704 16396 9716
rect 15580 9676 16396 9704
rect 11238 9596 11244 9648
rect 11296 9636 11302 9648
rect 13538 9636 13544 9648
rect 11296 9608 13544 9636
rect 11296 9596 11302 9608
rect 13538 9596 13544 9608
rect 13596 9636 13602 9648
rect 15102 9636 15108 9648
rect 13596 9608 13676 9636
rect 13596 9596 13602 9608
rect 1578 9568 1584 9580
rect 1539 9540 1584 9568
rect 1578 9528 1584 9540
rect 1636 9528 1642 9580
rect 13354 9568 13360 9580
rect 13315 9540 13360 9568
rect 13354 9528 13360 9540
rect 13412 9528 13418 9580
rect 13446 9528 13452 9580
rect 13504 9568 13510 9580
rect 13648 9577 13676 9608
rect 13740 9608 15108 9636
rect 13740 9577 13768 9608
rect 15102 9596 15108 9608
rect 15160 9596 15166 9648
rect 15580 9580 15608 9676
rect 16390 9664 16396 9676
rect 16448 9704 16454 9716
rect 17402 9704 17408 9716
rect 16448 9676 17408 9704
rect 16448 9664 16454 9676
rect 17402 9664 17408 9676
rect 17460 9664 17466 9716
rect 18598 9664 18604 9716
rect 18656 9704 18662 9716
rect 18782 9704 18788 9716
rect 18656 9676 18788 9704
rect 18656 9664 18662 9676
rect 18782 9664 18788 9676
rect 18840 9664 18846 9716
rect 22005 9707 22063 9713
rect 22005 9673 22017 9707
rect 22051 9673 22063 9707
rect 22005 9667 22063 9673
rect 22373 9707 22431 9713
rect 22373 9673 22385 9707
rect 22419 9704 22431 9707
rect 22419 9676 22692 9704
rect 22419 9673 22431 9676
rect 22373 9667 22431 9673
rect 20064 9639 20122 9645
rect 16316 9608 18092 9636
rect 13633 9571 13691 9577
rect 13504 9540 13549 9568
rect 13504 9528 13510 9540
rect 13633 9537 13645 9571
rect 13679 9537 13691 9571
rect 13633 9531 13691 9537
rect 13725 9571 13783 9577
rect 13725 9537 13737 9571
rect 13771 9537 13783 9571
rect 14182 9568 14188 9580
rect 14143 9540 14188 9568
rect 13725 9531 13783 9537
rect 14182 9528 14188 9540
rect 14240 9528 14246 9580
rect 15289 9571 15347 9577
rect 15289 9568 15301 9571
rect 14844 9540 15301 9568
rect 1762 9500 1768 9512
rect 1723 9472 1768 9500
rect 1762 9460 1768 9472
rect 1820 9460 1826 9512
rect 8754 9500 8760 9512
rect 8715 9472 8760 9500
rect 8754 9460 8760 9472
rect 8812 9460 8818 9512
rect 9217 9503 9275 9509
rect 9217 9469 9229 9503
rect 9263 9500 9275 9503
rect 9674 9500 9680 9512
rect 9263 9472 9680 9500
rect 9263 9469 9275 9472
rect 9217 9463 9275 9469
rect 9674 9460 9680 9472
rect 9732 9460 9738 9512
rect 13262 9460 13268 9512
rect 13320 9500 13326 9512
rect 14274 9500 14280 9512
rect 13320 9472 14280 9500
rect 13320 9460 13326 9472
rect 14274 9460 14280 9472
rect 14332 9460 14338 9512
rect 7190 9392 7196 9444
rect 7248 9432 7254 9444
rect 9033 9435 9091 9441
rect 9033 9432 9045 9435
rect 7248 9404 9045 9432
rect 7248 9392 7254 9404
rect 9033 9401 9045 9404
rect 9079 9401 9091 9435
rect 9033 9395 9091 9401
rect 12710 9324 12716 9376
rect 12768 9364 12774 9376
rect 13170 9364 13176 9376
rect 12768 9336 13176 9364
rect 12768 9324 12774 9336
rect 13170 9324 13176 9336
rect 13228 9324 13234 9376
rect 13630 9324 13636 9376
rect 13688 9364 13694 9376
rect 14844 9364 14872 9540
rect 15289 9537 15301 9540
rect 15335 9537 15347 9571
rect 15562 9568 15568 9580
rect 15475 9540 15568 9568
rect 15289 9531 15347 9537
rect 15562 9528 15568 9540
rect 15620 9528 15626 9580
rect 15657 9571 15715 9577
rect 15657 9537 15669 9571
rect 15703 9537 15715 9571
rect 15930 9568 15936 9580
rect 15891 9540 15936 9568
rect 15657 9531 15715 9537
rect 15672 9500 15700 9531
rect 15930 9528 15936 9540
rect 15988 9528 15994 9580
rect 16206 9568 16212 9580
rect 16167 9540 16212 9568
rect 16206 9528 16212 9540
rect 16264 9568 16270 9580
rect 16316 9568 16344 9608
rect 16264 9540 16344 9568
rect 17037 9571 17095 9577
rect 16264 9528 16270 9540
rect 17037 9537 17049 9571
rect 17083 9568 17095 9571
rect 17586 9568 17592 9580
rect 17083 9540 17592 9568
rect 17083 9537 17095 9540
rect 17037 9531 17095 9537
rect 17586 9528 17592 9540
rect 17644 9528 17650 9580
rect 17494 9500 17500 9512
rect 15672 9472 17500 9500
rect 17494 9460 17500 9472
rect 17552 9460 17558 9512
rect 18064 9509 18092 9608
rect 20064 9605 20076 9639
rect 20110 9636 20122 9639
rect 22020 9636 22048 9667
rect 20110 9608 22048 9636
rect 22664 9636 22692 9676
rect 23014 9664 23020 9716
rect 23072 9704 23078 9716
rect 24670 9704 24676 9716
rect 23072 9676 24676 9704
rect 23072 9664 23078 9676
rect 24670 9664 24676 9676
rect 24728 9664 24734 9716
rect 24946 9664 24952 9716
rect 25004 9704 25010 9716
rect 27525 9707 27583 9713
rect 27525 9704 27537 9707
rect 25004 9676 27537 9704
rect 25004 9664 25010 9676
rect 27525 9673 27537 9676
rect 27571 9704 27583 9707
rect 28166 9704 28172 9716
rect 27571 9676 28172 9704
rect 27571 9673 27583 9676
rect 27525 9667 27583 9673
rect 28166 9664 28172 9676
rect 28224 9664 28230 9716
rect 28442 9664 28448 9716
rect 28500 9704 28506 9716
rect 29273 9707 29331 9713
rect 29273 9704 29285 9707
rect 28500 9676 29285 9704
rect 28500 9664 28506 9676
rect 29273 9673 29285 9676
rect 29319 9673 29331 9707
rect 29454 9704 29460 9716
rect 29415 9676 29460 9704
rect 29273 9667 29331 9673
rect 29454 9664 29460 9676
rect 29512 9664 29518 9716
rect 29546 9664 29552 9716
rect 29604 9704 29610 9716
rect 31938 9704 31944 9716
rect 29604 9676 29649 9704
rect 30300 9676 31944 9704
rect 29604 9664 29610 9676
rect 23566 9636 23572 9648
rect 22664 9608 23572 9636
rect 20110 9605 20122 9608
rect 20064 9599 20122 9605
rect 23566 9596 23572 9608
rect 23624 9596 23630 9648
rect 23661 9639 23719 9645
rect 23661 9605 23673 9639
rect 23707 9636 23719 9639
rect 27341 9639 27399 9645
rect 23707 9608 26004 9636
rect 23707 9605 23719 9608
rect 23661 9599 23719 9605
rect 25976 9580 26004 9608
rect 27341 9605 27353 9639
rect 27387 9605 27399 9639
rect 28350 9636 28356 9648
rect 28311 9608 28356 9636
rect 27341 9599 27399 9605
rect 18877 9571 18935 9577
rect 18877 9537 18889 9571
rect 18923 9568 18935 9571
rect 21174 9568 21180 9580
rect 18923 9540 21180 9568
rect 18923 9537 18935 9540
rect 18877 9531 18935 9537
rect 21174 9528 21180 9540
rect 21232 9528 21238 9580
rect 21726 9528 21732 9580
rect 21784 9568 21790 9580
rect 21784 9540 22600 9568
rect 21784 9528 21790 9540
rect 18049 9503 18107 9509
rect 18049 9469 18061 9503
rect 18095 9500 18107 9503
rect 18782 9500 18788 9512
rect 18095 9472 18788 9500
rect 18095 9469 18107 9472
rect 18049 9463 18107 9469
rect 18782 9460 18788 9472
rect 18840 9460 18846 9512
rect 19150 9500 19156 9512
rect 19111 9472 19156 9500
rect 19150 9460 19156 9472
rect 19208 9460 19214 9512
rect 19426 9460 19432 9512
rect 19484 9500 19490 9512
rect 19797 9503 19855 9509
rect 19797 9500 19809 9503
rect 19484 9472 19809 9500
rect 19484 9460 19490 9472
rect 19797 9469 19809 9472
rect 19843 9469 19855 9503
rect 19797 9463 19855 9469
rect 21082 9460 21088 9512
rect 21140 9500 21146 9512
rect 22572 9509 22600 9540
rect 23934 9528 23940 9580
rect 23992 9568 23998 9580
rect 24029 9571 24087 9577
rect 24029 9568 24041 9571
rect 23992 9540 24041 9568
rect 23992 9528 23998 9540
rect 24029 9537 24041 9540
rect 24075 9537 24087 9571
rect 24029 9531 24087 9537
rect 24121 9571 24179 9577
rect 24121 9537 24133 9571
rect 24167 9537 24179 9571
rect 24121 9531 24179 9537
rect 24213 9571 24271 9577
rect 24213 9537 24225 9571
rect 24259 9568 24271 9571
rect 25038 9568 25044 9580
rect 24259 9540 25044 9568
rect 24259 9537 24271 9540
rect 24213 9531 24271 9537
rect 22465 9503 22523 9509
rect 22465 9500 22477 9503
rect 21140 9472 22477 9500
rect 21140 9460 21146 9472
rect 22465 9469 22477 9472
rect 22511 9469 22523 9503
rect 22465 9463 22523 9469
rect 22557 9503 22615 9509
rect 22557 9469 22569 9503
rect 22603 9469 22615 9503
rect 23474 9500 23480 9512
rect 23435 9472 23480 9500
rect 22557 9463 22615 9469
rect 23474 9460 23480 9472
rect 23532 9460 23538 9512
rect 24136 9500 24164 9531
rect 25038 9528 25044 9540
rect 25096 9568 25102 9580
rect 25225 9571 25283 9577
rect 25225 9568 25237 9571
rect 25096 9540 25237 9568
rect 25096 9528 25102 9540
rect 25225 9537 25237 9540
rect 25271 9537 25283 9571
rect 25406 9568 25412 9580
rect 25367 9540 25412 9568
rect 25225 9531 25283 9537
rect 25406 9528 25412 9540
rect 25464 9528 25470 9580
rect 25498 9528 25504 9580
rect 25556 9568 25562 9580
rect 25593 9571 25651 9577
rect 25593 9568 25605 9571
rect 25556 9540 25605 9568
rect 25556 9528 25562 9540
rect 25593 9537 25605 9540
rect 25639 9537 25651 9571
rect 25866 9568 25872 9580
rect 25827 9540 25872 9568
rect 25593 9531 25651 9537
rect 25866 9528 25872 9540
rect 25924 9528 25930 9580
rect 25958 9528 25964 9580
rect 26016 9568 26022 9580
rect 26145 9571 26203 9577
rect 26145 9568 26157 9571
rect 26016 9540 26157 9568
rect 26016 9528 26022 9540
rect 26145 9537 26157 9540
rect 26191 9537 26203 9571
rect 26145 9531 26203 9537
rect 24302 9500 24308 9512
rect 24136 9472 24308 9500
rect 24302 9460 24308 9472
rect 24360 9460 24366 9512
rect 24765 9503 24823 9509
rect 24765 9469 24777 9503
rect 24811 9500 24823 9503
rect 26602 9500 26608 9512
rect 24811 9472 26608 9500
rect 24811 9469 24823 9472
rect 24765 9463 24823 9469
rect 26602 9460 26608 9472
rect 26660 9460 26666 9512
rect 14921 9435 14979 9441
rect 14921 9401 14933 9435
rect 14967 9432 14979 9435
rect 15194 9432 15200 9444
rect 14967 9404 15200 9432
rect 14967 9401 14979 9404
rect 14921 9395 14979 9401
rect 15194 9392 15200 9404
rect 15252 9432 15258 9444
rect 16298 9432 16304 9444
rect 15252 9404 16304 9432
rect 15252 9392 15258 9404
rect 16298 9392 16304 9404
rect 16356 9392 16362 9444
rect 16482 9392 16488 9444
rect 16540 9432 16546 9444
rect 19168 9432 19196 9460
rect 27157 9435 27215 9441
rect 27157 9432 27169 9435
rect 16540 9404 19196 9432
rect 20732 9404 27169 9432
rect 16540 9392 16546 9404
rect 13688 9336 14872 9364
rect 13688 9324 13694 9336
rect 15654 9324 15660 9376
rect 15712 9364 15718 9376
rect 20732 9364 20760 9404
rect 27157 9401 27169 9404
rect 27203 9401 27215 9435
rect 27356 9432 27384 9599
rect 28350 9596 28356 9608
rect 28408 9596 28414 9648
rect 29730 9636 29736 9648
rect 29691 9608 29736 9636
rect 29730 9596 29736 9608
rect 29788 9596 29794 9648
rect 30300 9580 30328 9676
rect 31938 9664 31944 9676
rect 31996 9664 32002 9716
rect 32122 9664 32128 9716
rect 32180 9704 32186 9716
rect 32493 9707 32551 9713
rect 32493 9704 32505 9707
rect 32180 9676 32505 9704
rect 32180 9664 32186 9676
rect 32493 9673 32505 9676
rect 32539 9673 32551 9707
rect 32493 9667 32551 9673
rect 32674 9664 32680 9716
rect 32732 9704 32738 9716
rect 32950 9704 32956 9716
rect 32732 9676 32956 9704
rect 32732 9664 32738 9676
rect 32950 9664 32956 9676
rect 33008 9664 33014 9716
rect 33318 9704 33324 9716
rect 33376 9713 33382 9716
rect 33285 9676 33324 9704
rect 33318 9664 33324 9676
rect 33376 9667 33385 9713
rect 33376 9664 33382 9667
rect 33686 9664 33692 9716
rect 33744 9704 33750 9716
rect 38378 9704 38384 9716
rect 33744 9676 38384 9704
rect 33744 9664 33750 9676
rect 38378 9664 38384 9676
rect 38436 9664 38442 9716
rect 46569 9707 46627 9713
rect 46569 9673 46581 9707
rect 46615 9704 46627 9707
rect 46658 9704 46664 9716
rect 46615 9676 46664 9704
rect 46615 9673 46627 9676
rect 46569 9667 46627 9673
rect 46658 9664 46664 9676
rect 46716 9664 46722 9716
rect 31294 9596 31300 9648
rect 31352 9636 31358 9648
rect 33962 9636 33968 9648
rect 31352 9608 33968 9636
rect 31352 9596 31358 9608
rect 33962 9596 33968 9608
rect 34020 9636 34026 9648
rect 37737 9639 37795 9645
rect 37737 9636 37749 9639
rect 34020 9608 37749 9636
rect 34020 9596 34026 9608
rect 37737 9605 37749 9608
rect 37783 9605 37795 9639
rect 37737 9599 37795 9605
rect 38933 9639 38991 9645
rect 38933 9605 38945 9639
rect 38979 9636 38991 9639
rect 39206 9636 39212 9648
rect 38979 9608 39212 9636
rect 38979 9605 38991 9608
rect 38933 9599 38991 9605
rect 39206 9596 39212 9608
rect 39264 9596 39270 9648
rect 43993 9639 44051 9645
rect 43993 9605 44005 9639
rect 44039 9636 44051 9639
rect 44266 9636 44272 9648
rect 44039 9608 44272 9636
rect 44039 9605 44051 9608
rect 43993 9599 44051 9605
rect 44266 9596 44272 9608
rect 44324 9596 44330 9648
rect 45462 9645 45468 9648
rect 45456 9636 45468 9645
rect 45423 9608 45468 9636
rect 45456 9599 45468 9608
rect 45462 9596 45468 9599
rect 45520 9596 45526 9648
rect 27479 9571 27537 9577
rect 27479 9537 27491 9571
rect 27525 9568 27537 9571
rect 27614 9568 27620 9580
rect 27525 9540 27620 9568
rect 27525 9537 27537 9540
rect 27479 9531 27537 9537
rect 27614 9528 27620 9540
rect 27672 9528 27678 9580
rect 27709 9571 27767 9577
rect 27709 9537 27721 9571
rect 27755 9537 27767 9571
rect 27709 9531 27767 9537
rect 28169 9571 28227 9577
rect 28169 9537 28181 9571
rect 28215 9537 28227 9571
rect 28169 9531 28227 9537
rect 27522 9432 27528 9444
rect 27356 9404 27528 9432
rect 27157 9395 27215 9401
rect 27522 9392 27528 9404
rect 27580 9392 27586 9444
rect 15712 9336 20760 9364
rect 15712 9324 15718 9336
rect 21082 9324 21088 9376
rect 21140 9364 21146 9376
rect 21177 9367 21235 9373
rect 21177 9364 21189 9367
rect 21140 9336 21189 9364
rect 21140 9324 21146 9336
rect 21177 9333 21189 9336
rect 21223 9333 21235 9367
rect 21177 9327 21235 9333
rect 23014 9324 23020 9376
rect 23072 9364 23078 9376
rect 23934 9364 23940 9376
rect 23072 9336 23940 9364
rect 23072 9324 23078 9336
rect 23934 9324 23940 9336
rect 23992 9324 23998 9376
rect 24762 9324 24768 9376
rect 24820 9364 24826 9376
rect 27724 9364 27752 9531
rect 28184 9500 28212 9531
rect 28442 9528 28448 9580
rect 28500 9568 28506 9580
rect 28583 9571 28641 9577
rect 28500 9540 28545 9568
rect 28500 9528 28506 9540
rect 28583 9537 28595 9571
rect 28629 9568 28641 9571
rect 29270 9568 29276 9580
rect 28629 9540 29276 9568
rect 28629 9537 28641 9540
rect 28583 9531 28641 9537
rect 29104 9512 29132 9540
rect 29270 9528 29276 9540
rect 29328 9528 29334 9580
rect 29365 9571 29423 9577
rect 29365 9537 29377 9571
rect 29411 9537 29423 9571
rect 29365 9531 29423 9537
rect 30193 9571 30251 9577
rect 30193 9537 30205 9571
rect 30239 9568 30251 9571
rect 30282 9568 30288 9580
rect 30239 9540 30288 9568
rect 30239 9537 30251 9540
rect 30193 9531 30251 9537
rect 28810 9500 28816 9512
rect 28184 9472 28816 9500
rect 28810 9460 28816 9472
rect 28868 9460 28874 9512
rect 28920 9472 29045 9500
rect 28721 9435 28779 9441
rect 28721 9401 28733 9435
rect 28767 9432 28779 9435
rect 28920 9432 28948 9472
rect 28767 9404 28948 9432
rect 28767 9401 28779 9404
rect 28721 9395 28779 9401
rect 29017 9376 29045 9472
rect 29086 9460 29092 9512
rect 29144 9460 29150 9512
rect 29380 9500 29408 9531
rect 30282 9528 30288 9540
rect 30340 9568 30346 9580
rect 31018 9568 31024 9580
rect 30340 9540 30433 9568
rect 30979 9540 31024 9568
rect 30340 9528 30346 9540
rect 31018 9528 31024 9540
rect 31076 9528 31082 9580
rect 31754 9528 31760 9580
rect 31812 9568 31818 9580
rect 32585 9571 32643 9577
rect 32585 9568 32597 9571
rect 31812 9540 32597 9568
rect 31812 9528 31818 9540
rect 32585 9537 32597 9540
rect 32631 9537 32643 9571
rect 32585 9531 32643 9537
rect 32600 9500 32628 9531
rect 32674 9528 32680 9580
rect 32732 9568 32738 9580
rect 32769 9571 32827 9577
rect 32769 9568 32781 9571
rect 32732 9540 32781 9568
rect 32732 9528 32738 9540
rect 32769 9537 32781 9540
rect 32815 9537 32827 9571
rect 32769 9531 32827 9537
rect 33229 9571 33287 9577
rect 33229 9537 33241 9571
rect 33275 9537 33287 9571
rect 33410 9568 33416 9580
rect 33371 9540 33416 9568
rect 33229 9531 33287 9537
rect 33134 9500 33140 9512
rect 29380 9472 29868 9500
rect 32600 9472 33140 9500
rect 29840 9376 29868 9472
rect 33134 9460 33140 9472
rect 33192 9460 33198 9512
rect 33244 9500 33272 9531
rect 33410 9528 33416 9540
rect 33468 9528 33474 9580
rect 33505 9571 33563 9577
rect 33505 9537 33517 9571
rect 33551 9568 33563 9571
rect 33686 9568 33692 9580
rect 33551 9540 33692 9568
rect 33551 9537 33563 9540
rect 33505 9531 33563 9537
rect 33686 9528 33692 9540
rect 33744 9528 33750 9580
rect 35986 9568 35992 9580
rect 35947 9540 35992 9568
rect 35986 9528 35992 9540
rect 36044 9528 36050 9580
rect 36173 9571 36231 9577
rect 36173 9537 36185 9571
rect 36219 9568 36231 9571
rect 36538 9568 36544 9580
rect 36219 9540 36544 9568
rect 36219 9537 36231 9540
rect 36173 9531 36231 9537
rect 36538 9528 36544 9540
rect 36596 9528 36602 9580
rect 37458 9568 37464 9580
rect 37419 9540 37464 9568
rect 37458 9528 37464 9540
rect 37516 9528 37522 9580
rect 37609 9571 37667 9577
rect 37609 9537 37621 9571
rect 37655 9568 37667 9571
rect 37655 9540 37780 9568
rect 37655 9537 37667 9540
rect 37609 9531 37667 9537
rect 33870 9500 33876 9512
rect 33244 9472 33876 9500
rect 33870 9460 33876 9472
rect 33928 9460 33934 9512
rect 37752 9500 37780 9540
rect 37826 9528 37832 9580
rect 37884 9568 37890 9580
rect 37967 9571 38025 9577
rect 37884 9540 37929 9568
rect 37884 9528 37890 9540
rect 37967 9537 37979 9571
rect 38013 9568 38025 9571
rect 38102 9568 38108 9580
rect 38013 9540 38108 9568
rect 38013 9537 38025 9540
rect 37967 9531 38025 9537
rect 38102 9528 38108 9540
rect 38160 9528 38166 9580
rect 38562 9568 38568 9580
rect 38523 9540 38568 9568
rect 38562 9528 38568 9540
rect 38620 9528 38626 9580
rect 38654 9528 38660 9580
rect 38712 9568 38718 9580
rect 38838 9568 38844 9580
rect 38712 9540 38757 9568
rect 38799 9540 38844 9568
rect 38712 9528 38718 9540
rect 38838 9528 38844 9540
rect 38896 9528 38902 9580
rect 39071 9571 39129 9577
rect 39071 9537 39083 9571
rect 39117 9568 39129 9571
rect 40586 9568 40592 9580
rect 39117 9540 40592 9568
rect 39117 9537 39129 9540
rect 39071 9531 39129 9537
rect 40586 9528 40592 9540
rect 40644 9528 40650 9580
rect 40770 9528 40776 9580
rect 40828 9568 40834 9580
rect 42426 9568 42432 9580
rect 40828 9540 42432 9568
rect 40828 9528 40834 9540
rect 42426 9528 42432 9540
rect 42484 9528 42490 9580
rect 44085 9571 44143 9577
rect 44085 9537 44097 9571
rect 44131 9537 44143 9571
rect 44085 9531 44143 9537
rect 37752 9472 38884 9500
rect 38856 9444 38884 9472
rect 43990 9460 43996 9512
rect 44048 9500 44054 9512
rect 44100 9500 44128 9531
rect 44174 9528 44180 9580
rect 44232 9568 44238 9580
rect 45186 9568 45192 9580
rect 44232 9540 44277 9568
rect 45147 9540 45192 9568
rect 44232 9528 44238 9540
rect 45186 9528 45192 9540
rect 45244 9528 45250 9580
rect 46290 9568 46296 9580
rect 45296 9540 46296 9568
rect 45296 9500 45324 9540
rect 46290 9528 46296 9540
rect 46348 9528 46354 9580
rect 56962 9568 56968 9580
rect 56923 9540 56968 9568
rect 56962 9528 56968 9540
rect 57020 9528 57026 9580
rect 57054 9528 57060 9580
rect 57112 9568 57118 9580
rect 57149 9571 57207 9577
rect 57149 9568 57161 9571
rect 57112 9540 57161 9568
rect 57112 9528 57118 9540
rect 57149 9537 57161 9540
rect 57195 9537 57207 9571
rect 57149 9531 57207 9537
rect 44048 9472 45324 9500
rect 44048 9460 44054 9472
rect 31662 9392 31668 9444
rect 31720 9432 31726 9444
rect 34514 9432 34520 9444
rect 31720 9404 34520 9432
rect 31720 9392 31726 9404
rect 34514 9392 34520 9404
rect 34572 9392 34578 9444
rect 35158 9392 35164 9444
rect 35216 9432 35222 9444
rect 35216 9404 38792 9432
rect 35216 9392 35222 9404
rect 24820 9336 27752 9364
rect 24820 9324 24826 9336
rect 28994 9324 29000 9376
rect 29052 9324 29058 9376
rect 29822 9324 29828 9376
rect 29880 9364 29886 9376
rect 30377 9367 30435 9373
rect 30377 9364 30389 9367
rect 29880 9336 30389 9364
rect 29880 9324 29886 9336
rect 30377 9333 30389 9336
rect 30423 9364 30435 9367
rect 31018 9364 31024 9376
rect 30423 9336 31024 9364
rect 30423 9333 30435 9336
rect 30377 9327 30435 9333
rect 31018 9324 31024 9336
rect 31076 9324 31082 9376
rect 31297 9367 31355 9373
rect 31297 9333 31309 9367
rect 31343 9364 31355 9367
rect 31570 9364 31576 9376
rect 31343 9336 31576 9364
rect 31343 9333 31355 9336
rect 31297 9327 31355 9333
rect 31570 9324 31576 9336
rect 31628 9324 31634 9376
rect 32309 9367 32367 9373
rect 32309 9333 32321 9367
rect 32355 9364 32367 9367
rect 32582 9364 32588 9376
rect 32355 9336 32588 9364
rect 32355 9333 32367 9336
rect 32309 9327 32367 9333
rect 32582 9324 32588 9336
rect 32640 9364 32646 9376
rect 35894 9364 35900 9376
rect 32640 9336 35900 9364
rect 32640 9324 32646 9336
rect 35894 9324 35900 9336
rect 35952 9324 35958 9376
rect 35989 9367 36047 9373
rect 35989 9333 36001 9367
rect 36035 9364 36047 9367
rect 36262 9364 36268 9376
rect 36035 9336 36268 9364
rect 36035 9333 36047 9336
rect 35989 9327 36047 9333
rect 36262 9324 36268 9336
rect 36320 9324 36326 9376
rect 37550 9324 37556 9376
rect 37608 9364 37614 9376
rect 38105 9367 38163 9373
rect 38105 9364 38117 9367
rect 37608 9336 38117 9364
rect 37608 9324 37614 9336
rect 38105 9333 38117 9336
rect 38151 9333 38163 9367
rect 38764 9364 38792 9404
rect 38838 9392 38844 9444
rect 38896 9392 38902 9444
rect 39209 9435 39267 9441
rect 39209 9432 39221 9435
rect 38948 9404 39221 9432
rect 38948 9364 38976 9404
rect 39209 9401 39221 9404
rect 39255 9401 39267 9435
rect 39209 9395 39267 9401
rect 39298 9392 39304 9444
rect 39356 9432 39362 9444
rect 43809 9435 43867 9441
rect 43809 9432 43821 9435
rect 39356 9404 43821 9432
rect 39356 9392 39362 9404
rect 43809 9401 43821 9404
rect 43855 9432 43867 9435
rect 44450 9432 44456 9444
rect 43855 9404 44456 9432
rect 43855 9401 43867 9404
rect 43809 9395 43867 9401
rect 44450 9392 44456 9404
rect 44508 9392 44514 9444
rect 38764 9336 38976 9364
rect 38105 9327 38163 9333
rect 40310 9324 40316 9376
rect 40368 9364 40374 9376
rect 44361 9367 44419 9373
rect 44361 9364 44373 9367
rect 40368 9336 44373 9364
rect 40368 9324 40374 9336
rect 44361 9333 44373 9336
rect 44407 9333 44419 9367
rect 44361 9327 44419 9333
rect 56318 9324 56324 9376
rect 56376 9364 56382 9376
rect 57057 9367 57115 9373
rect 57057 9364 57069 9367
rect 56376 9336 57069 9364
rect 56376 9324 56382 9336
rect 57057 9333 57069 9336
rect 57103 9333 57115 9367
rect 57057 9327 57115 9333
rect 1104 9274 58880 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 58880 9274
rect 1104 9200 58880 9222
rect 13357 9163 13415 9169
rect 13357 9129 13369 9163
rect 13403 9160 13415 9163
rect 13814 9160 13820 9172
rect 13403 9132 13820 9160
rect 13403 9129 13415 9132
rect 13357 9123 13415 9129
rect 13814 9120 13820 9132
rect 13872 9120 13878 9172
rect 15194 9160 15200 9172
rect 13924 9132 15200 9160
rect 13262 9092 13268 9104
rect 13223 9064 13268 9092
rect 13262 9052 13268 9064
rect 13320 9052 13326 9104
rect 13924 9092 13952 9132
rect 15194 9120 15200 9132
rect 15252 9120 15258 9172
rect 16206 9120 16212 9172
rect 16264 9160 16270 9172
rect 21082 9160 21088 9172
rect 16264 9132 21088 9160
rect 16264 9120 16270 9132
rect 21082 9120 21088 9132
rect 21140 9120 21146 9172
rect 21266 9160 21272 9172
rect 21227 9132 21272 9160
rect 21266 9120 21272 9132
rect 21324 9120 21330 9172
rect 23658 9120 23664 9172
rect 23716 9160 23722 9172
rect 27062 9160 27068 9172
rect 23716 9132 27068 9160
rect 23716 9120 23722 9132
rect 27062 9120 27068 9132
rect 27120 9120 27126 9172
rect 27982 9120 27988 9172
rect 28040 9160 28046 9172
rect 28445 9163 28503 9169
rect 28445 9160 28457 9163
rect 28040 9132 28457 9160
rect 28040 9120 28046 9132
rect 28445 9129 28457 9132
rect 28491 9129 28503 9163
rect 30282 9160 30288 9172
rect 28445 9123 28503 9129
rect 29656 9132 30288 9160
rect 13372 9064 13952 9092
rect 14737 9095 14795 9101
rect 10686 8984 10692 9036
rect 10744 9024 10750 9036
rect 13372 9024 13400 9064
rect 14737 9061 14749 9095
rect 14783 9092 14795 9095
rect 23566 9092 23572 9104
rect 14783 9064 23572 9092
rect 14783 9061 14795 9064
rect 14737 9055 14795 9061
rect 23566 9052 23572 9064
rect 23624 9052 23630 9104
rect 24026 9052 24032 9104
rect 24084 9092 24090 9104
rect 24394 9092 24400 9104
rect 24084 9064 24400 9092
rect 24084 9052 24090 9064
rect 24394 9052 24400 9064
rect 24452 9052 24458 9104
rect 25866 9092 25872 9104
rect 24688 9064 25872 9092
rect 10744 8996 13400 9024
rect 10744 8984 10750 8996
rect 13538 8984 13544 9036
rect 13596 9024 13602 9036
rect 13596 8996 15332 9024
rect 13596 8984 13602 8996
rect 1581 8959 1639 8965
rect 1581 8925 1593 8959
rect 1627 8956 1639 8959
rect 8294 8956 8300 8968
rect 1627 8928 8300 8956
rect 1627 8925 1639 8928
rect 1581 8919 1639 8925
rect 8294 8916 8300 8928
rect 8352 8916 8358 8968
rect 14274 8916 14280 8968
rect 14332 8956 14338 8968
rect 15304 8965 15332 8996
rect 17586 8984 17592 9036
rect 17644 9024 17650 9036
rect 18325 9027 18383 9033
rect 18325 9024 18337 9027
rect 17644 8996 18337 9024
rect 17644 8984 17650 8996
rect 18325 8993 18337 8996
rect 18371 8993 18383 9027
rect 18325 8987 18383 8993
rect 15289 8959 15347 8965
rect 14332 8928 15148 8956
rect 14332 8916 14338 8928
rect 1854 8888 1860 8900
rect 1815 8860 1860 8888
rect 1854 8848 1860 8860
rect 1912 8848 1918 8900
rect 12434 8848 12440 8900
rect 12492 8888 12498 8900
rect 12897 8891 12955 8897
rect 12897 8888 12909 8891
rect 12492 8860 12909 8888
rect 12492 8848 12498 8860
rect 12897 8857 12909 8860
rect 12943 8857 12955 8891
rect 12897 8851 12955 8857
rect 13630 8848 13636 8900
rect 13688 8888 13694 8900
rect 14918 8888 14924 8900
rect 13688 8860 14924 8888
rect 13688 8848 13694 8860
rect 14918 8848 14924 8860
rect 14976 8848 14982 8900
rect 15120 8832 15148 8928
rect 15289 8925 15301 8959
rect 15335 8956 15347 8959
rect 17034 8956 17040 8968
rect 15335 8928 17040 8956
rect 15335 8925 15347 8928
rect 15289 8919 15347 8925
rect 17034 8916 17040 8928
rect 17092 8916 17098 8968
rect 18049 8959 18107 8965
rect 18049 8934 18061 8959
rect 18095 8934 18107 8959
rect 15749 8891 15807 8897
rect 15749 8857 15761 8891
rect 15795 8888 15807 8891
rect 17494 8888 17500 8900
rect 15795 8860 17356 8888
rect 17455 8860 17500 8888
rect 15795 8857 15807 8860
rect 15749 8851 15807 8857
rect 13446 8780 13452 8832
rect 13504 8820 13510 8832
rect 15013 8823 15071 8829
rect 15013 8820 15025 8823
rect 13504 8792 15025 8820
rect 13504 8780 13510 8792
rect 15013 8789 15025 8792
rect 15059 8789 15071 8823
rect 15013 8783 15071 8789
rect 15102 8780 15108 8832
rect 15160 8820 15166 8832
rect 17328 8820 17356 8860
rect 17494 8848 17500 8860
rect 17552 8848 17558 8900
rect 18046 8882 18052 8934
rect 18104 8882 18110 8934
rect 18340 8888 18368 8987
rect 18782 8984 18788 9036
rect 18840 9024 18846 9036
rect 24688 9033 24716 9064
rect 25866 9052 25872 9064
rect 25924 9052 25930 9104
rect 28166 9052 28172 9104
rect 28224 9092 28230 9104
rect 29656 9092 29684 9132
rect 30282 9120 30288 9132
rect 30340 9160 30346 9172
rect 30340 9132 30788 9160
rect 30340 9120 30346 9132
rect 28224 9064 29684 9092
rect 28224 9052 28230 9064
rect 29730 9052 29736 9104
rect 29788 9092 29794 9104
rect 30650 9092 30656 9104
rect 29788 9064 30656 9092
rect 29788 9052 29794 9064
rect 30650 9052 30656 9064
rect 30708 9052 30714 9104
rect 24673 9027 24731 9033
rect 18840 8996 24624 9024
rect 18840 8984 18846 8996
rect 19889 8959 19947 8965
rect 19889 8925 19901 8959
rect 19935 8956 19947 8959
rect 19935 8928 22094 8956
rect 19935 8925 19947 8928
rect 19889 8919 19947 8925
rect 21542 8888 21548 8900
rect 18340 8860 21548 8888
rect 21542 8848 21548 8860
rect 21600 8848 21606 8900
rect 22066 8888 22094 8928
rect 22462 8916 22468 8968
rect 22520 8956 22526 8968
rect 23477 8959 23535 8965
rect 23477 8956 23489 8959
rect 22520 8928 23489 8956
rect 22520 8916 22526 8928
rect 23477 8925 23489 8928
rect 23523 8925 23535 8959
rect 23658 8956 23664 8968
rect 23619 8928 23664 8956
rect 23477 8919 23535 8925
rect 23658 8916 23664 8928
rect 23716 8916 23722 8968
rect 24118 8956 24124 8968
rect 23768 8928 24124 8956
rect 23382 8888 23388 8900
rect 22066 8860 23388 8888
rect 23382 8848 23388 8860
rect 23440 8848 23446 8900
rect 18782 8820 18788 8832
rect 15160 8792 15253 8820
rect 17328 8792 18788 8820
rect 15160 8780 15166 8792
rect 18782 8780 18788 8792
rect 18840 8820 18846 8832
rect 19058 8820 19064 8832
rect 18840 8792 19064 8820
rect 18840 8780 18846 8792
rect 19058 8780 19064 8792
rect 19116 8780 19122 8832
rect 21174 8780 21180 8832
rect 21232 8820 21238 8832
rect 23014 8820 23020 8832
rect 21232 8792 23020 8820
rect 21232 8780 21238 8792
rect 23014 8780 23020 8792
rect 23072 8780 23078 8832
rect 23768 8829 23796 8928
rect 24118 8916 24124 8928
rect 24176 8916 24182 8968
rect 24596 8956 24624 8996
rect 24673 8993 24685 9027
rect 24719 8993 24731 9027
rect 25958 9024 25964 9036
rect 24673 8987 24731 8993
rect 25148 8996 25964 9024
rect 24765 8959 24823 8965
rect 24596 8928 24716 8956
rect 24026 8888 24032 8900
rect 23987 8860 24032 8888
rect 24026 8848 24032 8860
rect 24084 8848 24090 8900
rect 24688 8888 24716 8928
rect 24765 8925 24777 8959
rect 24811 8956 24823 8959
rect 25148 8956 25176 8996
rect 25958 8984 25964 8996
rect 26016 8984 26022 9036
rect 27430 9024 27436 9036
rect 26252 8996 27436 9024
rect 24811 8928 25176 8956
rect 25225 8959 25283 8965
rect 24811 8925 24823 8928
rect 24765 8919 24823 8925
rect 25225 8925 25237 8959
rect 25271 8956 25283 8959
rect 25314 8956 25320 8968
rect 25271 8928 25320 8956
rect 25271 8925 25283 8928
rect 25225 8919 25283 8925
rect 25314 8916 25320 8928
rect 25372 8916 25378 8968
rect 25682 8956 25688 8968
rect 25643 8928 25688 8956
rect 25682 8916 25688 8928
rect 25740 8916 25746 8968
rect 25774 8916 25780 8968
rect 25832 8956 25838 8968
rect 26252 8965 26280 8996
rect 27430 8984 27436 8996
rect 27488 8984 27494 9036
rect 27890 9024 27896 9036
rect 27851 8996 27896 9024
rect 27890 8984 27896 8996
rect 27948 8984 27954 9036
rect 29089 9027 29147 9033
rect 29089 8993 29101 9027
rect 29135 9024 29147 9027
rect 29178 9024 29184 9036
rect 29135 8996 29184 9024
rect 29135 8993 29147 8996
rect 29089 8987 29147 8993
rect 29178 8984 29184 8996
rect 29236 9024 29242 9036
rect 30098 9024 30104 9036
rect 29236 8996 30104 9024
rect 29236 8984 29242 8996
rect 30098 8984 30104 8996
rect 30156 8984 30162 9036
rect 30760 9033 30788 9132
rect 32490 9120 32496 9172
rect 32548 9160 32554 9172
rect 33686 9160 33692 9172
rect 32548 9132 33692 9160
rect 32548 9120 32554 9132
rect 33686 9120 33692 9132
rect 33744 9120 33750 9172
rect 34146 9120 34152 9172
rect 34204 9160 34210 9172
rect 35986 9160 35992 9172
rect 34204 9132 35992 9160
rect 34204 9120 34210 9132
rect 35986 9120 35992 9132
rect 36044 9160 36050 9172
rect 38930 9160 38936 9172
rect 36044 9132 38936 9160
rect 36044 9120 36050 9132
rect 38930 9120 38936 9132
rect 38988 9160 38994 9172
rect 39025 9163 39083 9169
rect 39025 9160 39037 9163
rect 38988 9132 39037 9160
rect 38988 9120 38994 9132
rect 39025 9129 39037 9132
rect 39071 9129 39083 9163
rect 41322 9160 41328 9172
rect 39025 9123 39083 9129
rect 39408 9132 41328 9160
rect 31386 9092 31392 9104
rect 31347 9064 31392 9092
rect 31386 9052 31392 9064
rect 31444 9052 31450 9104
rect 32582 9052 32588 9104
rect 32640 9092 32646 9104
rect 32861 9095 32919 9101
rect 32861 9092 32873 9095
rect 32640 9064 32873 9092
rect 32640 9052 32646 9064
rect 32861 9061 32873 9064
rect 32907 9061 32919 9095
rect 32861 9055 32919 9061
rect 33134 9052 33140 9104
rect 33192 9092 33198 9104
rect 34164 9092 34192 9120
rect 36446 9092 36452 9104
rect 33192 9064 34192 9092
rect 36096 9064 36452 9092
rect 33192 9052 33198 9064
rect 30745 9027 30803 9033
rect 30745 8993 30757 9027
rect 30791 8993 30803 9027
rect 34422 9024 34428 9036
rect 30745 8987 30803 8993
rect 33796 8996 34428 9024
rect 25869 8959 25927 8965
rect 25869 8956 25881 8959
rect 25832 8928 25881 8956
rect 25832 8916 25838 8928
rect 25869 8925 25881 8928
rect 25915 8925 25927 8959
rect 25869 8919 25927 8925
rect 26237 8959 26295 8965
rect 26237 8925 26249 8959
rect 26283 8925 26295 8959
rect 26418 8956 26424 8968
rect 26379 8928 26424 8956
rect 26237 8919 26295 8925
rect 26418 8916 26424 8928
rect 26476 8916 26482 8968
rect 26605 8959 26663 8965
rect 26605 8925 26617 8959
rect 26651 8925 26663 8959
rect 26605 8919 26663 8925
rect 27617 8959 27675 8965
rect 27617 8925 27629 8959
rect 27663 8925 27675 8959
rect 27798 8956 27804 8968
rect 27759 8928 27804 8956
rect 27617 8919 27675 8925
rect 26326 8888 26332 8900
rect 24688 8860 26332 8888
rect 26326 8848 26332 8860
rect 26384 8888 26390 8900
rect 26620 8888 26648 8919
rect 26384 8860 27384 8888
rect 26384 8848 26390 8860
rect 23753 8823 23811 8829
rect 23753 8789 23765 8823
rect 23799 8789 23811 8823
rect 23753 8783 23811 8789
rect 23842 8780 23848 8832
rect 23900 8820 23906 8832
rect 24946 8820 24952 8832
rect 23900 8792 24952 8820
rect 23900 8780 23906 8792
rect 24946 8780 24952 8792
rect 25004 8780 25010 8832
rect 26510 8780 26516 8832
rect 26568 8820 26574 8832
rect 26970 8820 26976 8832
rect 26568 8792 26976 8820
rect 26568 8780 26574 8792
rect 26970 8780 26976 8792
rect 27028 8820 27034 8832
rect 27065 8823 27123 8829
rect 27065 8820 27077 8823
rect 27028 8792 27077 8820
rect 27028 8780 27034 8792
rect 27065 8789 27077 8792
rect 27111 8789 27123 8823
rect 27356 8820 27384 8860
rect 27430 8848 27436 8900
rect 27488 8888 27494 8900
rect 27632 8888 27660 8919
rect 27798 8916 27804 8928
rect 27856 8916 27862 8968
rect 27982 8916 27988 8968
rect 28040 8956 28046 8968
rect 30009 8959 30067 8965
rect 30009 8956 30021 8959
rect 28040 8928 30021 8956
rect 28040 8916 28046 8928
rect 30009 8925 30021 8928
rect 30055 8956 30067 8959
rect 31478 8956 31484 8968
rect 30055 8928 31484 8956
rect 30055 8925 30067 8928
rect 30009 8919 30067 8925
rect 31478 8916 31484 8928
rect 31536 8916 31542 8968
rect 31570 8916 31576 8968
rect 31628 8956 31634 8968
rect 32214 8956 32220 8968
rect 31628 8928 32220 8956
rect 31628 8916 31634 8928
rect 32214 8916 32220 8928
rect 32272 8916 32278 8968
rect 33134 8956 33140 8968
rect 33095 8928 33140 8956
rect 33134 8916 33140 8928
rect 33192 8916 33198 8968
rect 33796 8965 33824 8996
rect 34422 8984 34428 8996
rect 34480 9024 34486 9036
rect 36096 9024 36124 9064
rect 36446 9052 36452 9064
rect 36504 9052 36510 9104
rect 36262 9024 36268 9036
rect 34480 8996 36124 9024
rect 36223 8996 36268 9024
rect 34480 8984 34486 8996
rect 36262 8984 36268 8996
rect 36320 8984 36326 9036
rect 37182 8984 37188 9036
rect 37240 9024 37246 9036
rect 38562 9024 38568 9036
rect 37240 8996 37872 9024
rect 37240 8984 37246 8996
rect 33321 8959 33379 8965
rect 33321 8925 33333 8959
rect 33367 8925 33379 8959
rect 33321 8919 33379 8925
rect 33781 8959 33839 8965
rect 33781 8925 33793 8959
rect 33827 8925 33839 8959
rect 33781 8919 33839 8925
rect 27488 8860 27660 8888
rect 27488 8848 27494 8860
rect 28442 8848 28448 8900
rect 28500 8888 28506 8900
rect 28905 8891 28963 8897
rect 28905 8888 28917 8891
rect 28500 8860 28917 8888
rect 28500 8848 28506 8860
rect 28905 8857 28917 8860
rect 28951 8857 28963 8891
rect 28905 8851 28963 8857
rect 29086 8848 29092 8900
rect 29144 8888 29150 8900
rect 30098 8888 30104 8900
rect 29144 8860 30104 8888
rect 29144 8848 29150 8860
rect 30098 8848 30104 8860
rect 30156 8848 30162 8900
rect 31938 8888 31944 8900
rect 31496 8860 31800 8888
rect 31899 8860 31944 8888
rect 27982 8820 27988 8832
rect 27356 8792 27988 8820
rect 27065 8783 27123 8789
rect 27982 8780 27988 8792
rect 28040 8780 28046 8832
rect 28813 8823 28871 8829
rect 28813 8789 28825 8823
rect 28859 8820 28871 8823
rect 29730 8820 29736 8832
rect 28859 8792 29736 8820
rect 28859 8789 28871 8792
rect 28813 8783 28871 8789
rect 29730 8780 29736 8792
rect 29788 8780 29794 8832
rect 30006 8780 30012 8832
rect 30064 8820 30070 8832
rect 31386 8820 31392 8832
rect 30064 8792 31392 8820
rect 30064 8780 30070 8792
rect 31386 8780 31392 8792
rect 31444 8820 31450 8832
rect 31496 8820 31524 8860
rect 31662 8820 31668 8832
rect 31444 8792 31524 8820
rect 31623 8792 31668 8820
rect 31444 8780 31450 8792
rect 31662 8780 31668 8792
rect 31720 8780 31726 8832
rect 31772 8829 31800 8860
rect 31938 8848 31944 8860
rect 31996 8848 32002 8900
rect 33336 8888 33364 8919
rect 34238 8916 34244 8968
rect 34296 8956 34302 8968
rect 35805 8959 35863 8965
rect 35805 8956 35817 8959
rect 34296 8928 35817 8956
rect 34296 8916 34302 8928
rect 35805 8925 35817 8928
rect 35851 8925 35863 8959
rect 35805 8919 35863 8925
rect 35894 8916 35900 8968
rect 35952 8956 35958 8968
rect 36357 8959 36415 8965
rect 36357 8956 36369 8959
rect 35952 8928 36369 8956
rect 35952 8916 35958 8928
rect 36357 8925 36369 8928
rect 36403 8956 36415 8959
rect 37090 8956 37096 8968
rect 36403 8928 37096 8956
rect 36403 8925 36415 8928
rect 36357 8919 36415 8925
rect 37090 8916 37096 8928
rect 37148 8916 37154 8968
rect 37734 8956 37740 8968
rect 37695 8928 37740 8956
rect 37734 8916 37740 8928
rect 37792 8916 37798 8968
rect 37844 8965 37872 8996
rect 38236 8996 38568 9024
rect 38236 8965 38264 8996
rect 38562 8984 38568 8996
rect 38620 9024 38626 9036
rect 39298 9024 39304 9036
rect 38620 8996 39304 9024
rect 38620 8984 38626 8996
rect 39298 8984 39304 8996
rect 39356 8984 39362 9036
rect 37830 8959 37888 8965
rect 37830 8925 37842 8959
rect 37876 8925 37888 8959
rect 38105 8959 38163 8965
rect 38105 8956 38117 8959
rect 37830 8919 37888 8925
rect 37936 8928 38117 8956
rect 32508 8860 33364 8888
rect 31757 8823 31815 8829
rect 31757 8789 31769 8823
rect 31803 8820 31815 8823
rect 32508 8820 32536 8860
rect 33152 8832 33180 8860
rect 33686 8848 33692 8900
rect 33744 8888 33750 8900
rect 34057 8891 34115 8897
rect 34057 8888 34069 8891
rect 33744 8860 34069 8888
rect 33744 8848 33750 8860
rect 34057 8857 34069 8860
rect 34103 8857 34115 8891
rect 34057 8851 34115 8857
rect 37458 8848 37464 8900
rect 37516 8888 37522 8900
rect 37936 8888 37964 8928
rect 38105 8925 38117 8928
rect 38151 8925 38163 8959
rect 38105 8919 38163 8925
rect 38221 8959 38279 8965
rect 38221 8925 38233 8959
rect 38267 8925 38279 8959
rect 38221 8919 38279 8925
rect 38470 8916 38476 8968
rect 38528 8956 38534 8968
rect 39025 8959 39083 8965
rect 39025 8956 39037 8959
rect 38528 8928 39037 8956
rect 38528 8916 38534 8928
rect 39025 8925 39037 8928
rect 39071 8956 39083 8959
rect 39408 8956 39436 9132
rect 41322 9120 41328 9132
rect 41380 9120 41386 9172
rect 46201 9163 46259 9169
rect 46201 9129 46213 9163
rect 46247 9160 46259 9163
rect 46750 9160 46756 9172
rect 46247 9132 46756 9160
rect 46247 9129 46259 9132
rect 46201 9123 46259 9129
rect 46750 9120 46756 9132
rect 46808 9120 46814 9172
rect 40034 9092 40040 9104
rect 39995 9064 40040 9092
rect 40034 9052 40040 9064
rect 40092 9052 40098 9104
rect 41782 9092 41788 9104
rect 40604 9064 41788 9092
rect 40604 9024 40632 9064
rect 41782 9052 41788 9064
rect 41840 9092 41846 9104
rect 56137 9095 56195 9101
rect 41840 9064 55214 9092
rect 41840 9052 41846 9064
rect 44082 9024 44088 9036
rect 40052 8996 40632 9024
rect 40696 8996 44088 9024
rect 40052 8965 40080 8996
rect 39071 8928 39436 8956
rect 40037 8959 40095 8965
rect 39071 8925 39083 8928
rect 39025 8919 39083 8925
rect 40037 8925 40049 8959
rect 40083 8925 40095 8959
rect 40037 8919 40095 8925
rect 40218 8916 40224 8968
rect 40276 8956 40282 8968
rect 40313 8959 40371 8965
rect 40313 8956 40325 8959
rect 40276 8928 40325 8956
rect 40276 8916 40282 8928
rect 40313 8925 40325 8928
rect 40359 8956 40371 8959
rect 40696 8956 40724 8996
rect 44082 8984 44088 8996
rect 44140 8984 44146 9036
rect 44450 9024 44456 9036
rect 44411 8996 44456 9024
rect 44450 8984 44456 8996
rect 44508 8984 44514 9036
rect 45002 8984 45008 9036
rect 45060 9024 45066 9036
rect 46198 9024 46204 9036
rect 45060 8996 46204 9024
rect 45060 8984 45066 8996
rect 46198 8984 46204 8996
rect 46256 8984 46262 9036
rect 40359 8928 40724 8956
rect 40773 8959 40831 8965
rect 40359 8925 40371 8928
rect 40313 8919 40371 8925
rect 40773 8925 40785 8959
rect 40819 8956 40831 8959
rect 40862 8956 40868 8968
rect 40819 8928 40868 8956
rect 40819 8925 40831 8928
rect 40773 8919 40831 8925
rect 40862 8916 40868 8928
rect 40920 8916 40926 8968
rect 45094 8916 45100 8968
rect 45152 8956 45158 8968
rect 45189 8959 45247 8965
rect 45189 8956 45201 8959
rect 45152 8928 45201 8956
rect 45152 8916 45158 8928
rect 45189 8925 45201 8928
rect 45235 8925 45247 8959
rect 46106 8956 46112 8968
rect 46067 8928 46112 8956
rect 45189 8919 45247 8925
rect 46106 8916 46112 8928
rect 46164 8916 46170 8968
rect 46290 8916 46296 8968
rect 46348 8956 46354 8968
rect 46842 8956 46848 8968
rect 46348 8928 46848 8956
rect 46348 8916 46354 8928
rect 46842 8916 46848 8928
rect 46900 8916 46906 8968
rect 55186 8956 55214 9064
rect 56137 9061 56149 9095
rect 56183 9061 56195 9095
rect 56137 9055 56195 9061
rect 56152 9024 56180 9055
rect 56870 9024 56876 9036
rect 56152 8996 56640 9024
rect 56831 8996 56876 9024
rect 56134 8956 56140 8968
rect 55186 8928 56140 8956
rect 56134 8916 56140 8928
rect 56192 8916 56198 8968
rect 56318 8956 56324 8968
rect 56279 8928 56324 8956
rect 56318 8916 56324 8928
rect 56376 8916 56382 8968
rect 56413 8959 56471 8965
rect 56413 8925 56425 8959
rect 56459 8925 56471 8959
rect 56612 8956 56640 8996
rect 56870 8984 56876 8996
rect 56928 8984 56934 9036
rect 57129 8959 57187 8965
rect 57129 8956 57141 8959
rect 56612 8928 57141 8956
rect 56413 8919 56471 8925
rect 57129 8925 57141 8928
rect 57175 8925 57187 8959
rect 57129 8919 57187 8925
rect 37516 8860 37964 8888
rect 37516 8848 37522 8860
rect 38010 8848 38016 8900
rect 38068 8888 38074 8900
rect 41230 8888 41236 8900
rect 38068 8860 38113 8888
rect 38212 8860 41236 8888
rect 38068 8848 38074 8860
rect 31803 8792 32536 8820
rect 31803 8789 31815 8792
rect 31757 8783 31815 8789
rect 32582 8780 32588 8832
rect 32640 8820 32646 8832
rect 33045 8823 33103 8829
rect 33045 8820 33057 8823
rect 32640 8792 33057 8820
rect 32640 8780 32646 8792
rect 33045 8789 33057 8792
rect 33091 8789 33103 8823
rect 33045 8783 33103 8789
rect 33134 8780 33140 8832
rect 33192 8780 33198 8832
rect 35986 8820 35992 8832
rect 35947 8792 35992 8820
rect 35986 8780 35992 8792
rect 36044 8780 36050 8832
rect 37274 8780 37280 8832
rect 37332 8820 37338 8832
rect 38212 8820 38240 8860
rect 41230 8848 41236 8860
rect 41288 8848 41294 8900
rect 41322 8848 41328 8900
rect 41380 8888 41386 8900
rect 43438 8888 43444 8900
rect 41380 8860 43444 8888
rect 41380 8848 41386 8860
rect 43438 8848 43444 8860
rect 43496 8848 43502 8900
rect 43714 8888 43720 8900
rect 43675 8860 43720 8888
rect 43714 8848 43720 8860
rect 43772 8848 43778 8900
rect 44082 8848 44088 8900
rect 44140 8888 44146 8900
rect 45465 8891 45523 8897
rect 45465 8888 45477 8891
rect 44140 8860 45477 8888
rect 44140 8848 44146 8860
rect 45465 8857 45477 8860
rect 45511 8857 45523 8891
rect 45465 8851 45523 8857
rect 46124 8860 55214 8888
rect 38378 8820 38384 8832
rect 37332 8792 38240 8820
rect 38339 8792 38384 8820
rect 37332 8780 37338 8792
rect 38378 8780 38384 8792
rect 38436 8780 38442 8832
rect 40221 8823 40279 8829
rect 40221 8789 40233 8823
rect 40267 8820 40279 8823
rect 40865 8823 40923 8829
rect 40865 8820 40877 8823
rect 40267 8792 40877 8820
rect 40267 8789 40279 8792
rect 40221 8783 40279 8789
rect 40865 8789 40877 8792
rect 40911 8789 40923 8823
rect 40865 8783 40923 8789
rect 40954 8780 40960 8832
rect 41012 8820 41018 8832
rect 46124 8820 46152 8860
rect 41012 8792 46152 8820
rect 55186 8820 55214 8860
rect 56428 8820 56456 8919
rect 55186 8792 56456 8820
rect 41012 8780 41018 8792
rect 57054 8780 57060 8832
rect 57112 8820 57118 8832
rect 58253 8823 58311 8829
rect 58253 8820 58265 8823
rect 57112 8792 58265 8820
rect 57112 8780 57118 8792
rect 58253 8789 58265 8792
rect 58299 8789 58311 8823
rect 58253 8783 58311 8789
rect 1104 8730 58880 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 58880 8730
rect 1104 8656 58880 8678
rect 13446 8576 13452 8628
rect 13504 8616 13510 8628
rect 14093 8619 14151 8625
rect 14093 8616 14105 8619
rect 13504 8588 14105 8616
rect 13504 8576 13510 8588
rect 14093 8585 14105 8588
rect 14139 8585 14151 8619
rect 14093 8579 14151 8585
rect 14918 8576 14924 8628
rect 14976 8616 14982 8628
rect 16209 8619 16267 8625
rect 16209 8616 16221 8619
rect 14976 8588 16221 8616
rect 14976 8576 14982 8588
rect 16209 8585 16221 8588
rect 16255 8585 16267 8619
rect 16209 8579 16267 8585
rect 16574 8576 16580 8628
rect 16632 8616 16638 8628
rect 17218 8616 17224 8628
rect 16632 8588 17224 8616
rect 16632 8576 16638 8588
rect 17218 8576 17224 8588
rect 17276 8616 17282 8628
rect 17276 8588 17540 8616
rect 17276 8576 17282 8588
rect 15102 8508 15108 8560
rect 15160 8548 15166 8560
rect 17034 8548 17040 8560
rect 15160 8520 15424 8548
rect 16995 8520 17040 8548
rect 15160 8508 15166 8520
rect 1581 8483 1639 8489
rect 1581 8449 1593 8483
rect 1627 8480 1639 8483
rect 10594 8480 10600 8492
rect 1627 8452 10600 8480
rect 1627 8449 1639 8452
rect 1581 8443 1639 8449
rect 10594 8440 10600 8452
rect 10652 8440 10658 8492
rect 13998 8480 14004 8492
rect 13959 8452 14004 8480
rect 13998 8440 14004 8452
rect 14056 8440 14062 8492
rect 15197 8483 15255 8489
rect 15197 8449 15209 8483
rect 15243 8480 15255 8483
rect 15286 8480 15292 8492
rect 15243 8452 15292 8480
rect 15243 8449 15255 8452
rect 15197 8443 15255 8449
rect 15286 8440 15292 8452
rect 15344 8440 15350 8492
rect 15396 8489 15424 8520
rect 17034 8508 17040 8520
rect 17092 8508 17098 8560
rect 17512 8548 17540 8588
rect 19150 8576 19156 8628
rect 19208 8576 19214 8628
rect 19242 8576 19248 8628
rect 19300 8616 19306 8628
rect 19429 8619 19487 8625
rect 19429 8616 19441 8619
rect 19300 8588 19441 8616
rect 19300 8576 19306 8588
rect 19429 8585 19441 8588
rect 19475 8585 19487 8619
rect 19429 8579 19487 8585
rect 19886 8576 19892 8628
rect 19944 8616 19950 8628
rect 22738 8616 22744 8628
rect 19944 8588 22744 8616
rect 19944 8576 19950 8588
rect 22738 8576 22744 8588
rect 22796 8576 22802 8628
rect 23032 8588 23244 8616
rect 17512 8520 17632 8548
rect 15381 8483 15439 8489
rect 15381 8449 15393 8483
rect 15427 8449 15439 8483
rect 15381 8443 15439 8449
rect 15470 8440 15476 8492
rect 15528 8480 15534 8492
rect 16117 8483 16175 8489
rect 16117 8480 16129 8483
rect 15528 8452 16129 8480
rect 15528 8440 15534 8452
rect 16117 8449 16129 8452
rect 16163 8480 16175 8483
rect 16666 8480 16672 8492
rect 16163 8452 16672 8480
rect 16163 8449 16175 8452
rect 16117 8443 16175 8449
rect 16666 8440 16672 8452
rect 16724 8480 16730 8492
rect 16945 8483 17003 8489
rect 16945 8480 16957 8483
rect 16724 8452 16957 8480
rect 16724 8440 16730 8452
rect 16945 8449 16957 8452
rect 16991 8449 17003 8483
rect 16945 8443 17003 8449
rect 17126 8440 17132 8492
rect 17184 8480 17190 8492
rect 17604 8489 17632 8520
rect 17954 8508 17960 8560
rect 18012 8548 18018 8560
rect 19168 8548 19196 8576
rect 23032 8548 23060 8588
rect 18012 8520 19104 8548
rect 19168 8520 23060 8548
rect 23216 8548 23244 8588
rect 23290 8576 23296 8628
rect 23348 8616 23354 8628
rect 23385 8619 23443 8625
rect 23385 8616 23397 8619
rect 23348 8588 23397 8616
rect 23348 8576 23354 8588
rect 23385 8585 23397 8588
rect 23431 8585 23443 8619
rect 23385 8579 23443 8585
rect 23477 8619 23535 8625
rect 23477 8585 23489 8619
rect 23523 8616 23535 8619
rect 23842 8616 23848 8628
rect 23523 8588 23848 8616
rect 23523 8585 23535 8588
rect 23477 8579 23535 8585
rect 23842 8576 23848 8588
rect 23900 8576 23906 8628
rect 25130 8576 25136 8628
rect 25188 8616 25194 8628
rect 25317 8619 25375 8625
rect 25317 8616 25329 8619
rect 25188 8588 25329 8616
rect 25188 8576 25194 8588
rect 25317 8585 25329 8588
rect 25363 8585 25375 8619
rect 25317 8579 25375 8585
rect 28350 8576 28356 8628
rect 28408 8616 28414 8628
rect 28718 8616 28724 8628
rect 28408 8588 28724 8616
rect 28408 8576 28414 8588
rect 28718 8576 28724 8588
rect 28776 8616 28782 8628
rect 31570 8616 31576 8628
rect 28776 8588 31576 8616
rect 28776 8576 28782 8588
rect 31570 8576 31576 8588
rect 31628 8576 31634 8628
rect 33413 8619 33471 8625
rect 33413 8585 33425 8619
rect 33459 8616 33471 8619
rect 34238 8616 34244 8628
rect 33459 8588 34244 8616
rect 33459 8585 33471 8588
rect 33413 8579 33471 8585
rect 34238 8576 34244 8588
rect 34296 8576 34302 8628
rect 35342 8616 35348 8628
rect 34339 8588 35348 8616
rect 23661 8551 23719 8557
rect 23661 8548 23673 8551
rect 23216 8520 23673 8548
rect 18012 8508 18018 8520
rect 17405 8483 17463 8489
rect 17405 8480 17417 8483
rect 17184 8452 17417 8480
rect 17184 8440 17190 8452
rect 17405 8449 17417 8452
rect 17451 8449 17463 8483
rect 17405 8443 17463 8449
rect 17497 8483 17555 8489
rect 17497 8449 17509 8483
rect 17543 8449 17555 8483
rect 17497 8443 17555 8449
rect 17589 8483 17647 8489
rect 17589 8449 17601 8483
rect 17635 8449 17647 8483
rect 17589 8443 17647 8449
rect 1762 8412 1768 8424
rect 1723 8384 1768 8412
rect 1762 8372 1768 8384
rect 1820 8372 1826 8424
rect 17310 8372 17316 8424
rect 17368 8412 17374 8424
rect 17512 8412 17540 8443
rect 17368 8384 17540 8412
rect 17604 8412 17632 8443
rect 17862 8440 17868 8492
rect 17920 8480 17926 8492
rect 19076 8489 19104 8520
rect 23661 8517 23673 8520
rect 23707 8517 23719 8551
rect 29546 8548 29552 8560
rect 23661 8511 23719 8517
rect 24136 8520 29552 8548
rect 24136 8492 24164 8520
rect 29546 8508 29552 8520
rect 29604 8508 29610 8560
rect 30929 8551 30987 8557
rect 30929 8548 30941 8551
rect 29748 8520 30941 8548
rect 18325 8483 18383 8489
rect 18693 8486 18751 8489
rect 18325 8480 18337 8483
rect 17920 8452 18337 8480
rect 17920 8440 17926 8452
rect 18325 8449 18337 8452
rect 18371 8449 18383 8483
rect 18524 8483 18751 8486
rect 18524 8480 18705 8483
rect 18325 8443 18383 8449
rect 18432 8458 18705 8480
rect 18432 8452 18552 8458
rect 18432 8412 18460 8452
rect 18693 8449 18705 8458
rect 18739 8449 18751 8483
rect 18693 8443 18751 8449
rect 19061 8483 19119 8489
rect 19061 8449 19073 8483
rect 19107 8449 19119 8483
rect 19061 8443 19119 8449
rect 19889 8483 19947 8489
rect 19889 8449 19901 8483
rect 19935 8480 19947 8483
rect 20346 8480 20352 8492
rect 19935 8452 20352 8480
rect 19935 8449 19947 8452
rect 19889 8443 19947 8449
rect 19904 8412 19932 8443
rect 20346 8440 20352 8452
rect 20404 8440 20410 8492
rect 22370 8480 22376 8492
rect 22331 8452 22376 8480
rect 22370 8440 22376 8452
rect 22428 8440 22434 8492
rect 23293 8483 23351 8489
rect 23293 8449 23305 8483
rect 23339 8480 23351 8483
rect 24118 8480 24124 8492
rect 23339 8452 23428 8480
rect 24079 8452 24124 8480
rect 23339 8449 23351 8452
rect 23293 8443 23351 8449
rect 17604 8384 18460 8412
rect 19010 8384 19932 8412
rect 17368 8372 17374 8384
rect 19010 8356 19038 8384
rect 19978 8372 19984 8424
rect 20036 8412 20042 8424
rect 22278 8412 22284 8424
rect 20036 8384 22284 8412
rect 20036 8372 20042 8384
rect 22278 8372 22284 8384
rect 22336 8372 22342 8424
rect 13354 8304 13360 8356
rect 13412 8344 13418 8356
rect 15565 8347 15623 8353
rect 15565 8344 15577 8347
rect 13412 8316 15577 8344
rect 13412 8304 13418 8316
rect 15565 8313 15577 8316
rect 15611 8313 15623 8347
rect 17862 8344 17868 8356
rect 15565 8307 15623 8313
rect 17696 8316 17868 8344
rect 15381 8279 15439 8285
rect 15381 8245 15393 8279
rect 15427 8276 15439 8279
rect 15654 8276 15660 8288
rect 15427 8248 15660 8276
rect 15427 8245 15439 8248
rect 15381 8239 15439 8245
rect 15654 8236 15660 8248
rect 15712 8236 15718 8288
rect 17402 8236 17408 8288
rect 17460 8276 17466 8288
rect 17696 8276 17724 8316
rect 17862 8304 17868 8316
rect 17920 8304 17926 8356
rect 18966 8344 18972 8356
rect 18616 8316 18972 8344
rect 18616 8294 18644 8316
rect 18966 8304 18972 8316
rect 19024 8316 19038 8356
rect 19886 8344 19892 8356
rect 19076 8316 19892 8344
rect 19024 8304 19030 8316
rect 18524 8288 18644 8294
rect 19076 8288 19104 8316
rect 19886 8304 19892 8316
rect 19944 8304 19950 8356
rect 20254 8304 20260 8356
rect 20312 8344 20318 8356
rect 23109 8347 23167 8353
rect 23109 8344 23121 8347
rect 20312 8316 23121 8344
rect 20312 8304 20318 8316
rect 23109 8313 23121 8316
rect 23155 8313 23167 8347
rect 23400 8344 23428 8452
rect 24118 8440 24124 8452
rect 24176 8440 24182 8492
rect 27154 8480 27160 8492
rect 27115 8452 27160 8480
rect 27154 8440 27160 8452
rect 27212 8440 27218 8492
rect 27522 8440 27528 8492
rect 27580 8480 27586 8492
rect 28994 8480 29000 8492
rect 27580 8452 29000 8480
rect 27580 8440 27586 8452
rect 28994 8440 29000 8452
rect 29052 8440 29058 8492
rect 29454 8480 29460 8492
rect 29415 8452 29460 8480
rect 29454 8440 29460 8452
rect 29512 8440 29518 8492
rect 23934 8372 23940 8424
rect 23992 8412 23998 8424
rect 25406 8412 25412 8424
rect 23992 8384 25412 8412
rect 23992 8372 23998 8384
rect 25406 8372 25412 8384
rect 25464 8372 25470 8424
rect 25774 8372 25780 8424
rect 25832 8412 25838 8424
rect 27617 8415 27675 8421
rect 27617 8412 27629 8415
rect 25832 8384 27629 8412
rect 25832 8372 25838 8384
rect 27617 8381 27629 8384
rect 27663 8412 27675 8415
rect 27706 8412 27712 8424
rect 27663 8384 27712 8412
rect 27663 8381 27675 8384
rect 27617 8375 27675 8381
rect 27706 8372 27712 8384
rect 27764 8412 27770 8424
rect 28534 8412 28540 8424
rect 27764 8384 28540 8412
rect 27764 8372 27770 8384
rect 28534 8372 28540 8384
rect 28592 8372 28598 8424
rect 29012 8412 29040 8440
rect 29748 8424 29776 8520
rect 30929 8517 30941 8520
rect 30975 8548 30987 8551
rect 31018 8548 31024 8560
rect 30975 8520 31024 8548
rect 30975 8517 30987 8520
rect 30929 8511 30987 8517
rect 31018 8508 31024 8520
rect 31076 8508 31082 8560
rect 33045 8551 33103 8557
rect 33045 8517 33057 8551
rect 33091 8548 33103 8551
rect 33502 8548 33508 8560
rect 33091 8520 33508 8548
rect 33091 8517 33103 8520
rect 33045 8511 33103 8517
rect 33502 8508 33508 8520
rect 33560 8508 33566 8560
rect 34149 8551 34207 8557
rect 34149 8548 34161 8551
rect 34072 8520 34161 8548
rect 30190 8480 30196 8492
rect 30024 8452 30196 8480
rect 29730 8412 29736 8424
rect 29012 8384 29736 8412
rect 29730 8372 29736 8384
rect 29788 8372 29794 8424
rect 24486 8344 24492 8356
rect 23400 8316 24492 8344
rect 23109 8307 23167 8313
rect 24486 8304 24492 8316
rect 24544 8344 24550 8356
rect 30024 8344 30052 8452
rect 30190 8440 30196 8452
rect 30248 8440 30254 8492
rect 30650 8440 30656 8492
rect 30708 8480 30714 8492
rect 31665 8483 31723 8489
rect 31665 8480 31677 8483
rect 30708 8452 31677 8480
rect 30708 8440 30714 8452
rect 31665 8449 31677 8452
rect 31711 8449 31723 8483
rect 32766 8480 32772 8492
rect 32727 8452 32772 8480
rect 31665 8443 31723 8449
rect 32766 8440 32772 8452
rect 32824 8440 32830 8492
rect 32862 8483 32920 8489
rect 32862 8449 32874 8483
rect 32908 8449 32920 8483
rect 33134 8480 33140 8492
rect 33095 8452 33140 8480
rect 32862 8443 32920 8449
rect 30098 8372 30104 8424
rect 30156 8412 30162 8424
rect 31294 8412 31300 8424
rect 30156 8384 30201 8412
rect 31255 8384 31300 8412
rect 30156 8372 30162 8384
rect 31294 8372 31300 8384
rect 31352 8372 31358 8424
rect 31754 8372 31760 8424
rect 31812 8412 31818 8424
rect 32877 8412 32905 8443
rect 33134 8440 33140 8452
rect 33192 8440 33198 8492
rect 33275 8483 33333 8489
rect 33275 8449 33287 8483
rect 33321 8480 33333 8483
rect 33686 8480 33692 8492
rect 33321 8452 33692 8480
rect 33321 8449 33333 8452
rect 33275 8443 33333 8449
rect 33686 8440 33692 8452
rect 33744 8440 33750 8492
rect 33870 8480 33876 8492
rect 33831 8452 33876 8480
rect 33870 8440 33876 8452
rect 33928 8440 33934 8492
rect 33966 8483 34024 8489
rect 33966 8449 33978 8483
rect 34012 8449 34024 8483
rect 33966 8443 34024 8449
rect 33981 8412 34009 8443
rect 31812 8384 34009 8412
rect 31812 8372 31818 8384
rect 24544 8316 30052 8344
rect 24544 8304 24550 8316
rect 30190 8304 30196 8356
rect 30248 8344 30254 8356
rect 30466 8344 30472 8356
rect 30248 8316 30472 8344
rect 30248 8304 30254 8316
rect 30466 8304 30472 8316
rect 30524 8304 30530 8356
rect 31202 8344 31208 8356
rect 31163 8316 31208 8344
rect 31202 8304 31208 8316
rect 31260 8304 31266 8356
rect 33410 8304 33416 8356
rect 33468 8344 33474 8356
rect 34072 8344 34100 8520
rect 34149 8517 34161 8520
rect 34195 8548 34207 8551
rect 34339 8548 34367 8588
rect 35342 8576 35348 8588
rect 35400 8576 35406 8628
rect 40954 8616 40960 8628
rect 37384 8588 40960 8616
rect 37384 8548 37412 8588
rect 40954 8576 40960 8588
rect 41012 8576 41018 8628
rect 44269 8619 44327 8625
rect 44269 8585 44281 8619
rect 44315 8616 44327 8619
rect 46106 8616 46112 8628
rect 44315 8588 46112 8616
rect 44315 8585 44327 8588
rect 44269 8579 44327 8585
rect 46106 8576 46112 8588
rect 46164 8576 46170 8628
rect 46198 8576 46204 8628
rect 46256 8616 46262 8628
rect 56321 8619 56379 8625
rect 56321 8616 56333 8619
rect 46256 8588 56333 8616
rect 46256 8576 46262 8588
rect 56321 8585 56333 8588
rect 56367 8585 56379 8619
rect 56321 8579 56379 8585
rect 37642 8548 37648 8560
rect 34195 8520 34367 8548
rect 35728 8520 37412 8548
rect 37476 8520 37648 8548
rect 34195 8517 34207 8520
rect 34149 8511 34207 8517
rect 34422 8489 34428 8492
rect 34249 8483 34307 8489
rect 34249 8449 34261 8483
rect 34295 8449 34307 8483
rect 34249 8443 34307 8449
rect 34379 8483 34428 8489
rect 34379 8449 34391 8483
rect 34425 8449 34428 8483
rect 34379 8443 34428 8449
rect 33468 8316 34100 8344
rect 33468 8304 33474 8316
rect 17460 8248 17724 8276
rect 17460 8236 17466 8248
rect 18506 8236 18512 8288
rect 18564 8266 18644 8288
rect 18564 8236 18570 8266
rect 19058 8236 19064 8288
rect 19116 8236 19122 8288
rect 19242 8236 19248 8288
rect 19300 8276 19306 8288
rect 20806 8276 20812 8288
rect 19300 8248 20812 8276
rect 19300 8236 19306 8248
rect 20806 8236 20812 8248
rect 20864 8236 20870 8288
rect 22557 8279 22615 8285
rect 22557 8245 22569 8279
rect 22603 8276 22615 8279
rect 23014 8276 23020 8288
rect 22603 8248 23020 8276
rect 22603 8245 22615 8248
rect 22557 8239 22615 8245
rect 23014 8236 23020 8248
rect 23072 8236 23078 8288
rect 23566 8236 23572 8288
rect 23624 8276 23630 8288
rect 27614 8276 27620 8288
rect 23624 8248 27620 8276
rect 23624 8236 23630 8248
rect 27614 8236 27620 8248
rect 27672 8236 27678 8288
rect 29086 8236 29092 8288
rect 29144 8276 29150 8288
rect 31094 8279 31152 8285
rect 31094 8276 31106 8279
rect 29144 8248 31106 8276
rect 29144 8236 29150 8248
rect 31094 8245 31106 8248
rect 31140 8276 31152 8279
rect 31294 8276 31300 8288
rect 31140 8248 31300 8276
rect 31140 8245 31152 8248
rect 31094 8239 31152 8245
rect 31294 8236 31300 8248
rect 31352 8236 31358 8288
rect 33962 8236 33968 8288
rect 34020 8276 34026 8288
rect 34256 8276 34284 8443
rect 34422 8440 34428 8443
rect 34480 8440 34486 8492
rect 35728 8480 35756 8520
rect 35894 8480 35900 8492
rect 35636 8452 35756 8480
rect 35855 8452 35900 8480
rect 35636 8421 35664 8452
rect 35894 8440 35900 8452
rect 35952 8440 35958 8492
rect 36722 8480 36728 8492
rect 36683 8452 36728 8480
rect 36722 8440 36728 8452
rect 36780 8440 36786 8492
rect 37274 8480 37280 8492
rect 37016 8452 37280 8480
rect 35345 8415 35403 8421
rect 35345 8412 35357 8415
rect 34532 8384 35357 8412
rect 34532 8353 34560 8384
rect 35345 8381 35357 8384
rect 35391 8381 35403 8415
rect 35345 8375 35403 8381
rect 35621 8415 35679 8421
rect 35621 8381 35633 8415
rect 35667 8381 35679 8415
rect 35802 8412 35808 8424
rect 35763 8384 35808 8412
rect 35621 8375 35679 8381
rect 35802 8372 35808 8384
rect 35860 8372 35866 8424
rect 36541 8415 36599 8421
rect 36541 8381 36553 8415
rect 36587 8412 36599 8415
rect 37016 8412 37044 8452
rect 37274 8440 37280 8452
rect 37332 8440 37338 8492
rect 37476 8489 37504 8520
rect 37642 8508 37648 8520
rect 37700 8508 37706 8560
rect 39942 8548 39948 8560
rect 39132 8520 39948 8548
rect 37461 8483 37519 8489
rect 37461 8449 37473 8483
rect 37507 8449 37519 8483
rect 37461 8443 37519 8449
rect 37550 8440 37556 8492
rect 37608 8480 37614 8492
rect 37737 8483 37795 8489
rect 37608 8452 37653 8480
rect 37608 8440 37614 8452
rect 37737 8449 37749 8483
rect 37783 8449 37795 8483
rect 37737 8443 37795 8449
rect 36587 8384 37044 8412
rect 36587 8381 36599 8384
rect 36541 8375 36599 8381
rect 37090 8372 37096 8424
rect 37148 8412 37154 8424
rect 37752 8412 37780 8443
rect 39132 8424 39160 8520
rect 39942 8508 39948 8520
rect 40000 8548 40006 8560
rect 45186 8548 45192 8560
rect 40000 8520 45192 8548
rect 40000 8508 40006 8520
rect 45186 8508 45192 8520
rect 45244 8508 45250 8560
rect 53098 8548 53104 8560
rect 45296 8520 53104 8548
rect 39206 8440 39212 8492
rect 39264 8480 39270 8492
rect 39373 8483 39431 8489
rect 39373 8480 39385 8483
rect 39264 8452 39385 8480
rect 39264 8440 39270 8452
rect 39373 8449 39385 8452
rect 39419 8449 39431 8483
rect 39373 8443 39431 8449
rect 42889 8483 42947 8489
rect 42889 8449 42901 8483
rect 42935 8480 42947 8483
rect 42978 8480 42984 8492
rect 42935 8452 42984 8480
rect 42935 8449 42947 8452
rect 42889 8443 42947 8449
rect 42978 8440 42984 8452
rect 43036 8440 43042 8492
rect 44266 8440 44272 8492
rect 44324 8480 44330 8492
rect 44453 8483 44511 8489
rect 44453 8480 44465 8483
rect 44324 8452 44465 8480
rect 44324 8440 44330 8452
rect 44453 8449 44465 8452
rect 44499 8449 44511 8483
rect 44453 8443 44511 8449
rect 44542 8440 44548 8492
rect 44600 8480 44606 8492
rect 44729 8483 44787 8489
rect 44600 8452 44645 8480
rect 44600 8440 44606 8452
rect 44729 8449 44741 8483
rect 44775 8449 44787 8483
rect 44729 8443 44787 8449
rect 37148 8384 37780 8412
rect 37921 8415 37979 8421
rect 37148 8372 37154 8384
rect 37921 8381 37933 8415
rect 37967 8412 37979 8415
rect 38010 8412 38016 8424
rect 37967 8384 38016 8412
rect 37967 8381 37979 8384
rect 37921 8375 37979 8381
rect 34517 8347 34575 8353
rect 34517 8313 34529 8347
rect 34563 8313 34575 8347
rect 37936 8344 37964 8375
rect 38010 8372 38016 8384
rect 38068 8372 38074 8424
rect 39114 8412 39120 8424
rect 39075 8384 39120 8412
rect 39114 8372 39120 8384
rect 39172 8372 39178 8424
rect 42518 8372 42524 8424
rect 42576 8412 42582 8424
rect 43165 8415 43223 8421
rect 43165 8412 43177 8415
rect 42576 8384 43177 8412
rect 42576 8372 42582 8384
rect 43165 8381 43177 8384
rect 43211 8381 43223 8415
rect 43165 8375 43223 8381
rect 43898 8372 43904 8424
rect 43956 8412 43962 8424
rect 44744 8412 44772 8443
rect 44818 8440 44824 8492
rect 44876 8480 44882 8492
rect 45296 8489 45324 8520
rect 53098 8508 53104 8520
rect 53156 8508 53162 8560
rect 57330 8548 57336 8560
rect 57291 8520 57336 8548
rect 57330 8508 57336 8520
rect 57388 8508 57394 8560
rect 45281 8483 45339 8489
rect 44876 8452 44921 8480
rect 44876 8440 44882 8452
rect 45281 8449 45293 8483
rect 45327 8449 45339 8483
rect 46382 8480 46388 8492
rect 46343 8452 46388 8480
rect 45281 8443 45339 8449
rect 46382 8440 46388 8452
rect 46440 8440 46446 8492
rect 56226 8480 56232 8492
rect 56187 8452 56232 8480
rect 56226 8440 56232 8452
rect 56284 8440 56290 8492
rect 57054 8480 57060 8492
rect 57015 8452 57060 8480
rect 57054 8440 57060 8452
rect 57112 8440 57118 8492
rect 45370 8412 45376 8424
rect 43956 8384 45376 8412
rect 43956 8372 43962 8384
rect 45370 8372 45376 8384
rect 45428 8372 45434 8424
rect 45462 8372 45468 8424
rect 45520 8412 45526 8424
rect 46566 8412 46572 8424
rect 45520 8384 45565 8412
rect 46527 8384 46572 8412
rect 45520 8372 45526 8384
rect 46566 8372 46572 8384
rect 46624 8372 46630 8424
rect 34517 8307 34575 8313
rect 36745 8316 37964 8344
rect 40497 8347 40555 8353
rect 34020 8248 34284 8276
rect 34020 8236 34026 8248
rect 34422 8236 34428 8288
rect 34480 8276 34486 8288
rect 36745 8276 36773 8316
rect 40497 8313 40509 8347
rect 40543 8344 40555 8347
rect 40862 8344 40868 8356
rect 40543 8316 40868 8344
rect 40543 8313 40555 8316
rect 40497 8307 40555 8313
rect 40862 8304 40868 8316
rect 40920 8344 40926 8356
rect 56502 8344 56508 8356
rect 40920 8316 56508 8344
rect 40920 8304 40926 8316
rect 56502 8304 56508 8316
rect 56560 8304 56566 8356
rect 36906 8276 36912 8288
rect 34480 8248 36773 8276
rect 36867 8248 36912 8276
rect 34480 8236 34486 8248
rect 36906 8236 36912 8248
rect 36964 8236 36970 8288
rect 38838 8236 38844 8288
rect 38896 8276 38902 8288
rect 43162 8276 43168 8288
rect 38896 8248 43168 8276
rect 38896 8236 38902 8248
rect 43162 8236 43168 8248
rect 43220 8236 43226 8288
rect 43438 8236 43444 8288
rect 43496 8276 43502 8288
rect 44818 8276 44824 8288
rect 43496 8248 44824 8276
rect 43496 8236 43502 8248
rect 44818 8236 44824 8248
rect 44876 8276 44882 8288
rect 45462 8276 45468 8288
rect 44876 8248 45468 8276
rect 44876 8236 44882 8248
rect 45462 8236 45468 8248
rect 45520 8236 45526 8288
rect 55490 8236 55496 8288
rect 55548 8276 55554 8288
rect 56962 8276 56968 8288
rect 55548 8248 56968 8276
rect 55548 8236 55554 8248
rect 56962 8236 56968 8248
rect 57020 8236 57026 8288
rect 1104 8186 58880 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 58880 8186
rect 1104 8112 58880 8134
rect 2682 8032 2688 8084
rect 2740 8072 2746 8084
rect 2740 8032 2774 8072
rect 10042 8032 10048 8084
rect 10100 8072 10106 8084
rect 26234 8072 26240 8084
rect 10100 8044 26240 8072
rect 10100 8032 10106 8044
rect 26234 8032 26240 8044
rect 26292 8032 26298 8084
rect 32398 8072 32404 8084
rect 26344 8044 32404 8072
rect 2746 7936 2774 8032
rect 12710 7964 12716 8016
rect 12768 8004 12774 8016
rect 12805 8007 12863 8013
rect 12805 8004 12817 8007
rect 12768 7976 12817 8004
rect 12768 7964 12774 7976
rect 12805 7973 12817 7976
rect 12851 7973 12863 8007
rect 12805 7967 12863 7973
rect 13998 7964 14004 8016
rect 14056 8004 14062 8016
rect 15194 8004 15200 8016
rect 14056 7976 15200 8004
rect 14056 7964 14062 7976
rect 15194 7964 15200 7976
rect 15252 8004 15258 8016
rect 16482 8004 16488 8016
rect 15252 7976 16488 8004
rect 15252 7964 15258 7976
rect 16482 7964 16488 7976
rect 16540 7964 16546 8016
rect 16666 7964 16672 8016
rect 16724 8004 16730 8016
rect 17494 8004 17500 8016
rect 16724 7976 17500 8004
rect 16724 7964 16730 7976
rect 17494 7964 17500 7976
rect 17552 7964 17558 8016
rect 17586 7964 17592 8016
rect 17644 8004 17650 8016
rect 17770 8004 17776 8016
rect 17644 7976 17776 8004
rect 17644 7964 17650 7976
rect 17770 7964 17776 7976
rect 17828 7964 17834 8016
rect 18690 7964 18696 8016
rect 18748 8004 18754 8016
rect 19150 8004 19156 8016
rect 18748 7976 19156 8004
rect 18748 7964 18754 7976
rect 19150 7964 19156 7976
rect 19208 7964 19214 8016
rect 20806 8004 20812 8016
rect 20767 7976 20812 8004
rect 20806 7964 20812 7976
rect 20864 7964 20870 8016
rect 26145 8007 26203 8013
rect 26145 8004 26157 8007
rect 22066 7976 26157 8004
rect 11149 7939 11207 7945
rect 11149 7936 11161 7939
rect 2746 7908 11161 7936
rect 1578 7868 1584 7880
rect 1539 7840 1584 7868
rect 1578 7828 1584 7840
rect 1636 7828 1642 7880
rect 5994 7828 6000 7880
rect 6052 7868 6058 7880
rect 7837 7871 7895 7877
rect 7837 7868 7849 7871
rect 6052 7840 7849 7868
rect 6052 7828 6058 7840
rect 7837 7837 7849 7840
rect 7883 7837 7895 7871
rect 7837 7831 7895 7837
rect 7926 7828 7932 7880
rect 7984 7868 7990 7880
rect 8113 7871 8171 7877
rect 7984 7840 8029 7868
rect 7984 7828 7990 7840
rect 8113 7837 8125 7871
rect 8159 7868 8171 7871
rect 8754 7868 8760 7880
rect 8159 7840 8760 7868
rect 8159 7837 8171 7840
rect 8113 7831 8171 7837
rect 8754 7828 8760 7840
rect 8812 7828 8818 7880
rect 9953 7871 10011 7877
rect 9953 7837 9965 7871
rect 9999 7868 10011 7871
rect 10042 7868 10048 7880
rect 9999 7840 10048 7868
rect 9999 7837 10011 7840
rect 9953 7831 10011 7837
rect 10042 7828 10048 7840
rect 10100 7828 10106 7880
rect 10244 7877 10272 7908
rect 11149 7905 11161 7908
rect 11195 7936 11207 7939
rect 16298 7936 16304 7948
rect 11195 7908 16304 7936
rect 11195 7905 11207 7908
rect 11149 7899 11207 7905
rect 16298 7896 16304 7908
rect 16356 7896 16362 7948
rect 17310 7936 17316 7948
rect 17052 7908 17316 7936
rect 10229 7871 10287 7877
rect 10229 7837 10241 7871
rect 10275 7837 10287 7871
rect 10229 7831 10287 7837
rect 10873 7871 10931 7877
rect 10873 7837 10885 7871
rect 10919 7868 10931 7871
rect 15010 7868 15016 7880
rect 10919 7840 15016 7868
rect 10919 7837 10931 7840
rect 10873 7831 10931 7837
rect 15010 7828 15016 7840
rect 15068 7828 15074 7880
rect 15194 7868 15200 7880
rect 15155 7840 15200 7868
rect 15194 7828 15200 7840
rect 15252 7828 15258 7880
rect 15470 7868 15476 7880
rect 15431 7840 15476 7868
rect 15470 7828 15476 7840
rect 15528 7828 15534 7880
rect 16022 7828 16028 7880
rect 16080 7868 16086 7880
rect 17052 7877 17080 7908
rect 17310 7896 17316 7908
rect 17368 7896 17374 7948
rect 19426 7936 19432 7948
rect 19387 7908 19432 7936
rect 19426 7896 19432 7908
rect 19484 7896 19490 7948
rect 20714 7896 20720 7948
rect 20772 7936 20778 7948
rect 22066 7936 22094 7976
rect 26145 7973 26157 7976
rect 26191 7973 26203 8007
rect 26145 7967 26203 7973
rect 20772 7908 22094 7936
rect 23293 7939 23351 7945
rect 20772 7896 20778 7908
rect 23293 7905 23305 7939
rect 23339 7936 23351 7939
rect 23750 7936 23756 7948
rect 23339 7908 23756 7936
rect 23339 7905 23351 7908
rect 23293 7899 23351 7905
rect 23750 7896 23756 7908
rect 23808 7896 23814 7948
rect 26344 7936 26372 8044
rect 32398 8032 32404 8044
rect 32456 8072 32462 8084
rect 33962 8072 33968 8084
rect 32456 8044 33968 8072
rect 32456 8032 32462 8044
rect 33962 8032 33968 8044
rect 34020 8032 34026 8084
rect 34149 8075 34207 8081
rect 34149 8041 34161 8075
rect 34195 8072 34207 8075
rect 35802 8072 35808 8084
rect 34195 8044 35808 8072
rect 34195 8041 34207 8044
rect 34149 8035 34207 8041
rect 35802 8032 35808 8044
rect 35860 8032 35866 8084
rect 37734 8072 37740 8084
rect 36280 8044 37740 8072
rect 27338 7964 27344 8016
rect 27396 8004 27402 8016
rect 30466 8004 30472 8016
rect 27396 7976 30472 8004
rect 27396 7964 27402 7976
rect 30466 7964 30472 7976
rect 30524 7964 30530 8016
rect 30926 8004 30932 8016
rect 30887 7976 30932 8004
rect 30926 7964 30932 7976
rect 30984 7964 30990 8016
rect 31294 7964 31300 8016
rect 31352 8004 31358 8016
rect 31481 8007 31539 8013
rect 31481 8004 31493 8007
rect 31352 7976 31493 8004
rect 31352 7964 31358 7976
rect 31481 7973 31493 7976
rect 31527 7973 31539 8007
rect 31481 7967 31539 7973
rect 31662 7964 31668 8016
rect 31720 8004 31726 8016
rect 31846 8004 31852 8016
rect 31720 7976 31852 8004
rect 31720 7964 31726 7976
rect 31846 7964 31852 7976
rect 31904 7964 31910 8016
rect 32490 7964 32496 8016
rect 32548 8004 32554 8016
rect 32585 8007 32643 8013
rect 32585 8004 32597 8007
rect 32548 7976 32597 8004
rect 32548 7964 32554 7976
rect 32585 7973 32597 7976
rect 32631 7973 32643 8007
rect 32585 7967 32643 7973
rect 33134 7964 33140 8016
rect 33192 8004 33198 8016
rect 33318 8004 33324 8016
rect 33192 7976 33324 8004
rect 33192 7964 33198 7976
rect 33318 7964 33324 7976
rect 33376 7964 33382 8016
rect 34606 7964 34612 8016
rect 34664 8004 34670 8016
rect 35253 8007 35311 8013
rect 35253 8004 35265 8007
rect 34664 7976 35265 8004
rect 34664 7964 34670 7976
rect 35253 7973 35265 7976
rect 35299 8004 35311 8007
rect 35618 8004 35624 8016
rect 35299 7976 35624 8004
rect 35299 7973 35311 7976
rect 35253 7967 35311 7973
rect 35618 7964 35624 7976
rect 35676 7964 35682 8016
rect 35710 7964 35716 8016
rect 35768 8004 35774 8016
rect 36280 8004 36308 8044
rect 37734 8032 37740 8044
rect 37792 8032 37798 8084
rect 38657 8075 38715 8081
rect 38657 8041 38669 8075
rect 38703 8072 38715 8075
rect 39206 8072 39212 8084
rect 38703 8044 39212 8072
rect 38703 8041 38715 8044
rect 38657 8035 38715 8041
rect 39206 8032 39212 8044
rect 39264 8032 39270 8084
rect 42889 8075 42947 8081
rect 42889 8041 42901 8075
rect 42935 8072 42947 8075
rect 43714 8072 43720 8084
rect 42935 8044 43720 8072
rect 42935 8041 42947 8044
rect 42889 8035 42947 8041
rect 43714 8032 43720 8044
rect 43772 8032 43778 8084
rect 45373 8075 45431 8081
rect 45373 8041 45385 8075
rect 45419 8072 45431 8075
rect 46382 8072 46388 8084
rect 45419 8044 46388 8072
rect 45419 8041 45431 8044
rect 45373 8035 45431 8041
rect 46382 8032 46388 8044
rect 46440 8032 46446 8084
rect 57790 8072 57796 8084
rect 56060 8044 57796 8072
rect 35768 7976 36308 8004
rect 35768 7964 35774 7976
rect 37274 7964 37280 8016
rect 37332 8004 37338 8016
rect 38838 8004 38844 8016
rect 37332 7976 38844 8004
rect 37332 7964 37338 7976
rect 38838 7964 38844 7976
rect 38896 7964 38902 8016
rect 38930 7964 38936 8016
rect 38988 8004 38994 8016
rect 38988 7976 39033 8004
rect 38988 7964 38994 7976
rect 43162 7964 43168 8016
rect 43220 8004 43226 8016
rect 55950 8004 55956 8016
rect 43220 7976 55956 8004
rect 43220 7964 43226 7976
rect 55950 7964 55956 7976
rect 56008 7964 56014 8016
rect 28718 7936 28724 7948
rect 24964 7908 26372 7936
rect 28679 7908 28724 7936
rect 24964 7880 24992 7908
rect 28718 7896 28724 7908
rect 28776 7896 28782 7948
rect 29822 7936 29828 7948
rect 29783 7908 29828 7936
rect 29822 7896 29828 7908
rect 29880 7896 29886 7948
rect 30116 7908 36400 7936
rect 16485 7871 16543 7877
rect 16485 7868 16497 7871
rect 16080 7840 16497 7868
rect 16080 7828 16086 7840
rect 16485 7837 16497 7840
rect 16531 7837 16543 7871
rect 16485 7831 16543 7837
rect 17037 7871 17095 7877
rect 17037 7837 17049 7871
rect 17083 7837 17095 7871
rect 17218 7868 17224 7880
rect 17179 7840 17224 7868
rect 17037 7831 17095 7837
rect 17218 7828 17224 7840
rect 17276 7828 17282 7880
rect 17402 7828 17408 7880
rect 17460 7868 17466 7880
rect 17954 7868 17960 7880
rect 17460 7840 17960 7868
rect 17460 7828 17466 7840
rect 17954 7828 17960 7840
rect 18012 7868 18018 7880
rect 19058 7868 19064 7880
rect 18012 7840 19064 7868
rect 18012 7828 18018 7840
rect 19058 7828 19064 7840
rect 19116 7828 19122 7880
rect 19628 7840 19840 7868
rect 1854 7800 1860 7812
rect 1815 7772 1860 7800
rect 1854 7760 1860 7772
rect 1912 7760 1918 7812
rect 8570 7800 8576 7812
rect 8531 7772 8576 7800
rect 8570 7760 8576 7772
rect 8628 7760 8634 7812
rect 9766 7800 9772 7812
rect 9727 7772 9772 7800
rect 9766 7760 9772 7772
rect 9824 7760 9830 7812
rect 12434 7760 12440 7812
rect 12492 7800 12498 7812
rect 12529 7803 12587 7809
rect 12529 7800 12541 7803
rect 12492 7772 12541 7800
rect 12492 7760 12498 7772
rect 12529 7769 12541 7772
rect 12575 7769 12587 7803
rect 12529 7763 12587 7769
rect 15657 7803 15715 7809
rect 15657 7769 15669 7803
rect 15703 7800 15715 7803
rect 15746 7800 15752 7812
rect 15703 7772 15752 7800
rect 15703 7769 15715 7772
rect 15657 7763 15715 7769
rect 15746 7760 15752 7772
rect 15804 7760 15810 7812
rect 15933 7803 15991 7809
rect 15933 7769 15945 7803
rect 15979 7800 15991 7803
rect 19628 7800 19656 7840
rect 15979 7772 19656 7800
rect 19696 7803 19754 7809
rect 15979 7769 15991 7772
rect 15933 7763 15991 7769
rect 19696 7769 19708 7803
rect 19742 7769 19754 7803
rect 19812 7800 19840 7840
rect 19978 7828 19984 7880
rect 20036 7868 20042 7880
rect 24026 7868 24032 7880
rect 20036 7840 24032 7868
rect 20036 7828 20042 7840
rect 24026 7828 24032 7840
rect 24084 7828 24090 7880
rect 24946 7868 24952 7880
rect 24907 7840 24952 7868
rect 24946 7828 24952 7840
rect 25004 7828 25010 7880
rect 28258 7828 28264 7880
rect 28316 7868 28322 7880
rect 28353 7871 28411 7877
rect 28353 7868 28365 7871
rect 28316 7840 28365 7868
rect 28316 7828 28322 7840
rect 28353 7837 28365 7840
rect 28399 7837 28411 7871
rect 29454 7868 29460 7880
rect 28353 7831 28411 7837
rect 28460 7840 29460 7868
rect 28460 7800 28488 7840
rect 29454 7828 29460 7840
rect 29512 7828 29518 7880
rect 30006 7868 30012 7880
rect 29967 7840 30012 7868
rect 30006 7828 30012 7840
rect 30064 7828 30070 7880
rect 30116 7877 30144 7908
rect 30101 7871 30159 7877
rect 30101 7837 30113 7871
rect 30147 7837 30159 7871
rect 30101 7831 30159 7837
rect 31018 7828 31024 7880
rect 31076 7868 31082 7880
rect 31389 7871 31447 7877
rect 31389 7868 31401 7871
rect 31076 7840 31401 7868
rect 31076 7828 31082 7840
rect 31389 7837 31401 7840
rect 31435 7837 31447 7871
rect 31389 7831 31447 7837
rect 31665 7871 31723 7877
rect 31665 7837 31677 7871
rect 31711 7837 31723 7871
rect 31665 7831 31723 7837
rect 19812 7772 28488 7800
rect 19696 7763 19754 7769
rect 9950 7692 9956 7744
rect 10008 7732 10014 7744
rect 10137 7735 10195 7741
rect 10137 7732 10149 7735
rect 10008 7704 10149 7732
rect 10008 7692 10014 7704
rect 10137 7701 10149 7704
rect 10183 7701 10195 7735
rect 10137 7695 10195 7701
rect 12989 7735 13047 7741
rect 12989 7701 13001 7735
rect 13035 7732 13047 7735
rect 15286 7732 15292 7744
rect 13035 7704 15292 7732
rect 13035 7701 13047 7704
rect 12989 7695 13047 7701
rect 15286 7692 15292 7704
rect 15344 7692 15350 7744
rect 15565 7735 15623 7741
rect 15565 7701 15577 7735
rect 15611 7732 15623 7735
rect 16022 7732 16028 7744
rect 15611 7704 16028 7732
rect 15611 7701 15623 7704
rect 15565 7695 15623 7701
rect 16022 7692 16028 7704
rect 16080 7692 16086 7744
rect 16485 7735 16543 7741
rect 16485 7701 16497 7735
rect 16531 7732 16543 7735
rect 16758 7732 16764 7744
rect 16531 7704 16764 7732
rect 16531 7701 16543 7704
rect 16485 7695 16543 7701
rect 16758 7692 16764 7704
rect 16816 7692 16822 7744
rect 17954 7692 17960 7744
rect 18012 7732 18018 7744
rect 18506 7732 18512 7744
rect 18012 7704 18512 7732
rect 18012 7692 18018 7704
rect 18506 7692 18512 7704
rect 18564 7692 18570 7744
rect 19334 7692 19340 7744
rect 19392 7732 19398 7744
rect 19720 7732 19748 7763
rect 28718 7760 28724 7812
rect 28776 7800 28782 7812
rect 30469 7803 30527 7809
rect 30469 7800 30481 7803
rect 28776 7772 30481 7800
rect 28776 7760 28782 7772
rect 30469 7769 30481 7772
rect 30515 7769 30527 7803
rect 30469 7763 30527 7769
rect 31202 7760 31208 7812
rect 31260 7800 31266 7812
rect 31680 7800 31708 7831
rect 32214 7828 32220 7880
rect 32272 7868 32278 7880
rect 32769 7871 32827 7877
rect 32769 7868 32781 7871
rect 32272 7840 32781 7868
rect 32272 7828 32278 7840
rect 32769 7837 32781 7840
rect 32815 7837 32827 7871
rect 33594 7868 33600 7880
rect 32769 7831 32827 7837
rect 32876 7840 33600 7868
rect 31260 7772 31708 7800
rect 31260 7760 31266 7772
rect 19392 7704 19748 7732
rect 19392 7692 19398 7704
rect 20162 7692 20168 7744
rect 20220 7732 20226 7744
rect 20346 7732 20352 7744
rect 20220 7704 20352 7732
rect 20220 7692 20226 7704
rect 20346 7692 20352 7704
rect 20404 7732 20410 7744
rect 21450 7732 21456 7744
rect 20404 7704 21456 7732
rect 20404 7692 20410 7704
rect 21450 7692 21456 7704
rect 21508 7692 21514 7744
rect 22278 7692 22284 7744
rect 22336 7732 22342 7744
rect 22649 7735 22707 7741
rect 22649 7732 22661 7735
rect 22336 7704 22661 7732
rect 22336 7692 22342 7704
rect 22649 7701 22661 7704
rect 22695 7701 22707 7735
rect 23014 7732 23020 7744
rect 22975 7704 23020 7732
rect 22649 7695 22707 7701
rect 23014 7692 23020 7704
rect 23072 7692 23078 7744
rect 23106 7692 23112 7744
rect 23164 7732 23170 7744
rect 23164 7704 23209 7732
rect 23164 7692 23170 7704
rect 23474 7692 23480 7744
rect 23532 7732 23538 7744
rect 31110 7732 31116 7744
rect 23532 7704 31116 7732
rect 23532 7692 23538 7704
rect 31110 7692 31116 7704
rect 31168 7692 31174 7744
rect 31846 7732 31852 7744
rect 31807 7704 31852 7732
rect 31846 7692 31852 7704
rect 31904 7692 31910 7744
rect 32876 7741 32904 7840
rect 33594 7828 33600 7840
rect 33652 7828 33658 7880
rect 34146 7868 34152 7880
rect 34107 7840 34152 7868
rect 34146 7828 34152 7840
rect 34204 7828 34210 7880
rect 34333 7871 34391 7877
rect 34333 7837 34345 7871
rect 34379 7837 34391 7871
rect 34333 7831 34391 7837
rect 33134 7800 33140 7812
rect 33095 7772 33140 7800
rect 33134 7760 33140 7772
rect 33192 7760 33198 7812
rect 34348 7800 34376 7831
rect 35158 7828 35164 7880
rect 35216 7868 35222 7880
rect 36265 7871 36323 7877
rect 36265 7868 36277 7871
rect 35216 7840 36277 7868
rect 35216 7828 35222 7840
rect 36265 7837 36277 7840
rect 36311 7837 36323 7871
rect 36265 7831 36323 7837
rect 34164 7772 34376 7800
rect 34164 7744 34192 7772
rect 34698 7760 34704 7812
rect 34756 7800 34762 7812
rect 34977 7803 35035 7809
rect 34977 7800 34989 7803
rect 34756 7772 34989 7800
rect 34756 7760 34762 7772
rect 34977 7769 34989 7772
rect 35023 7769 35035 7803
rect 36372 7800 36400 7908
rect 38378 7896 38384 7948
rect 38436 7936 38442 7948
rect 38654 7936 38660 7948
rect 38436 7908 38660 7936
rect 38436 7896 38442 7908
rect 38654 7896 38660 7908
rect 38712 7896 38718 7948
rect 39025 7939 39083 7945
rect 39025 7905 39037 7939
rect 39071 7936 39083 7939
rect 39390 7936 39396 7948
rect 39071 7908 39396 7936
rect 39071 7905 39083 7908
rect 39025 7899 39083 7905
rect 39390 7896 39396 7908
rect 39448 7896 39454 7948
rect 39666 7896 39672 7948
rect 39724 7936 39730 7948
rect 46566 7936 46572 7948
rect 39724 7908 46572 7936
rect 39724 7896 39730 7908
rect 36532 7871 36590 7877
rect 36532 7837 36544 7871
rect 36578 7868 36590 7871
rect 36906 7868 36912 7880
rect 36578 7840 36912 7868
rect 36578 7837 36590 7840
rect 36532 7831 36590 7837
rect 36906 7828 36912 7840
rect 36964 7828 36970 7880
rect 38850 7871 38908 7877
rect 38850 7868 38862 7871
rect 38847 7846 38862 7868
rect 38654 7800 38660 7812
rect 36372 7772 38660 7800
rect 34977 7763 35035 7769
rect 38654 7760 38660 7772
rect 38712 7760 38718 7812
rect 38829 7794 38835 7846
rect 38896 7837 38908 7871
rect 38887 7831 38908 7837
rect 39117 7871 39175 7877
rect 39117 7837 39129 7871
rect 39163 7868 39175 7871
rect 39206 7868 39212 7880
rect 39163 7840 39212 7868
rect 39163 7837 39175 7840
rect 39117 7831 39175 7837
rect 38887 7794 38893 7831
rect 39206 7828 39212 7840
rect 39264 7828 39270 7880
rect 39301 7871 39359 7877
rect 39301 7837 39313 7871
rect 39347 7868 39359 7871
rect 40034 7868 40040 7880
rect 39347 7840 40040 7868
rect 39347 7837 39359 7840
rect 39301 7831 39359 7837
rect 40034 7828 40040 7840
rect 40092 7828 40098 7880
rect 42518 7828 42524 7880
rect 42576 7868 42582 7880
rect 42797 7871 42855 7877
rect 42797 7868 42809 7871
rect 42576 7840 42809 7868
rect 42576 7828 42582 7840
rect 42797 7837 42809 7840
rect 42843 7837 42855 7871
rect 42797 7831 42855 7837
rect 43438 7828 43444 7880
rect 43496 7868 43502 7880
rect 43717 7871 43775 7877
rect 43717 7868 43729 7871
rect 43496 7840 43729 7868
rect 43496 7828 43502 7840
rect 43717 7837 43729 7840
rect 43763 7837 43775 7871
rect 43990 7868 43996 7880
rect 43951 7840 43996 7868
rect 43717 7831 43775 7837
rect 43990 7828 43996 7840
rect 44048 7828 44054 7880
rect 44174 7828 44180 7880
rect 44232 7868 44238 7880
rect 45278 7868 45284 7880
rect 44232 7840 45284 7868
rect 44232 7828 44238 7840
rect 45278 7828 45284 7840
rect 45336 7828 45342 7880
rect 45370 7828 45376 7880
rect 45428 7868 45434 7880
rect 46308 7877 46336 7908
rect 46566 7896 46572 7908
rect 46624 7896 46630 7948
rect 46658 7896 46664 7948
rect 46716 7936 46722 7948
rect 56060 7936 56088 8044
rect 57790 8032 57796 8044
rect 57848 8072 57854 8084
rect 58253 8075 58311 8081
rect 58253 8072 58265 8075
rect 57848 8044 58265 8072
rect 57848 8032 57854 8044
rect 58253 8041 58265 8044
rect 58299 8041 58311 8075
rect 58253 8035 58311 8041
rect 56137 8007 56195 8013
rect 56137 7973 56149 8007
rect 56183 7973 56195 8007
rect 56137 7967 56195 7973
rect 46716 7908 46761 7936
rect 55692 7908 56088 7936
rect 56152 7936 56180 7967
rect 56870 7936 56876 7948
rect 56152 7908 56640 7936
rect 56831 7908 56876 7936
rect 46716 7896 46722 7908
rect 45557 7871 45615 7877
rect 45557 7868 45569 7871
rect 45428 7840 45569 7868
rect 45428 7828 45434 7840
rect 45557 7837 45569 7840
rect 45603 7837 45615 7871
rect 45557 7831 45615 7837
rect 46293 7871 46351 7877
rect 46293 7837 46305 7871
rect 46339 7837 46351 7871
rect 55490 7868 55496 7880
rect 55451 7840 55496 7868
rect 46293 7831 46351 7837
rect 55490 7828 55496 7840
rect 55548 7828 55554 7880
rect 55692 7877 55720 7908
rect 55677 7871 55735 7877
rect 55677 7837 55689 7871
rect 55723 7837 55735 7871
rect 55677 7831 55735 7837
rect 55766 7828 55772 7880
rect 55824 7868 55830 7880
rect 56413 7871 56471 7877
rect 56413 7868 56425 7871
rect 55824 7840 56425 7868
rect 55824 7828 55830 7840
rect 56413 7837 56425 7840
rect 56459 7837 56471 7871
rect 56612 7868 56640 7908
rect 56870 7896 56876 7908
rect 56928 7896 56934 7948
rect 57129 7871 57187 7877
rect 57129 7868 57141 7871
rect 56612 7840 57141 7868
rect 56413 7831 56471 7837
rect 57129 7837 57141 7840
rect 57175 7837 57187 7871
rect 57129 7831 57187 7837
rect 43898 7800 43904 7812
rect 43859 7772 43904 7800
rect 43898 7760 43904 7772
rect 43956 7760 43962 7812
rect 44450 7800 44456 7812
rect 44411 7772 44456 7800
rect 44450 7760 44456 7772
rect 44508 7760 44514 7812
rect 45465 7803 45523 7809
rect 45465 7769 45477 7803
rect 45511 7800 45523 7803
rect 46750 7800 46756 7812
rect 45511 7772 46756 7800
rect 45511 7769 45523 7772
rect 45465 7763 45523 7769
rect 46750 7760 46756 7772
rect 46808 7760 46814 7812
rect 56134 7800 56140 7812
rect 56095 7772 56140 7800
rect 56134 7760 56140 7772
rect 56192 7760 56198 7812
rect 32861 7735 32919 7741
rect 32861 7701 32873 7735
rect 32907 7701 32919 7735
rect 32861 7695 32919 7701
rect 32953 7735 33011 7741
rect 32953 7701 32965 7735
rect 32999 7732 33011 7735
rect 33042 7732 33048 7744
rect 32999 7704 33048 7732
rect 32999 7701 33011 7704
rect 32953 7695 33011 7701
rect 33042 7692 33048 7704
rect 33100 7692 33106 7744
rect 34146 7692 34152 7744
rect 34204 7692 34210 7744
rect 36538 7692 36544 7744
rect 36596 7732 36602 7744
rect 37645 7735 37703 7741
rect 37645 7732 37657 7735
rect 36596 7704 37657 7732
rect 36596 7692 36602 7704
rect 37645 7701 37657 7704
rect 37691 7701 37703 7735
rect 37645 7695 37703 7701
rect 37734 7692 37740 7744
rect 37792 7732 37798 7744
rect 39666 7732 39672 7744
rect 37792 7704 39672 7732
rect 37792 7692 37798 7704
rect 39666 7692 39672 7704
rect 39724 7692 39730 7744
rect 55677 7735 55735 7741
rect 55677 7701 55689 7735
rect 55723 7732 55735 7735
rect 56321 7735 56379 7741
rect 56321 7732 56333 7735
rect 55723 7704 56333 7732
rect 55723 7701 55735 7704
rect 55677 7695 55735 7701
rect 56321 7701 56333 7704
rect 56367 7701 56379 7735
rect 56321 7695 56379 7701
rect 1104 7642 58880 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 58880 7642
rect 1104 7568 58880 7590
rect 10594 7528 10600 7540
rect 10555 7500 10600 7528
rect 10594 7488 10600 7500
rect 10652 7488 10658 7540
rect 15010 7488 15016 7540
rect 15068 7528 15074 7540
rect 16758 7528 16764 7540
rect 15068 7500 16764 7528
rect 15068 7488 15074 7500
rect 16758 7488 16764 7500
rect 16816 7488 16822 7540
rect 17236 7500 17816 7528
rect 17236 7472 17264 7500
rect 1578 7420 1584 7472
rect 1636 7460 1642 7472
rect 10778 7460 10784 7472
rect 1636 7432 10784 7460
rect 1636 7420 1642 7432
rect 10778 7420 10784 7432
rect 10836 7420 10842 7472
rect 11977 7463 12035 7469
rect 11977 7460 11989 7463
rect 11440 7432 11989 7460
rect 11440 7404 11468 7432
rect 11977 7429 11989 7432
rect 12023 7429 12035 7463
rect 11977 7423 12035 7429
rect 15289 7463 15347 7469
rect 15289 7429 15301 7463
rect 15335 7460 15347 7463
rect 15470 7460 15476 7472
rect 15335 7432 15476 7460
rect 15335 7429 15347 7432
rect 15289 7423 15347 7429
rect 15470 7420 15476 7432
rect 15528 7420 15534 7472
rect 15654 7420 15660 7472
rect 15712 7460 15718 7472
rect 15841 7463 15899 7469
rect 15841 7460 15853 7463
rect 15712 7432 15853 7460
rect 15712 7420 15718 7432
rect 15841 7429 15853 7432
rect 15887 7429 15899 7463
rect 15841 7423 15899 7429
rect 9490 7392 9496 7404
rect 9451 7364 9496 7392
rect 9490 7352 9496 7364
rect 9548 7352 9554 7404
rect 9582 7352 9588 7404
rect 9640 7392 9646 7404
rect 10965 7395 11023 7401
rect 10965 7392 10977 7395
rect 9640 7364 10977 7392
rect 9640 7352 9646 7364
rect 10965 7361 10977 7364
rect 11011 7392 11023 7395
rect 11422 7392 11428 7404
rect 11011 7364 11428 7392
rect 11011 7361 11023 7364
rect 10965 7355 11023 7361
rect 11422 7352 11428 7364
rect 11480 7352 11486 7404
rect 11793 7395 11851 7401
rect 11793 7361 11805 7395
rect 11839 7392 11851 7395
rect 15746 7392 15752 7404
rect 11839 7364 12434 7392
rect 15707 7364 15752 7392
rect 11839 7361 11851 7364
rect 11793 7355 11851 7361
rect 12406 7336 12434 7364
rect 15746 7352 15752 7364
rect 15804 7352 15810 7404
rect 15856 7392 15884 7423
rect 16298 7420 16304 7472
rect 16356 7460 16362 7472
rect 16945 7463 17003 7469
rect 16945 7460 16957 7463
rect 16356 7432 16957 7460
rect 16356 7420 16362 7432
rect 16945 7429 16957 7432
rect 16991 7460 17003 7463
rect 17218 7460 17224 7472
rect 16991 7432 17224 7460
rect 16991 7429 17003 7432
rect 16945 7423 17003 7429
rect 17218 7420 17224 7432
rect 17276 7420 17282 7472
rect 17494 7420 17500 7472
rect 17552 7460 17558 7472
rect 17552 7432 17597 7460
rect 17552 7420 17558 7432
rect 16022 7392 16028 7404
rect 15856 7364 16028 7392
rect 16022 7352 16028 7364
rect 16080 7392 16086 7404
rect 17126 7392 17132 7404
rect 16080 7364 17132 7392
rect 16080 7352 16086 7364
rect 17126 7352 17132 7364
rect 17184 7392 17190 7404
rect 17359 7395 17417 7401
rect 17359 7392 17371 7395
rect 17184 7364 17371 7392
rect 17184 7352 17190 7364
rect 17359 7361 17371 7364
rect 17405 7361 17417 7395
rect 17788 7392 17816 7500
rect 18046 7488 18052 7540
rect 18104 7528 18110 7540
rect 19245 7531 19303 7537
rect 19245 7528 19257 7531
rect 18104 7500 19257 7528
rect 18104 7488 18110 7500
rect 19245 7497 19257 7500
rect 19291 7497 19303 7531
rect 19245 7491 19303 7497
rect 21450 7488 21456 7540
rect 21508 7528 21514 7540
rect 23474 7528 23480 7540
rect 21508 7500 23336 7528
rect 23435 7500 23480 7528
rect 21508 7488 21514 7500
rect 17862 7420 17868 7472
rect 17920 7460 17926 7472
rect 18509 7463 18567 7469
rect 18509 7460 18521 7463
rect 17920 7432 18521 7460
rect 17920 7420 17926 7432
rect 18509 7429 18521 7432
rect 18555 7429 18567 7463
rect 19058 7460 19064 7472
rect 19019 7432 19064 7460
rect 18509 7423 18567 7429
rect 19058 7420 19064 7432
rect 19116 7420 19122 7472
rect 19518 7420 19524 7472
rect 19576 7460 19582 7472
rect 19576 7432 21312 7460
rect 19576 7420 19582 7432
rect 18966 7392 18972 7404
rect 17788 7364 18972 7392
rect 17359 7355 17417 7361
rect 18966 7352 18972 7364
rect 19024 7352 19030 7404
rect 19426 7352 19432 7404
rect 19484 7392 19490 7404
rect 20073 7395 20131 7401
rect 20073 7392 20085 7395
rect 19484 7364 20085 7392
rect 19484 7352 19490 7364
rect 20073 7361 20085 7364
rect 20119 7361 20131 7395
rect 20073 7355 20131 7361
rect 20340 7395 20398 7401
rect 20340 7361 20352 7395
rect 20386 7392 20398 7395
rect 21174 7392 21180 7404
rect 20386 7364 21180 7392
rect 20386 7361 20398 7364
rect 20340 7355 20398 7361
rect 21174 7352 21180 7364
rect 21232 7352 21238 7404
rect 10686 7284 10692 7336
rect 10744 7324 10750 7336
rect 10781 7327 10839 7333
rect 10781 7324 10793 7327
rect 10744 7296 10793 7324
rect 10744 7284 10750 7296
rect 10781 7293 10793 7296
rect 10827 7293 10839 7327
rect 10781 7287 10839 7293
rect 10870 7284 10876 7336
rect 10928 7324 10934 7336
rect 10928 7296 10973 7324
rect 10928 7284 10934 7296
rect 11054 7284 11060 7336
rect 11112 7324 11118 7336
rect 11112 7296 11157 7324
rect 12406 7296 12440 7336
rect 11112 7284 11118 7296
rect 12434 7284 12440 7296
rect 12492 7324 12498 7336
rect 15381 7327 15439 7333
rect 12492 7296 12537 7324
rect 12492 7284 12498 7296
rect 15381 7293 15393 7327
rect 15427 7293 15439 7327
rect 16298 7324 16304 7336
rect 16259 7296 16304 7324
rect 15381 7287 15439 7293
rect 7374 7216 7380 7268
rect 7432 7256 7438 7268
rect 12713 7259 12771 7265
rect 12713 7256 12725 7259
rect 7432 7228 12725 7256
rect 7432 7216 7438 7228
rect 12713 7225 12725 7228
rect 12759 7225 12771 7259
rect 12713 7219 12771 7225
rect 12897 7259 12955 7265
rect 12897 7225 12909 7259
rect 12943 7256 12955 7259
rect 15194 7256 15200 7268
rect 12943 7228 15200 7256
rect 12943 7225 12955 7228
rect 12897 7219 12955 7225
rect 15194 7216 15200 7228
rect 15252 7216 15258 7268
rect 9398 7148 9404 7200
rect 9456 7188 9462 7200
rect 9677 7191 9735 7197
rect 9677 7188 9689 7191
rect 9456 7160 9689 7188
rect 9456 7148 9462 7160
rect 9677 7157 9689 7160
rect 9723 7157 9735 7191
rect 15396 7188 15424 7287
rect 16298 7284 16304 7296
rect 16356 7284 16362 7336
rect 17034 7284 17040 7336
rect 17092 7324 17098 7336
rect 17862 7324 17868 7336
rect 17092 7296 17137 7324
rect 17328 7296 17868 7324
rect 17092 7284 17098 7296
rect 17328 7268 17356 7296
rect 17862 7284 17868 7296
rect 17920 7324 17926 7336
rect 17957 7327 18015 7333
rect 17957 7324 17969 7327
rect 17920 7296 17969 7324
rect 17920 7284 17926 7296
rect 17957 7293 17969 7296
rect 18003 7293 18015 7327
rect 17957 7287 18015 7293
rect 19058 7284 19064 7336
rect 19116 7324 19122 7336
rect 19886 7324 19892 7336
rect 19116 7296 19892 7324
rect 19116 7284 19122 7296
rect 19886 7284 19892 7296
rect 19944 7284 19950 7336
rect 21284 7324 21312 7432
rect 23308 7401 23336 7500
rect 23474 7488 23480 7500
rect 23532 7488 23538 7540
rect 27798 7528 27804 7540
rect 23584 7500 27804 7528
rect 23293 7395 23351 7401
rect 23293 7361 23305 7395
rect 23339 7361 23351 7395
rect 23293 7355 23351 7361
rect 23584 7324 23612 7500
rect 27798 7488 27804 7500
rect 27856 7528 27862 7540
rect 27893 7531 27951 7537
rect 27893 7528 27905 7531
rect 27856 7500 27905 7528
rect 27856 7488 27862 7500
rect 27893 7497 27905 7500
rect 27939 7528 27951 7531
rect 29270 7528 29276 7540
rect 27939 7500 29276 7528
rect 27939 7497 27951 7500
rect 27893 7491 27951 7497
rect 29270 7488 29276 7500
rect 29328 7488 29334 7540
rect 29914 7528 29920 7540
rect 29875 7500 29920 7528
rect 29914 7488 29920 7500
rect 29972 7528 29978 7540
rect 30190 7528 30196 7540
rect 29972 7500 30196 7528
rect 29972 7488 29978 7500
rect 30190 7488 30196 7500
rect 30248 7488 30254 7540
rect 30466 7488 30472 7540
rect 30524 7528 30530 7540
rect 31570 7528 31576 7540
rect 30524 7500 31576 7528
rect 30524 7488 30530 7500
rect 31570 7488 31576 7500
rect 31628 7528 31634 7540
rect 35434 7528 35440 7540
rect 31628 7500 35296 7528
rect 35395 7500 35440 7528
rect 31628 7488 31634 7500
rect 27338 7460 27344 7472
rect 23676 7432 27344 7460
rect 23676 7401 23704 7432
rect 27338 7420 27344 7432
rect 27396 7420 27402 7472
rect 27614 7460 27620 7472
rect 27448 7432 27620 7460
rect 27448 7401 27476 7432
rect 27614 7420 27620 7432
rect 27672 7420 27678 7472
rect 28166 7420 28172 7472
rect 28224 7460 28230 7472
rect 30208 7460 30236 7488
rect 35158 7460 35164 7472
rect 28224 7432 28994 7460
rect 30208 7432 35164 7460
rect 28224 7420 28230 7432
rect 23661 7395 23719 7401
rect 23661 7361 23673 7395
rect 23707 7361 23719 7395
rect 23661 7355 23719 7361
rect 24305 7395 24363 7401
rect 24305 7361 24317 7395
rect 24351 7392 24363 7395
rect 27433 7395 27491 7401
rect 24351 7364 26004 7392
rect 24351 7361 24363 7364
rect 24305 7355 24363 7361
rect 21284 7296 23612 7324
rect 17310 7216 17316 7268
rect 17368 7216 17374 7268
rect 18046 7216 18052 7268
rect 18104 7256 18110 7268
rect 18491 7259 18549 7265
rect 18491 7256 18503 7259
rect 18104 7228 18503 7256
rect 18104 7216 18110 7228
rect 18491 7225 18503 7228
rect 18537 7225 18549 7259
rect 18491 7219 18549 7225
rect 19150 7216 19156 7268
rect 19208 7256 19214 7268
rect 19978 7256 19984 7268
rect 19208 7228 19984 7256
rect 19208 7216 19214 7228
rect 19978 7216 19984 7228
rect 20036 7216 20042 7268
rect 21082 7216 21088 7268
rect 21140 7256 21146 7268
rect 25501 7259 25559 7265
rect 25501 7256 25513 7259
rect 21140 7228 25513 7256
rect 21140 7216 21146 7228
rect 25501 7225 25513 7228
rect 25547 7225 25559 7259
rect 25501 7219 25559 7225
rect 21266 7188 21272 7200
rect 15396 7160 21272 7188
rect 9677 7151 9735 7157
rect 21266 7148 21272 7160
rect 21324 7148 21330 7200
rect 21450 7188 21456 7200
rect 21411 7160 21456 7188
rect 21450 7148 21456 7160
rect 21508 7148 21514 7200
rect 21542 7148 21548 7200
rect 21600 7188 21606 7200
rect 23845 7191 23903 7197
rect 23845 7188 23857 7191
rect 21600 7160 23857 7188
rect 21600 7148 21606 7160
rect 23845 7157 23857 7160
rect 23891 7188 23903 7191
rect 25682 7188 25688 7200
rect 23891 7160 25688 7188
rect 23891 7157 23903 7160
rect 23845 7151 23903 7157
rect 25682 7148 25688 7160
rect 25740 7148 25746 7200
rect 25976 7188 26004 7364
rect 27433 7361 27445 7395
rect 27479 7361 27491 7395
rect 27433 7355 27491 7361
rect 27522 7352 27528 7404
rect 27580 7392 27586 7404
rect 27709 7395 27767 7401
rect 27580 7364 27625 7392
rect 27580 7352 27586 7364
rect 27709 7361 27721 7395
rect 27755 7361 27767 7395
rect 28626 7392 28632 7404
rect 28587 7364 28632 7392
rect 27709 7355 27767 7361
rect 27724 7256 27752 7355
rect 28626 7352 28632 7364
rect 28684 7352 28690 7404
rect 28966 7392 28994 7432
rect 30837 7395 30895 7401
rect 30837 7392 30849 7395
rect 28966 7364 30849 7392
rect 30837 7361 30849 7364
rect 30883 7361 30895 7395
rect 32582 7392 32588 7404
rect 32543 7364 32588 7392
rect 30837 7355 30895 7361
rect 32582 7352 32588 7364
rect 32640 7352 32646 7404
rect 32766 7392 32772 7404
rect 32727 7364 32772 7392
rect 32766 7352 32772 7364
rect 32824 7352 32830 7404
rect 32861 7395 32919 7401
rect 32861 7361 32873 7395
rect 32907 7392 32919 7395
rect 33226 7392 33232 7404
rect 32907 7364 33232 7392
rect 32907 7361 32919 7364
rect 32861 7355 32919 7361
rect 33226 7352 33232 7364
rect 33284 7352 33290 7404
rect 34072 7401 34100 7432
rect 35158 7420 35164 7432
rect 35216 7420 35222 7472
rect 35268 7460 35296 7500
rect 35434 7488 35440 7500
rect 35492 7488 35498 7540
rect 36173 7531 36231 7537
rect 36173 7497 36185 7531
rect 36219 7528 36231 7531
rect 36722 7528 36728 7540
rect 36219 7500 36728 7528
rect 36219 7497 36231 7500
rect 36173 7491 36231 7497
rect 36722 7488 36728 7500
rect 36780 7488 36786 7540
rect 38562 7488 38568 7540
rect 38620 7528 38626 7540
rect 44450 7528 44456 7540
rect 38620 7500 44456 7528
rect 38620 7488 38626 7500
rect 44450 7488 44456 7500
rect 44508 7488 44514 7540
rect 52454 7488 52460 7540
rect 52512 7528 52518 7540
rect 56502 7528 56508 7540
rect 52512 7500 56508 7528
rect 52512 7488 52518 7500
rect 56502 7488 56508 7500
rect 56560 7488 56566 7540
rect 35342 7460 35348 7472
rect 35268 7432 35348 7460
rect 35342 7420 35348 7432
rect 35400 7420 35406 7472
rect 35986 7420 35992 7472
rect 36044 7460 36050 7472
rect 55766 7460 55772 7472
rect 36044 7432 55772 7460
rect 36044 7420 36050 7432
rect 55766 7420 55772 7432
rect 55824 7420 55830 7472
rect 55861 7463 55919 7469
rect 55861 7429 55873 7463
rect 55907 7460 55919 7463
rect 58161 7463 58219 7469
rect 58161 7460 58173 7463
rect 55907 7432 58173 7460
rect 55907 7429 55919 7432
rect 55861 7423 55919 7429
rect 58161 7429 58173 7432
rect 58207 7429 58219 7463
rect 58161 7423 58219 7429
rect 34330 7401 34336 7404
rect 34057 7395 34115 7401
rect 34057 7361 34069 7395
rect 34103 7361 34115 7395
rect 34057 7355 34115 7361
rect 34324 7355 34336 7401
rect 34388 7392 34394 7404
rect 34388 7364 34424 7392
rect 34330 7352 34336 7355
rect 34388 7352 34394 7364
rect 34698 7352 34704 7404
rect 34756 7392 34762 7404
rect 35710 7392 35716 7404
rect 34756 7364 35716 7392
rect 34756 7352 34762 7364
rect 35710 7352 35716 7364
rect 35768 7352 35774 7404
rect 36538 7392 36544 7404
rect 36499 7364 36544 7392
rect 36538 7352 36544 7364
rect 36596 7352 36602 7404
rect 36633 7395 36691 7401
rect 36633 7361 36645 7395
rect 36679 7392 36691 7395
rect 36906 7392 36912 7404
rect 36679 7364 36912 7392
rect 36679 7361 36691 7364
rect 36633 7355 36691 7361
rect 36906 7352 36912 7364
rect 36964 7352 36970 7404
rect 43898 7352 43904 7404
rect 43956 7392 43962 7404
rect 44361 7395 44419 7401
rect 44361 7392 44373 7395
rect 43956 7364 44373 7392
rect 43956 7352 43962 7364
rect 44361 7361 44373 7364
rect 44407 7361 44419 7395
rect 44361 7355 44419 7361
rect 44453 7395 44511 7401
rect 44453 7361 44465 7395
rect 44499 7392 44511 7395
rect 44542 7392 44548 7404
rect 44499 7364 44548 7392
rect 44499 7361 44511 7364
rect 44453 7355 44511 7361
rect 29086 7324 29092 7336
rect 28184 7296 29092 7324
rect 28184 7256 28212 7296
rect 29086 7284 29092 7296
rect 29144 7324 29150 7336
rect 30006 7324 30012 7336
rect 29144 7296 30012 7324
rect 29144 7284 29150 7296
rect 30006 7284 30012 7296
rect 30064 7284 30070 7336
rect 31021 7327 31079 7333
rect 31021 7324 31033 7327
rect 30116 7296 31033 7324
rect 27724 7228 28212 7256
rect 28258 7216 28264 7268
rect 28316 7256 28322 7268
rect 30116 7256 30144 7296
rect 31021 7293 31033 7296
rect 31067 7293 31079 7327
rect 33134 7324 33140 7336
rect 31021 7287 31079 7293
rect 31726 7296 33140 7324
rect 28316 7228 30144 7256
rect 28316 7216 28322 7228
rect 30374 7216 30380 7268
rect 30432 7256 30438 7268
rect 31726 7256 31754 7296
rect 33134 7284 33140 7296
rect 33192 7284 33198 7336
rect 35342 7284 35348 7336
rect 35400 7324 35406 7336
rect 36725 7327 36783 7333
rect 36725 7324 36737 7327
rect 35400 7296 36737 7324
rect 35400 7284 35406 7296
rect 36725 7293 36737 7296
rect 36771 7324 36783 7327
rect 38562 7324 38568 7336
rect 36771 7296 38568 7324
rect 36771 7293 36783 7296
rect 36725 7287 36783 7293
rect 38562 7284 38568 7296
rect 38620 7284 38626 7336
rect 40126 7284 40132 7336
rect 40184 7324 40190 7336
rect 43162 7324 43168 7336
rect 40184 7296 43168 7324
rect 40184 7284 40190 7296
rect 43162 7284 43168 7296
rect 43220 7284 43226 7336
rect 30432 7228 31754 7256
rect 30432 7216 30438 7228
rect 32214 7216 32220 7268
rect 32272 7256 32278 7268
rect 33870 7256 33876 7268
rect 32272 7228 33876 7256
rect 32272 7216 32278 7228
rect 33870 7216 33876 7228
rect 33928 7216 33934 7268
rect 37274 7256 37280 7268
rect 35360 7228 37280 7256
rect 30558 7188 30564 7200
rect 25976 7160 30564 7188
rect 30558 7148 30564 7160
rect 30616 7148 30622 7200
rect 32401 7191 32459 7197
rect 32401 7157 32413 7191
rect 32447 7188 32459 7191
rect 35360 7188 35388 7228
rect 37274 7216 37280 7228
rect 37332 7216 37338 7268
rect 32447 7160 35388 7188
rect 35897 7191 35955 7197
rect 32447 7157 32459 7160
rect 32401 7151 32459 7157
rect 35897 7157 35909 7191
rect 35943 7188 35955 7191
rect 35986 7188 35992 7200
rect 35943 7160 35992 7188
rect 35943 7157 35955 7160
rect 35897 7151 35955 7157
rect 35986 7148 35992 7160
rect 36044 7188 36050 7200
rect 36906 7188 36912 7200
rect 36044 7160 36912 7188
rect 36044 7148 36050 7160
rect 36906 7148 36912 7160
rect 36964 7148 36970 7200
rect 44376 7188 44404 7355
rect 44542 7352 44548 7364
rect 44600 7352 44606 7404
rect 45005 7395 45063 7401
rect 45005 7361 45017 7395
rect 45051 7392 45063 7395
rect 45094 7392 45100 7404
rect 45051 7364 45100 7392
rect 45051 7361 45063 7364
rect 45005 7355 45063 7361
rect 45094 7352 45100 7364
rect 45152 7352 45158 7404
rect 45272 7395 45330 7401
rect 45272 7361 45284 7395
rect 45318 7392 45330 7395
rect 45830 7392 45836 7404
rect 45318 7364 45836 7392
rect 45318 7361 45330 7364
rect 45272 7355 45330 7361
rect 45830 7352 45836 7364
rect 45888 7352 45894 7404
rect 55677 7395 55735 7401
rect 55677 7361 55689 7395
rect 55723 7361 55735 7395
rect 55950 7392 55956 7404
rect 55911 7364 55956 7392
rect 55677 7355 55735 7361
rect 55692 7324 55720 7355
rect 55950 7352 55956 7364
rect 56008 7352 56014 7404
rect 56502 7392 56508 7404
rect 56463 7364 56508 7392
rect 56502 7352 56508 7364
rect 56560 7352 56566 7404
rect 56962 7352 56968 7404
rect 57020 7392 57026 7404
rect 58069 7395 58127 7401
rect 58069 7392 58081 7395
rect 57020 7364 58081 7392
rect 57020 7352 57026 7364
rect 58069 7361 58081 7364
rect 58115 7361 58127 7395
rect 58250 7392 58256 7404
rect 58211 7364 58256 7392
rect 58069 7355 58127 7361
rect 58250 7352 58256 7364
rect 58308 7352 58314 7404
rect 56134 7324 56140 7336
rect 55692 7296 56140 7324
rect 56134 7284 56140 7296
rect 56192 7324 56198 7336
rect 56781 7327 56839 7333
rect 56781 7324 56793 7327
rect 56192 7296 56793 7324
rect 56192 7284 56198 7296
rect 56781 7293 56793 7296
rect 56827 7293 56839 7327
rect 56781 7287 56839 7293
rect 45922 7188 45928 7200
rect 44376 7160 45928 7188
rect 45922 7148 45928 7160
rect 45980 7148 45986 7200
rect 46382 7188 46388 7200
rect 46343 7160 46388 7188
rect 46382 7148 46388 7160
rect 46440 7148 46446 7200
rect 55677 7191 55735 7197
rect 55677 7157 55689 7191
rect 55723 7188 55735 7191
rect 56962 7188 56968 7200
rect 55723 7160 56968 7188
rect 55723 7157 55735 7160
rect 55677 7151 55735 7157
rect 56962 7148 56968 7160
rect 57020 7148 57026 7200
rect 1104 7098 58880 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 58880 7098
rect 1104 7024 58880 7046
rect 10870 6944 10876 6996
rect 10928 6984 10934 6996
rect 20530 6984 20536 6996
rect 10928 6956 20536 6984
rect 10928 6944 10934 6956
rect 20530 6944 20536 6956
rect 20588 6944 20594 6996
rect 21174 6984 21180 6996
rect 21135 6956 21180 6984
rect 21174 6944 21180 6956
rect 21232 6944 21238 6996
rect 21266 6944 21272 6996
rect 21324 6984 21330 6996
rect 27154 6984 27160 6996
rect 21324 6956 27160 6984
rect 21324 6944 21330 6956
rect 27154 6944 27160 6956
rect 27212 6944 27218 6996
rect 27706 6944 27712 6996
rect 27764 6944 27770 6996
rect 27890 6944 27896 6996
rect 27948 6984 27954 6996
rect 31846 6984 31852 6996
rect 27948 6956 31852 6984
rect 27948 6944 27954 6956
rect 31846 6944 31852 6956
rect 31904 6984 31910 6996
rect 34330 6984 34336 6996
rect 31904 6956 33364 6984
rect 34291 6956 34336 6984
rect 31904 6944 31910 6956
rect 18138 6876 18144 6928
rect 18196 6916 18202 6928
rect 20714 6916 20720 6928
rect 18196 6888 20720 6916
rect 18196 6876 18202 6888
rect 20714 6876 20720 6888
rect 20772 6876 20778 6928
rect 23842 6916 23848 6928
rect 23803 6888 23848 6916
rect 23842 6876 23848 6888
rect 23900 6876 23906 6928
rect 27724 6916 27752 6944
rect 30834 6916 30840 6928
rect 27172 6888 27752 6916
rect 30795 6888 30840 6916
rect 8754 6808 8760 6860
rect 8812 6848 8818 6860
rect 10778 6848 10784 6860
rect 8812 6820 9536 6848
rect 10739 6820 10784 6848
rect 8812 6808 8818 6820
rect 1581 6783 1639 6789
rect 1581 6749 1593 6783
rect 1627 6780 1639 6783
rect 9122 6780 9128 6792
rect 1627 6752 9128 6780
rect 1627 6749 1639 6752
rect 1581 6743 1639 6749
rect 9122 6740 9128 6752
rect 9180 6740 9186 6792
rect 9508 6780 9536 6820
rect 10778 6808 10784 6820
rect 10836 6808 10842 6860
rect 10870 6808 10876 6860
rect 10928 6848 10934 6860
rect 18598 6848 18604 6860
rect 10928 6820 18604 6848
rect 10928 6808 10934 6820
rect 18598 6808 18604 6820
rect 18656 6808 18662 6860
rect 18693 6851 18751 6857
rect 18693 6817 18705 6851
rect 18739 6817 18751 6851
rect 18693 6811 18751 6817
rect 9582 6780 9588 6792
rect 9495 6752 9588 6780
rect 9582 6740 9588 6752
rect 9640 6740 9646 6792
rect 10686 6740 10692 6792
rect 10744 6780 10750 6792
rect 10965 6783 11023 6789
rect 10965 6780 10977 6783
rect 10744 6752 10977 6780
rect 10744 6740 10750 6752
rect 10965 6749 10977 6752
rect 11011 6749 11023 6783
rect 10965 6743 11023 6749
rect 11057 6783 11115 6789
rect 11057 6749 11069 6783
rect 11103 6749 11115 6783
rect 11057 6743 11115 6749
rect 11149 6783 11207 6789
rect 11149 6749 11161 6783
rect 11195 6749 11207 6783
rect 11149 6743 11207 6749
rect 1854 6712 1860 6724
rect 1815 6684 1860 6712
rect 1854 6672 1860 6684
rect 1912 6672 1918 6724
rect 9490 6604 9496 6656
rect 9548 6644 9554 6656
rect 9674 6644 9680 6656
rect 9548 6616 9680 6644
rect 9548 6604 9554 6616
rect 9674 6604 9680 6616
rect 9732 6644 9738 6656
rect 9769 6647 9827 6653
rect 9769 6644 9781 6647
rect 9732 6616 9781 6644
rect 9732 6604 9738 6616
rect 9769 6613 9781 6616
rect 9815 6613 9827 6647
rect 11072 6644 11100 6743
rect 11164 6712 11192 6743
rect 11238 6740 11244 6792
rect 11296 6780 11302 6792
rect 16577 6783 16635 6789
rect 11296 6752 11341 6780
rect 11296 6740 11302 6752
rect 16577 6749 16589 6783
rect 16623 6780 16635 6783
rect 17402 6780 17408 6792
rect 16623 6752 17408 6780
rect 16623 6749 16635 6752
rect 16577 6743 16635 6749
rect 17402 6740 17408 6752
rect 17460 6740 17466 6792
rect 17770 6740 17776 6792
rect 17828 6780 17834 6792
rect 17954 6780 17960 6792
rect 17828 6752 17960 6780
rect 17828 6740 17834 6752
rect 17954 6740 17960 6752
rect 18012 6740 18018 6792
rect 18506 6740 18512 6792
rect 18564 6780 18570 6792
rect 18708 6780 18736 6811
rect 18966 6808 18972 6860
rect 19024 6848 19030 6860
rect 19797 6851 19855 6857
rect 19797 6848 19809 6851
rect 19024 6820 19809 6848
rect 19024 6808 19030 6820
rect 19797 6817 19809 6820
rect 19843 6817 19855 6851
rect 19797 6811 19855 6817
rect 21174 6808 21180 6860
rect 21232 6848 21238 6860
rect 21726 6848 21732 6860
rect 21232 6820 21732 6848
rect 21232 6808 21238 6820
rect 21726 6808 21732 6820
rect 21784 6808 21790 6860
rect 26513 6851 26571 6857
rect 26513 6817 26525 6851
rect 26559 6848 26571 6851
rect 26786 6848 26792 6860
rect 26559 6820 26792 6848
rect 26559 6817 26571 6820
rect 26513 6811 26571 6817
rect 26786 6808 26792 6820
rect 26844 6848 26850 6860
rect 27062 6848 27068 6860
rect 26844 6820 27068 6848
rect 26844 6808 26850 6820
rect 27062 6808 27068 6820
rect 27120 6808 27126 6860
rect 18564 6752 18736 6780
rect 18564 6740 18570 6752
rect 11422 6712 11428 6724
rect 11164 6684 11428 6712
rect 11422 6672 11428 6684
rect 11480 6672 11486 6724
rect 17313 6715 17371 6721
rect 17313 6681 17325 6715
rect 17359 6712 17371 6715
rect 17494 6712 17500 6724
rect 17359 6684 17500 6712
rect 17359 6681 17371 6684
rect 17313 6675 17371 6681
rect 17494 6672 17500 6684
rect 17552 6672 17558 6724
rect 17865 6715 17923 6721
rect 17865 6681 17877 6715
rect 17911 6712 17923 6715
rect 18708 6712 18736 6752
rect 19334 6740 19340 6792
rect 19392 6780 19398 6792
rect 19521 6783 19579 6789
rect 19521 6780 19533 6783
rect 19392 6752 19533 6780
rect 19392 6740 19398 6752
rect 19521 6749 19533 6752
rect 19567 6749 19579 6783
rect 19521 6743 19579 6749
rect 19610 6740 19616 6792
rect 19668 6780 19674 6792
rect 22465 6783 22523 6789
rect 22465 6780 22477 6783
rect 19668 6752 22477 6780
rect 19668 6740 19674 6752
rect 22465 6749 22477 6752
rect 22511 6780 22523 6783
rect 24670 6780 24676 6792
rect 22511 6752 24676 6780
rect 22511 6749 22523 6752
rect 22465 6743 22523 6749
rect 24670 6740 24676 6752
rect 24728 6740 24734 6792
rect 27172 6789 27200 6888
rect 30834 6876 30840 6888
rect 30892 6876 30898 6928
rect 31570 6876 31576 6928
rect 31628 6916 31634 6928
rect 33336 6916 33364 6956
rect 34330 6944 34336 6956
rect 34388 6944 34394 6996
rect 45189 6987 45247 6993
rect 34440 6956 36492 6984
rect 34440 6916 34468 6956
rect 31628 6888 31984 6916
rect 33336 6888 34468 6916
rect 34885 6919 34943 6925
rect 31628 6876 31634 6888
rect 27249 6851 27307 6857
rect 27249 6817 27261 6851
rect 27295 6848 27307 6851
rect 27706 6848 27712 6860
rect 27295 6820 27712 6848
rect 27295 6817 27307 6820
rect 27249 6811 27307 6817
rect 27706 6808 27712 6820
rect 27764 6808 27770 6860
rect 28074 6808 28080 6860
rect 28132 6848 28138 6860
rect 28534 6848 28540 6860
rect 28132 6820 28540 6848
rect 28132 6808 28138 6820
rect 28534 6808 28540 6820
rect 28592 6808 28598 6860
rect 29822 6808 29828 6860
rect 29880 6848 29886 6860
rect 30193 6851 30251 6857
rect 30193 6848 30205 6851
rect 29880 6820 30205 6848
rect 29880 6808 29886 6820
rect 30193 6817 30205 6820
rect 30239 6848 30251 6851
rect 31018 6848 31024 6860
rect 30239 6820 31024 6848
rect 30239 6817 30251 6820
rect 30193 6811 30251 6817
rect 31018 6808 31024 6820
rect 31076 6808 31082 6860
rect 31662 6808 31668 6860
rect 31720 6848 31726 6860
rect 31956 6857 31984 6888
rect 34885 6885 34897 6919
rect 34931 6885 34943 6919
rect 34885 6879 34943 6885
rect 31849 6851 31907 6857
rect 31849 6848 31861 6851
rect 31720 6820 31861 6848
rect 31720 6808 31726 6820
rect 31849 6817 31861 6820
rect 31895 6817 31907 6851
rect 31849 6811 31907 6817
rect 31941 6851 31999 6857
rect 31941 6817 31953 6851
rect 31987 6817 31999 6851
rect 31941 6811 31999 6817
rect 32585 6851 32643 6857
rect 32585 6817 32597 6851
rect 32631 6848 32643 6851
rect 33134 6848 33140 6860
rect 32631 6820 33140 6848
rect 32631 6817 32643 6820
rect 32585 6811 32643 6817
rect 33134 6808 33140 6820
rect 33192 6848 33198 6860
rect 33965 6851 34023 6857
rect 33965 6848 33977 6851
rect 33192 6820 33977 6848
rect 33192 6808 33198 6820
rect 33965 6817 33977 6820
rect 34011 6817 34023 6851
rect 34422 6848 34428 6860
rect 33965 6811 34023 6817
rect 34072 6820 34428 6848
rect 27157 6783 27215 6789
rect 27157 6749 27169 6783
rect 27203 6749 27215 6783
rect 27157 6743 27215 6749
rect 27491 6783 27549 6789
rect 27491 6749 27503 6783
rect 27537 6749 27549 6783
rect 27491 6743 27549 6749
rect 27617 6783 27675 6789
rect 27617 6749 27629 6783
rect 27663 6780 27675 6783
rect 27982 6780 27988 6792
rect 27663 6752 27988 6780
rect 27663 6749 27675 6752
rect 27617 6743 27675 6749
rect 21174 6712 21180 6724
rect 17911 6684 18552 6712
rect 18708 6684 21180 6712
rect 17911 6681 17923 6684
rect 17865 6675 17923 6681
rect 18524 6656 18552 6684
rect 21174 6672 21180 6684
rect 21232 6672 21238 6724
rect 21545 6715 21603 6721
rect 21545 6681 21557 6715
rect 21591 6712 21603 6715
rect 21591 6684 22094 6712
rect 21591 6681 21603 6684
rect 21545 6675 21603 6681
rect 16206 6644 16212 6656
rect 11072 6616 16212 6644
rect 9769 6607 9827 6613
rect 16206 6604 16212 6616
rect 16264 6604 16270 6656
rect 18138 6644 18144 6656
rect 18099 6616 18144 6644
rect 18138 6604 18144 6616
rect 18196 6604 18202 6656
rect 18506 6644 18512 6656
rect 18467 6616 18512 6644
rect 18506 6604 18512 6616
rect 18564 6604 18570 6656
rect 18598 6604 18604 6656
rect 18656 6644 18662 6656
rect 18656 6616 18701 6644
rect 18656 6604 18662 6616
rect 20714 6604 20720 6656
rect 20772 6644 20778 6656
rect 21450 6644 21456 6656
rect 20772 6616 21456 6644
rect 20772 6604 20778 6616
rect 21450 6604 21456 6616
rect 21508 6644 21514 6656
rect 21637 6647 21695 6653
rect 21637 6644 21649 6647
rect 21508 6616 21649 6644
rect 21508 6604 21514 6616
rect 21637 6613 21649 6616
rect 21683 6613 21695 6647
rect 22066 6644 22094 6684
rect 22278 6672 22284 6724
rect 22336 6712 22342 6724
rect 22732 6715 22790 6721
rect 22732 6712 22744 6715
rect 22336 6684 22744 6712
rect 22336 6672 22342 6684
rect 22732 6681 22744 6684
rect 22778 6681 22790 6715
rect 22732 6675 22790 6681
rect 23290 6672 23296 6724
rect 23348 6712 23354 6724
rect 24762 6712 24768 6724
rect 23348 6684 24768 6712
rect 23348 6672 23354 6684
rect 24762 6672 24768 6684
rect 24820 6672 24826 6724
rect 24940 6715 24998 6721
rect 24940 6681 24952 6715
rect 24986 6712 24998 6715
rect 25590 6712 25596 6724
rect 24986 6684 25596 6712
rect 24986 6681 24998 6684
rect 24940 6675 24998 6681
rect 25590 6672 25596 6684
rect 25648 6672 25654 6724
rect 26418 6672 26424 6724
rect 26476 6712 26482 6724
rect 27494 6712 27522 6743
rect 27982 6740 27988 6752
rect 28040 6740 28046 6792
rect 28166 6780 28172 6792
rect 28127 6752 28172 6780
rect 28166 6740 28172 6752
rect 28224 6740 28230 6792
rect 30009 6783 30067 6789
rect 30009 6749 30021 6783
rect 30055 6749 30067 6783
rect 30009 6743 30067 6749
rect 30101 6783 30159 6789
rect 30101 6749 30113 6783
rect 30147 6780 30159 6783
rect 31478 6780 31484 6792
rect 30147 6752 31484 6780
rect 30147 6749 30159 6752
rect 30101 6743 30159 6749
rect 27798 6712 27804 6724
rect 26476 6684 27804 6712
rect 26476 6672 26482 6684
rect 27798 6672 27804 6684
rect 27856 6672 27862 6724
rect 22922 6644 22928 6656
rect 22066 6616 22928 6644
rect 21637 6607 21695 6613
rect 22922 6604 22928 6616
rect 22980 6604 22986 6656
rect 25130 6604 25136 6656
rect 25188 6644 25194 6656
rect 26053 6647 26111 6653
rect 26053 6644 26065 6647
rect 25188 6616 26065 6644
rect 25188 6604 25194 6616
rect 26053 6613 26065 6616
rect 26099 6613 26111 6647
rect 26053 6607 26111 6613
rect 26510 6604 26516 6656
rect 26568 6644 26574 6656
rect 30024 6644 30052 6743
rect 31478 6740 31484 6752
rect 31536 6740 31542 6792
rect 31570 6740 31576 6792
rect 31628 6780 31634 6792
rect 31757 6783 31815 6789
rect 31757 6780 31769 6783
rect 31628 6752 31769 6780
rect 31628 6740 31634 6752
rect 31757 6749 31769 6752
rect 31803 6780 31815 6783
rect 32674 6780 32680 6792
rect 31803 6752 32680 6780
rect 31803 6749 31815 6752
rect 31757 6743 31815 6749
rect 32674 6740 32680 6752
rect 32732 6740 32738 6792
rect 32769 6783 32827 6789
rect 32769 6749 32781 6783
rect 32815 6780 32827 6783
rect 32815 6752 32904 6780
rect 32815 6749 32827 6752
rect 32769 6743 32827 6749
rect 30374 6672 30380 6724
rect 30432 6712 30438 6724
rect 30469 6715 30527 6721
rect 30469 6712 30481 6715
rect 30432 6684 30481 6712
rect 30432 6672 30438 6684
rect 30469 6681 30481 6684
rect 30515 6681 30527 6715
rect 30469 6675 30527 6681
rect 30282 6644 30288 6656
rect 26568 6616 30288 6644
rect 26568 6604 26574 6616
rect 30282 6604 30288 6616
rect 30340 6604 30346 6656
rect 31389 6647 31447 6653
rect 31389 6613 31401 6647
rect 31435 6644 31447 6647
rect 32876 6644 32904 6752
rect 32950 6740 32956 6792
rect 33008 6780 33014 6792
rect 33008 6752 33053 6780
rect 33008 6740 33014 6752
rect 33686 6740 33692 6792
rect 33744 6780 33750 6792
rect 34072 6780 34100 6820
rect 34422 6808 34428 6820
rect 34480 6808 34486 6860
rect 33744 6752 34100 6780
rect 34149 6783 34207 6789
rect 33744 6740 33750 6752
rect 34149 6749 34161 6783
rect 34195 6780 34207 6783
rect 34900 6780 34928 6879
rect 35342 6808 35348 6860
rect 35400 6848 35406 6860
rect 35437 6851 35495 6857
rect 35437 6848 35449 6851
rect 35400 6820 35449 6848
rect 35400 6808 35406 6820
rect 35437 6817 35449 6820
rect 35483 6817 35495 6851
rect 35437 6811 35495 6817
rect 36464 6789 36492 6956
rect 45189 6953 45201 6987
rect 45235 6984 45247 6987
rect 45278 6984 45284 6996
rect 45235 6956 45284 6984
rect 45235 6953 45247 6956
rect 45189 6947 45247 6953
rect 45278 6944 45284 6956
rect 45336 6944 45342 6996
rect 45830 6984 45836 6996
rect 45791 6956 45836 6984
rect 45830 6944 45836 6956
rect 45888 6944 45894 6996
rect 45922 6944 45928 6996
rect 45980 6984 45986 6996
rect 58342 6984 58348 6996
rect 45980 6956 58348 6984
rect 45980 6944 45986 6956
rect 58342 6944 58348 6956
rect 58400 6944 58406 6996
rect 36541 6851 36599 6857
rect 36541 6817 36553 6851
rect 36587 6848 36599 6851
rect 37182 6848 37188 6860
rect 36587 6820 37188 6848
rect 36587 6817 36599 6820
rect 36541 6811 36599 6817
rect 37182 6808 37188 6820
rect 37240 6808 37246 6860
rect 38654 6808 38660 6860
rect 38712 6848 38718 6860
rect 46293 6851 46351 6857
rect 46293 6848 46305 6851
rect 38712 6820 46305 6848
rect 38712 6808 38718 6820
rect 46293 6817 46305 6820
rect 46339 6848 46351 6851
rect 46382 6848 46388 6860
rect 46339 6820 46388 6848
rect 46339 6817 46351 6820
rect 46293 6811 46351 6817
rect 46382 6808 46388 6820
rect 46440 6808 46446 6860
rect 46477 6851 46535 6857
rect 46477 6817 46489 6851
rect 46523 6848 46535 6851
rect 46658 6848 46664 6860
rect 46523 6820 46664 6848
rect 46523 6817 46535 6820
rect 46477 6811 46535 6817
rect 46658 6808 46664 6820
rect 46716 6808 46722 6860
rect 48774 6808 48780 6860
rect 48832 6848 48838 6860
rect 48832 6820 56916 6848
rect 48832 6808 48838 6820
rect 56888 6792 56916 6820
rect 34195 6752 34928 6780
rect 36449 6783 36507 6789
rect 34195 6749 34207 6752
rect 34149 6743 34207 6749
rect 36449 6749 36461 6783
rect 36495 6749 36507 6783
rect 36449 6743 36507 6749
rect 36633 6783 36691 6789
rect 36633 6749 36645 6783
rect 36679 6780 36691 6783
rect 36722 6780 36728 6792
rect 36679 6752 36728 6780
rect 36679 6749 36691 6752
rect 36633 6743 36691 6749
rect 36722 6740 36728 6752
rect 36780 6740 36786 6792
rect 44542 6740 44548 6792
rect 44600 6780 44606 6792
rect 45189 6783 45247 6789
rect 45189 6780 45201 6783
rect 44600 6752 45201 6780
rect 44600 6740 44606 6752
rect 45189 6749 45201 6752
rect 45235 6749 45247 6783
rect 45189 6743 45247 6749
rect 45373 6783 45431 6789
rect 45373 6749 45385 6783
rect 45419 6780 45431 6783
rect 45462 6780 45468 6792
rect 45419 6752 45468 6780
rect 45419 6749 45431 6752
rect 45373 6743 45431 6749
rect 45462 6740 45468 6752
rect 45520 6740 45526 6792
rect 48222 6780 48228 6792
rect 45572 6752 48228 6780
rect 33226 6672 33232 6724
rect 33284 6712 33290 6724
rect 35345 6715 35403 6721
rect 35345 6712 35357 6715
rect 33284 6684 35357 6712
rect 33284 6672 33290 6684
rect 35345 6681 35357 6684
rect 35391 6712 35403 6715
rect 35618 6712 35624 6724
rect 35391 6684 35624 6712
rect 35391 6681 35403 6684
rect 35345 6675 35403 6681
rect 35618 6672 35624 6684
rect 35676 6672 35682 6724
rect 35802 6672 35808 6724
rect 35860 6712 35866 6724
rect 45572 6712 45600 6752
rect 48222 6740 48228 6752
rect 48280 6740 48286 6792
rect 56870 6780 56876 6792
rect 56831 6752 56876 6780
rect 56870 6740 56876 6752
rect 56928 6740 56934 6792
rect 56962 6740 56968 6792
rect 57020 6780 57026 6792
rect 57129 6783 57187 6789
rect 57129 6780 57141 6783
rect 57020 6752 57141 6780
rect 57020 6740 57026 6752
rect 57129 6749 57141 6752
rect 57175 6749 57187 6783
rect 57129 6743 57187 6749
rect 35860 6684 45600 6712
rect 46201 6715 46259 6721
rect 35860 6672 35866 6684
rect 46201 6681 46213 6715
rect 46247 6712 46259 6715
rect 58710 6712 58716 6724
rect 46247 6684 58716 6712
rect 46247 6681 46259 6684
rect 46201 6675 46259 6681
rect 58710 6672 58716 6684
rect 58768 6672 58774 6724
rect 31435 6616 32904 6644
rect 31435 6613 31447 6616
rect 31389 6607 31447 6613
rect 33042 6604 33048 6656
rect 33100 6644 33106 6656
rect 35253 6647 35311 6653
rect 35253 6644 35265 6647
rect 33100 6616 35265 6644
rect 33100 6604 33106 6616
rect 35253 6613 35265 6616
rect 35299 6644 35311 6647
rect 35894 6644 35900 6656
rect 35299 6616 35900 6644
rect 35299 6613 35311 6616
rect 35253 6607 35311 6613
rect 35894 6604 35900 6616
rect 35952 6604 35958 6656
rect 36446 6604 36452 6656
rect 36504 6644 36510 6656
rect 36722 6644 36728 6656
rect 36504 6616 36728 6644
rect 36504 6604 36510 6616
rect 36722 6604 36728 6616
rect 36780 6604 36786 6656
rect 57974 6604 57980 6656
rect 58032 6644 58038 6656
rect 58250 6644 58256 6656
rect 58032 6616 58256 6644
rect 58032 6604 58038 6616
rect 58250 6604 58256 6616
rect 58308 6604 58314 6656
rect 1104 6554 58880 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 58880 6554
rect 1104 6480 58880 6502
rect 9122 6440 9128 6452
rect 9083 6412 9128 6440
rect 9122 6400 9128 6412
rect 9180 6400 9186 6452
rect 14369 6443 14427 6449
rect 14369 6409 14381 6443
rect 14415 6409 14427 6443
rect 14369 6403 14427 6409
rect 10870 6372 10876 6384
rect 9324 6344 10876 6372
rect 9324 6316 9352 6344
rect 10870 6332 10876 6344
rect 10928 6332 10934 6384
rect 11698 6332 11704 6384
rect 11756 6372 11762 6384
rect 13541 6375 13599 6381
rect 13541 6372 13553 6375
rect 11756 6344 13553 6372
rect 11756 6332 11762 6344
rect 13541 6341 13553 6344
rect 13587 6372 13599 6375
rect 14384 6372 14412 6403
rect 17862 6400 17868 6452
rect 17920 6440 17926 6452
rect 24670 6440 24676 6452
rect 17920 6412 23339 6440
rect 24631 6412 24676 6440
rect 17920 6400 17926 6412
rect 13587 6344 14412 6372
rect 13587 6341 13599 6344
rect 13541 6335 13599 6341
rect 15378 6332 15384 6384
rect 15436 6372 15442 6384
rect 15436 6344 15481 6372
rect 15436 6332 15442 6344
rect 15654 6332 15660 6384
rect 15712 6372 15718 6384
rect 15712 6344 16344 6372
rect 15712 6332 15718 6344
rect 1581 6307 1639 6313
rect 1581 6273 1593 6307
rect 1627 6304 1639 6307
rect 9122 6304 9128 6316
rect 1627 6276 9128 6304
rect 1627 6273 1639 6276
rect 1581 6267 1639 6273
rect 9122 6264 9128 6276
rect 9180 6264 9186 6316
rect 9306 6304 9312 6316
rect 9219 6276 9312 6304
rect 9306 6264 9312 6276
rect 9364 6264 9370 6316
rect 9401 6307 9459 6313
rect 9401 6273 9413 6307
rect 9447 6304 9459 6307
rect 14277 6307 14335 6313
rect 9447 6276 14228 6304
rect 9447 6273 9459 6276
rect 9401 6267 9459 6273
rect 1762 6236 1768 6248
rect 1723 6208 1768 6236
rect 1762 6196 1768 6208
rect 1820 6196 1826 6248
rect 8938 6196 8944 6248
rect 8996 6236 9002 6248
rect 9490 6236 9496 6248
rect 8996 6208 9496 6236
rect 8996 6196 9002 6208
rect 9490 6196 9496 6208
rect 9548 6196 9554 6248
rect 9582 6196 9588 6248
rect 9640 6236 9646 6248
rect 9640 6208 9685 6236
rect 9640 6196 9646 6208
rect 12434 6128 12440 6180
rect 12492 6168 12498 6180
rect 13722 6168 13728 6180
rect 12492 6140 13728 6168
rect 12492 6128 12498 6140
rect 13722 6128 13728 6140
rect 13780 6128 13786 6180
rect 14200 6168 14228 6276
rect 14277 6273 14289 6307
rect 14323 6304 14335 6307
rect 15194 6304 15200 6316
rect 14323 6276 15200 6304
rect 14323 6273 14335 6276
rect 14277 6267 14335 6273
rect 15194 6264 15200 6276
rect 15252 6264 15258 6316
rect 15289 6307 15347 6313
rect 15289 6273 15301 6307
rect 15335 6304 15347 6307
rect 15470 6304 15476 6316
rect 15335 6276 15476 6304
rect 15335 6273 15347 6276
rect 15289 6267 15347 6273
rect 15470 6264 15476 6276
rect 15528 6264 15534 6316
rect 15746 6304 15752 6316
rect 15659 6276 15752 6304
rect 15746 6264 15752 6276
rect 15804 6264 15810 6316
rect 15841 6307 15899 6313
rect 15841 6273 15853 6307
rect 15887 6304 15899 6307
rect 16206 6304 16212 6316
rect 15887 6276 16212 6304
rect 15887 6273 15899 6276
rect 15841 6267 15899 6273
rect 16206 6264 16212 6276
rect 16264 6264 16270 6316
rect 16316 6313 16344 6344
rect 17770 6332 17776 6384
rect 17828 6372 17834 6384
rect 18233 6375 18291 6381
rect 18233 6372 18245 6375
rect 17828 6344 18245 6372
rect 17828 6332 17834 6344
rect 18233 6341 18245 6344
rect 18279 6341 18291 6375
rect 18233 6335 18291 6341
rect 18506 6332 18512 6384
rect 18564 6372 18570 6384
rect 19518 6372 19524 6384
rect 18564 6344 19524 6372
rect 18564 6332 18570 6344
rect 19518 6332 19524 6344
rect 19576 6332 19582 6384
rect 19794 6332 19800 6384
rect 19852 6372 19858 6384
rect 19852 6344 22784 6372
rect 19852 6332 19858 6344
rect 16301 6307 16359 6313
rect 16301 6273 16313 6307
rect 16347 6304 16359 6307
rect 17034 6304 17040 6316
rect 16347 6276 17040 6304
rect 16347 6273 16359 6276
rect 16301 6267 16359 6273
rect 17034 6264 17040 6276
rect 17092 6264 17098 6316
rect 17497 6307 17555 6313
rect 17497 6273 17509 6307
rect 17543 6304 17555 6307
rect 17954 6304 17960 6316
rect 17543 6276 17960 6304
rect 17543 6273 17555 6276
rect 17497 6267 17555 6273
rect 17954 6264 17960 6276
rect 18012 6304 18018 6316
rect 19242 6304 19248 6316
rect 18012 6276 19248 6304
rect 18012 6264 18018 6276
rect 19242 6264 19248 6276
rect 19300 6264 19306 6316
rect 19334 6264 19340 6316
rect 19392 6304 19398 6316
rect 19685 6307 19743 6313
rect 19685 6304 19697 6307
rect 19392 6276 19697 6304
rect 19392 6264 19398 6276
rect 19685 6273 19697 6276
rect 19731 6273 19743 6307
rect 19685 6267 19743 6273
rect 22373 6307 22431 6313
rect 22373 6273 22385 6307
rect 22419 6304 22431 6307
rect 22646 6304 22652 6316
rect 22419 6276 22652 6304
rect 22419 6273 22431 6276
rect 22373 6267 22431 6273
rect 22646 6264 22652 6276
rect 22704 6264 22710 6316
rect 15764 6236 15792 6264
rect 16390 6236 16396 6248
rect 15764 6208 16396 6236
rect 16390 6196 16396 6208
rect 16448 6196 16454 6248
rect 18506 6196 18512 6248
rect 18564 6236 18570 6248
rect 18782 6236 18788 6248
rect 18564 6208 18788 6236
rect 18564 6196 18570 6208
rect 18782 6196 18788 6208
rect 18840 6196 18846 6248
rect 19426 6236 19432 6248
rect 19387 6208 19432 6236
rect 19426 6196 19432 6208
rect 19484 6196 19490 6248
rect 18690 6168 18696 6180
rect 14200 6140 18696 6168
rect 18690 6128 18696 6140
rect 18748 6128 18754 6180
rect 21358 6128 21364 6180
rect 21416 6168 21422 6180
rect 22557 6171 22615 6177
rect 22557 6168 22569 6171
rect 21416 6140 22569 6168
rect 21416 6128 21422 6140
rect 22557 6137 22569 6140
rect 22603 6137 22615 6171
rect 22557 6131 22615 6137
rect 9398 6060 9404 6112
rect 9456 6100 9462 6112
rect 20714 6100 20720 6112
rect 9456 6072 20720 6100
rect 9456 6060 9462 6072
rect 20714 6060 20720 6072
rect 20772 6060 20778 6112
rect 20809 6103 20867 6109
rect 20809 6069 20821 6103
rect 20855 6100 20867 6103
rect 21450 6100 21456 6112
rect 20855 6072 21456 6100
rect 20855 6069 20867 6072
rect 20809 6063 20867 6069
rect 21450 6060 21456 6072
rect 21508 6060 21514 6112
rect 22756 6100 22784 6344
rect 23311 6304 23339 6412
rect 24670 6400 24676 6412
rect 24728 6400 24734 6452
rect 25590 6440 25596 6452
rect 25551 6412 25596 6440
rect 25590 6400 25596 6412
rect 25648 6400 25654 6452
rect 25682 6400 25688 6452
rect 25740 6440 25746 6452
rect 28258 6440 28264 6452
rect 25740 6412 28264 6440
rect 25740 6400 25746 6412
rect 28258 6400 28264 6412
rect 28316 6400 28322 6452
rect 30469 6443 30527 6449
rect 30469 6409 30481 6443
rect 30515 6440 30527 6443
rect 30558 6440 30564 6452
rect 30515 6412 30564 6440
rect 30515 6409 30527 6412
rect 30469 6403 30527 6409
rect 30558 6400 30564 6412
rect 30616 6400 30622 6452
rect 33778 6400 33784 6452
rect 33836 6440 33842 6452
rect 37645 6443 37703 6449
rect 37645 6440 37657 6443
rect 33836 6412 37657 6440
rect 33836 6400 33842 6412
rect 37645 6409 37657 6412
rect 37691 6409 37703 6443
rect 46750 6440 46756 6452
rect 46711 6412 46756 6440
rect 37645 6403 37703 6409
rect 46750 6400 46756 6412
rect 46808 6400 46814 6452
rect 23385 6375 23443 6381
rect 23385 6341 23397 6375
rect 23431 6372 23443 6375
rect 28626 6372 28632 6384
rect 23431 6344 28632 6372
rect 23431 6341 23443 6344
rect 23385 6335 23443 6341
rect 28626 6332 28632 6344
rect 28684 6332 28690 6384
rect 33686 6372 33692 6384
rect 28966 6344 33692 6372
rect 23311 6276 23428 6304
rect 23400 6168 23428 6276
rect 25038 6264 25044 6316
rect 25096 6304 25102 6316
rect 25961 6307 26019 6313
rect 25961 6304 25973 6307
rect 25096 6276 25973 6304
rect 25096 6264 25102 6276
rect 25961 6273 25973 6276
rect 26007 6273 26019 6307
rect 25961 6267 26019 6273
rect 26234 6264 26240 6316
rect 26292 6304 26298 6316
rect 26602 6304 26608 6316
rect 26292 6276 26608 6304
rect 26292 6264 26298 6276
rect 26602 6264 26608 6276
rect 26660 6264 26666 6316
rect 27154 6304 27160 6316
rect 27115 6276 27160 6304
rect 27154 6264 27160 6276
rect 27212 6264 27218 6316
rect 28966 6304 28994 6344
rect 33686 6332 33692 6344
rect 33744 6332 33750 6384
rect 51350 6372 51356 6384
rect 46492 6344 51356 6372
rect 27264 6276 28994 6304
rect 29089 6307 29147 6313
rect 26050 6236 26056 6248
rect 26011 6208 26056 6236
rect 26050 6196 26056 6208
rect 26108 6196 26114 6248
rect 26145 6239 26203 6245
rect 26145 6205 26157 6239
rect 26191 6236 26203 6239
rect 26418 6236 26424 6248
rect 26191 6208 26424 6236
rect 26191 6205 26203 6208
rect 26145 6199 26203 6205
rect 26418 6196 26424 6208
rect 26476 6236 26482 6248
rect 26878 6236 26884 6248
rect 26476 6208 26884 6236
rect 26476 6196 26482 6208
rect 26878 6196 26884 6208
rect 26936 6196 26942 6248
rect 27264 6168 27292 6276
rect 29089 6273 29101 6307
rect 29135 6273 29147 6307
rect 29089 6267 29147 6273
rect 27433 6239 27491 6245
rect 27433 6205 27445 6239
rect 27479 6236 27491 6239
rect 27522 6236 27528 6248
rect 27479 6208 27528 6236
rect 27479 6205 27491 6208
rect 27433 6199 27491 6205
rect 27522 6196 27528 6208
rect 27580 6196 27586 6248
rect 29104 6236 29132 6267
rect 30558 6264 30564 6316
rect 30616 6304 30622 6316
rect 32122 6304 32128 6316
rect 30616 6276 32128 6304
rect 30616 6264 30622 6276
rect 32122 6264 32128 6276
rect 32180 6264 32186 6316
rect 33870 6264 33876 6316
rect 33928 6304 33934 6316
rect 34517 6307 34575 6313
rect 33928 6276 33973 6304
rect 33928 6264 33934 6276
rect 34517 6273 34529 6307
rect 34563 6304 34575 6307
rect 34606 6304 34612 6316
rect 34563 6276 34612 6304
rect 34563 6273 34575 6276
rect 34517 6267 34575 6273
rect 34606 6264 34612 6276
rect 34664 6264 34670 6316
rect 35434 6264 35440 6316
rect 35492 6304 35498 6316
rect 35529 6307 35587 6313
rect 35529 6304 35541 6307
rect 35492 6276 35541 6304
rect 35492 6264 35498 6276
rect 35529 6273 35541 6276
rect 35575 6273 35587 6307
rect 35894 6304 35900 6316
rect 35855 6276 35900 6304
rect 35529 6267 35587 6273
rect 35894 6264 35900 6276
rect 35952 6264 35958 6316
rect 36449 6307 36507 6313
rect 36449 6273 36461 6307
rect 36495 6273 36507 6307
rect 36449 6267 36507 6273
rect 27623 6208 32904 6236
rect 27623 6168 27651 6208
rect 23400 6140 27292 6168
rect 27356 6140 27651 6168
rect 27709 6171 27767 6177
rect 27356 6100 27384 6140
rect 27709 6137 27721 6171
rect 27755 6168 27767 6171
rect 32766 6168 32772 6180
rect 27755 6140 32772 6168
rect 27755 6137 27767 6140
rect 27709 6131 27767 6137
rect 32766 6128 32772 6140
rect 32824 6128 32830 6180
rect 32876 6168 32904 6208
rect 33134 6196 33140 6248
rect 33192 6236 33198 6248
rect 34701 6239 34759 6245
rect 34701 6236 34713 6239
rect 33192 6208 34713 6236
rect 33192 6196 33198 6208
rect 34701 6205 34713 6208
rect 34747 6205 34759 6239
rect 34701 6199 34759 6205
rect 35802 6196 35808 6248
rect 35860 6236 35866 6248
rect 36464 6236 36492 6267
rect 37274 6264 37280 6316
rect 37332 6304 37338 6316
rect 46492 6313 46520 6344
rect 51350 6332 51356 6344
rect 51408 6332 51414 6384
rect 57146 6372 57152 6384
rect 57107 6344 57152 6372
rect 57146 6332 57152 6344
rect 57204 6332 57210 6384
rect 37553 6307 37611 6313
rect 37553 6304 37565 6307
rect 37332 6276 37565 6304
rect 37332 6264 37338 6276
rect 37553 6273 37565 6276
rect 37599 6273 37611 6307
rect 37553 6267 37611 6273
rect 46477 6307 46535 6313
rect 46477 6273 46489 6307
rect 46523 6273 46535 6307
rect 46477 6267 46535 6273
rect 46569 6307 46627 6313
rect 46569 6273 46581 6307
rect 46615 6304 46627 6307
rect 46842 6304 46848 6316
rect 46615 6276 46848 6304
rect 46615 6273 46627 6276
rect 46569 6267 46627 6273
rect 46842 6264 46848 6276
rect 46900 6264 46906 6316
rect 35860 6208 36860 6236
rect 35860 6196 35866 6208
rect 33318 6168 33324 6180
rect 32876 6140 33324 6168
rect 33318 6128 33324 6140
rect 33376 6128 33382 6180
rect 34057 6171 34115 6177
rect 34057 6137 34069 6171
rect 34103 6168 34115 6171
rect 36262 6168 36268 6180
rect 34103 6140 36268 6168
rect 34103 6137 34115 6140
rect 34057 6131 34115 6137
rect 36262 6128 36268 6140
rect 36320 6128 36326 6180
rect 22756 6072 27384 6100
rect 27522 6060 27528 6112
rect 27580 6100 27586 6112
rect 27580 6072 27625 6100
rect 27580 6060 27586 6072
rect 29086 6060 29092 6112
rect 29144 6100 29150 6112
rect 35434 6100 35440 6112
rect 29144 6072 35440 6100
rect 29144 6060 29150 6072
rect 35434 6060 35440 6072
rect 35492 6060 35498 6112
rect 35894 6060 35900 6112
rect 35952 6100 35958 6112
rect 36541 6103 36599 6109
rect 36541 6100 36553 6103
rect 35952 6072 36553 6100
rect 35952 6060 35958 6072
rect 36541 6069 36553 6072
rect 36587 6069 36599 6103
rect 36832 6100 36860 6208
rect 36906 6128 36912 6180
rect 36964 6168 36970 6180
rect 36964 6140 55214 6168
rect 36964 6128 36970 6140
rect 39298 6100 39304 6112
rect 36832 6072 39304 6100
rect 36541 6063 36599 6069
rect 39298 6060 39304 6072
rect 39356 6060 39362 6112
rect 55186 6100 55214 6140
rect 57241 6103 57299 6109
rect 57241 6100 57253 6103
rect 55186 6072 57253 6100
rect 57241 6069 57253 6072
rect 57287 6069 57299 6103
rect 57241 6063 57299 6069
rect 1104 6010 58880 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 58880 6010
rect 1104 5936 58880 5958
rect 9122 5896 9128 5908
rect 9083 5868 9128 5896
rect 9122 5856 9128 5868
rect 9180 5856 9186 5908
rect 10873 5899 10931 5905
rect 9232 5868 10824 5896
rect 7926 5788 7932 5840
rect 7984 5828 7990 5840
rect 9232 5828 9260 5868
rect 7984 5800 9260 5828
rect 10689 5831 10747 5837
rect 7984 5788 7990 5800
rect 10689 5797 10701 5831
rect 10735 5797 10747 5831
rect 10689 5791 10747 5797
rect 9398 5760 9404 5772
rect 9359 5732 9404 5760
rect 9398 5720 9404 5732
rect 9456 5720 9462 5772
rect 9493 5763 9551 5769
rect 9493 5729 9505 5763
rect 9539 5760 9551 5763
rect 9674 5760 9680 5772
rect 9539 5732 9680 5760
rect 9539 5729 9551 5732
rect 9493 5723 9551 5729
rect 9674 5720 9680 5732
rect 9732 5760 9738 5772
rect 9732 5732 9825 5760
rect 9732 5720 9738 5732
rect 1581 5695 1639 5701
rect 1581 5661 1593 5695
rect 1627 5692 1639 5695
rect 9306 5692 9312 5704
rect 1627 5664 2774 5692
rect 9267 5664 9312 5692
rect 1627 5661 1639 5664
rect 1581 5655 1639 5661
rect 1854 5624 1860 5636
rect 1815 5596 1860 5624
rect 1854 5584 1860 5596
rect 1912 5584 1918 5636
rect 2746 5624 2774 5664
rect 9306 5652 9312 5664
rect 9364 5652 9370 5704
rect 9582 5652 9588 5704
rect 9640 5692 9646 5704
rect 9784 5692 9812 5732
rect 9640 5664 9685 5692
rect 9784 5664 10456 5692
rect 9640 5652 9646 5664
rect 10428 5636 10456 5664
rect 10134 5624 10140 5636
rect 2746 5596 10140 5624
rect 10134 5584 10140 5596
rect 10192 5584 10198 5636
rect 10410 5624 10416 5636
rect 10371 5596 10416 5624
rect 10410 5584 10416 5596
rect 10468 5584 10474 5636
rect 7742 5516 7748 5568
rect 7800 5556 7806 5568
rect 10704 5556 10732 5791
rect 10796 5760 10824 5868
rect 10873 5865 10885 5899
rect 10919 5896 10931 5899
rect 11054 5896 11060 5908
rect 10919 5868 11060 5896
rect 10919 5865 10931 5868
rect 10873 5859 10931 5865
rect 11054 5856 11060 5868
rect 11112 5856 11118 5908
rect 12618 5856 12624 5908
rect 12676 5896 12682 5908
rect 13725 5899 13783 5905
rect 13725 5896 13737 5899
rect 12676 5868 13737 5896
rect 12676 5856 12682 5868
rect 13725 5865 13737 5868
rect 13771 5865 13783 5899
rect 13725 5859 13783 5865
rect 13814 5856 13820 5908
rect 13872 5896 13878 5908
rect 23017 5899 23075 5905
rect 13872 5868 22968 5896
rect 13872 5856 13878 5868
rect 11882 5788 11888 5840
rect 11940 5828 11946 5840
rect 13541 5831 13599 5837
rect 13541 5828 13553 5831
rect 11940 5800 13553 5828
rect 11940 5788 11946 5800
rect 13541 5797 13553 5800
rect 13587 5797 13599 5831
rect 13541 5791 13599 5797
rect 14553 5831 14611 5837
rect 14553 5797 14565 5831
rect 14599 5797 14611 5831
rect 14553 5791 14611 5797
rect 10796 5732 12434 5760
rect 12406 5692 12434 5732
rect 14568 5692 14596 5791
rect 16206 5788 16212 5840
rect 16264 5788 16270 5840
rect 16850 5788 16856 5840
rect 16908 5828 16914 5840
rect 19610 5828 19616 5840
rect 16908 5800 19616 5828
rect 16908 5788 16914 5800
rect 19610 5788 19616 5800
rect 19668 5788 19674 5840
rect 22940 5828 22968 5868
rect 23017 5865 23029 5899
rect 23063 5896 23075 5899
rect 23106 5896 23112 5908
rect 23063 5868 23112 5896
rect 23063 5865 23075 5868
rect 23017 5859 23075 5865
rect 23106 5856 23112 5868
rect 23164 5856 23170 5908
rect 23382 5856 23388 5908
rect 23440 5896 23446 5908
rect 26145 5899 26203 5905
rect 26145 5896 26157 5899
rect 23440 5868 26157 5896
rect 23440 5856 23446 5868
rect 26145 5865 26157 5868
rect 26191 5865 26203 5899
rect 26145 5859 26203 5865
rect 26234 5856 26240 5908
rect 26292 5896 26298 5908
rect 29638 5896 29644 5908
rect 26292 5868 29644 5896
rect 26292 5856 26298 5868
rect 29638 5856 29644 5868
rect 29696 5856 29702 5908
rect 29730 5856 29736 5908
rect 29788 5896 29794 5908
rect 29898 5899 29956 5905
rect 29898 5896 29910 5899
rect 29788 5868 29910 5896
rect 29788 5856 29794 5868
rect 29898 5865 29910 5868
rect 29944 5865 29956 5899
rect 29898 5859 29956 5865
rect 30006 5856 30012 5908
rect 30064 5896 30070 5908
rect 48314 5896 48320 5908
rect 30064 5868 30109 5896
rect 37752 5868 48320 5896
rect 30064 5856 30070 5868
rect 22940 5800 23888 5828
rect 15654 5760 15660 5772
rect 15615 5732 15660 5760
rect 15654 5720 15660 5732
rect 15712 5720 15718 5772
rect 15749 5763 15807 5769
rect 15749 5729 15761 5763
rect 15795 5760 15807 5763
rect 15838 5760 15844 5772
rect 15795 5732 15844 5760
rect 15795 5729 15807 5732
rect 15749 5723 15807 5729
rect 15838 5720 15844 5732
rect 15896 5720 15902 5772
rect 12406 5664 14596 5692
rect 15470 5652 15476 5704
rect 15528 5692 15534 5704
rect 16224 5701 16252 5788
rect 16868 5732 17172 5760
rect 16390 5701 16396 5704
rect 16117 5695 16175 5701
rect 16117 5692 16129 5695
rect 15528 5664 16129 5692
rect 15528 5652 15534 5664
rect 16117 5661 16129 5664
rect 16163 5661 16175 5695
rect 16117 5655 16175 5661
rect 16205 5695 16263 5701
rect 16205 5661 16217 5695
rect 16251 5661 16263 5695
rect 16205 5655 16263 5661
rect 16347 5695 16396 5701
rect 16347 5661 16359 5695
rect 16393 5661 16396 5695
rect 16347 5655 16396 5661
rect 16390 5652 16396 5655
rect 16448 5692 16454 5704
rect 16868 5692 16896 5732
rect 17034 5692 17040 5704
rect 16448 5664 16896 5692
rect 16995 5664 17040 5692
rect 16448 5652 16454 5664
rect 17034 5652 17040 5664
rect 17092 5652 17098 5704
rect 17144 5692 17172 5732
rect 17402 5720 17408 5772
rect 17460 5760 17466 5772
rect 17460 5732 17908 5760
rect 17460 5720 17466 5732
rect 17589 5695 17647 5701
rect 17589 5692 17601 5695
rect 17144 5664 17601 5692
rect 17589 5661 17601 5664
rect 17635 5692 17647 5695
rect 17770 5692 17776 5704
rect 17635 5664 17776 5692
rect 17635 5661 17647 5664
rect 17589 5655 17647 5661
rect 17770 5652 17776 5664
rect 17828 5652 17834 5704
rect 17880 5701 17908 5732
rect 18138 5720 18144 5772
rect 18196 5760 18202 5772
rect 21637 5763 21695 5769
rect 21637 5760 21649 5763
rect 18196 5732 19748 5760
rect 18196 5720 18202 5732
rect 17865 5695 17923 5701
rect 17865 5661 17877 5695
rect 17911 5661 17923 5695
rect 17865 5655 17923 5661
rect 18601 5695 18659 5701
rect 18601 5661 18613 5695
rect 18647 5692 18659 5695
rect 18966 5692 18972 5704
rect 18647 5664 18972 5692
rect 18647 5661 18659 5664
rect 18601 5655 18659 5661
rect 18966 5652 18972 5664
rect 19024 5652 19030 5704
rect 19426 5652 19432 5704
rect 19484 5692 19490 5704
rect 19610 5692 19616 5704
rect 19484 5664 19616 5692
rect 19484 5652 19490 5664
rect 19610 5652 19616 5664
rect 19668 5652 19674 5704
rect 19720 5692 19748 5732
rect 20640 5732 21649 5760
rect 19869 5695 19927 5701
rect 19869 5692 19881 5695
rect 19720 5664 19881 5692
rect 19869 5661 19881 5664
rect 19915 5661 19927 5695
rect 19869 5655 19927 5661
rect 20254 5652 20260 5704
rect 20312 5692 20318 5704
rect 20640 5692 20668 5732
rect 21637 5729 21649 5732
rect 21683 5729 21695 5763
rect 21637 5723 21695 5729
rect 23106 5720 23112 5772
rect 23164 5760 23170 5772
rect 23569 5763 23627 5769
rect 23164 5732 23336 5760
rect 23164 5720 23170 5732
rect 21450 5692 21456 5704
rect 20312 5664 20668 5692
rect 21411 5664 21456 5692
rect 20312 5652 20318 5664
rect 21450 5652 21456 5664
rect 21508 5652 21514 5704
rect 22557 5695 22615 5701
rect 22557 5661 22569 5695
rect 22603 5692 22615 5695
rect 23198 5692 23204 5704
rect 22603 5664 23204 5692
rect 22603 5661 22615 5664
rect 22557 5655 22615 5661
rect 23198 5652 23204 5664
rect 23256 5652 23262 5704
rect 23308 5692 23336 5732
rect 23569 5729 23581 5763
rect 23615 5729 23627 5763
rect 23860 5760 23888 5800
rect 26602 5788 26608 5840
rect 26660 5828 26666 5840
rect 28902 5828 28908 5840
rect 26660 5800 28908 5828
rect 26660 5788 26666 5800
rect 28902 5788 28908 5800
rect 28960 5828 28966 5840
rect 35802 5828 35808 5840
rect 28960 5800 29960 5828
rect 28960 5788 28966 5800
rect 23860 5732 29868 5760
rect 23569 5723 23627 5729
rect 23477 5695 23535 5701
rect 23477 5692 23489 5695
rect 23308 5664 23489 5692
rect 23477 5661 23489 5664
rect 23523 5661 23535 5695
rect 23477 5655 23535 5661
rect 13265 5627 13323 5633
rect 13265 5593 13277 5627
rect 13311 5624 13323 5627
rect 14274 5624 14280 5636
rect 13311 5596 14280 5624
rect 13311 5593 13323 5596
rect 13265 5587 13323 5593
rect 14274 5584 14280 5596
rect 14332 5584 14338 5636
rect 15562 5624 15568 5636
rect 14660 5596 15568 5624
rect 7800 5528 10732 5556
rect 7800 5516 7806 5528
rect 13906 5516 13912 5568
rect 13964 5556 13970 5568
rect 14660 5556 14688 5596
rect 15562 5584 15568 5596
rect 15620 5624 15626 5636
rect 16850 5624 16856 5636
rect 15620 5596 16856 5624
rect 15620 5584 15626 5596
rect 16850 5584 16856 5596
rect 16908 5584 16914 5636
rect 23290 5624 23296 5636
rect 16960 5596 23296 5624
rect 13964 5528 14688 5556
rect 14737 5559 14795 5565
rect 13964 5516 13970 5528
rect 14737 5525 14749 5559
rect 14783 5556 14795 5559
rect 16960 5556 16988 5596
rect 23290 5584 23296 5596
rect 23348 5584 23354 5636
rect 14783 5528 16988 5556
rect 18325 5559 18383 5565
rect 14783 5525 14795 5528
rect 14737 5519 14795 5525
rect 18325 5525 18337 5559
rect 18371 5556 18383 5559
rect 18506 5556 18512 5568
rect 18371 5528 18512 5556
rect 18371 5525 18383 5528
rect 18325 5519 18383 5525
rect 18506 5516 18512 5528
rect 18564 5516 18570 5568
rect 18598 5516 18604 5568
rect 18656 5556 18662 5568
rect 20993 5559 21051 5565
rect 20993 5556 21005 5559
rect 18656 5528 21005 5556
rect 18656 5516 18662 5528
rect 20993 5525 21005 5528
rect 21039 5525 21051 5559
rect 20993 5519 21051 5525
rect 21082 5516 21088 5568
rect 21140 5556 21146 5568
rect 23385 5559 23443 5565
rect 23385 5556 23397 5559
rect 21140 5528 23397 5556
rect 21140 5516 21146 5528
rect 23385 5525 23397 5528
rect 23431 5525 23443 5559
rect 23584 5556 23612 5723
rect 24854 5652 24860 5704
rect 24912 5692 24918 5704
rect 24949 5695 25007 5701
rect 24949 5692 24961 5695
rect 24912 5664 24961 5692
rect 24912 5652 24918 5664
rect 24949 5661 24961 5664
rect 24995 5661 25007 5695
rect 24949 5655 25007 5661
rect 26602 5652 26608 5704
rect 26660 5692 26666 5704
rect 27893 5695 27951 5701
rect 27893 5692 27905 5695
rect 26660 5664 27905 5692
rect 26660 5652 26666 5664
rect 27893 5661 27905 5664
rect 27939 5661 27951 5695
rect 28534 5692 28540 5704
rect 28495 5664 28540 5692
rect 27893 5655 27951 5661
rect 28534 5652 28540 5664
rect 28592 5652 28598 5704
rect 28810 5652 28816 5704
rect 28868 5692 28874 5704
rect 28905 5695 28963 5701
rect 28905 5692 28917 5695
rect 28868 5664 28917 5692
rect 28868 5652 28874 5664
rect 28905 5661 28917 5664
rect 28951 5661 28963 5695
rect 28905 5655 28963 5661
rect 23658 5584 23664 5636
rect 23716 5624 23722 5636
rect 28718 5624 28724 5636
rect 23716 5596 28724 5624
rect 23716 5584 23722 5596
rect 28718 5584 28724 5596
rect 28776 5584 28782 5636
rect 29733 5627 29791 5633
rect 29733 5593 29745 5627
rect 29779 5593 29791 5627
rect 29840 5624 29868 5732
rect 29932 5692 29960 5800
rect 34164 5800 35808 5828
rect 30098 5760 30104 5772
rect 30059 5732 30104 5760
rect 30098 5720 30104 5732
rect 30156 5720 30162 5772
rect 30190 5720 30196 5772
rect 30248 5760 30254 5772
rect 31205 5763 31263 5769
rect 31205 5760 31217 5763
rect 30248 5732 31217 5760
rect 30248 5720 30254 5732
rect 31205 5729 31217 5732
rect 31251 5729 31263 5763
rect 31205 5723 31263 5729
rect 30469 5695 30527 5701
rect 30469 5692 30481 5695
rect 29932 5664 30481 5692
rect 30469 5661 30481 5664
rect 30515 5661 30527 5695
rect 30469 5655 30527 5661
rect 31472 5695 31530 5701
rect 31472 5661 31484 5695
rect 31518 5692 31530 5695
rect 32950 5692 32956 5704
rect 31518 5664 32956 5692
rect 31518 5661 31530 5664
rect 31472 5655 31530 5661
rect 32950 5652 32956 5664
rect 33008 5652 33014 5704
rect 33413 5695 33471 5701
rect 33413 5661 33425 5695
rect 33459 5692 33471 5695
rect 33778 5692 33784 5704
rect 33459 5664 33784 5692
rect 33459 5661 33471 5664
rect 33413 5655 33471 5661
rect 33778 5652 33784 5664
rect 33836 5692 33842 5704
rect 34164 5701 34192 5800
rect 35802 5788 35808 5800
rect 35860 5788 35866 5840
rect 35989 5831 36047 5837
rect 35989 5797 36001 5831
rect 36035 5828 36047 5831
rect 37642 5828 37648 5840
rect 36035 5800 37648 5828
rect 36035 5797 36047 5800
rect 35989 5791 36047 5797
rect 37642 5788 37648 5800
rect 37700 5788 37706 5840
rect 35342 5720 35348 5772
rect 35400 5760 35406 5772
rect 36541 5763 36599 5769
rect 36541 5760 36553 5763
rect 35400 5732 36553 5760
rect 35400 5720 35406 5732
rect 36541 5729 36553 5732
rect 36587 5729 36599 5763
rect 37752 5760 37780 5868
rect 48314 5856 48320 5868
rect 48372 5856 48378 5908
rect 38378 5828 38384 5840
rect 38339 5800 38384 5828
rect 38378 5788 38384 5800
rect 38436 5788 38442 5840
rect 40313 5831 40371 5837
rect 40313 5797 40325 5831
rect 40359 5828 40371 5831
rect 40494 5828 40500 5840
rect 40359 5800 40500 5828
rect 40359 5797 40371 5800
rect 40313 5791 40371 5797
rect 40494 5788 40500 5800
rect 40552 5788 40558 5840
rect 41414 5788 41420 5840
rect 41472 5828 41478 5840
rect 41601 5831 41659 5837
rect 41601 5828 41613 5831
rect 41472 5800 41613 5828
rect 41472 5788 41478 5800
rect 41601 5797 41613 5800
rect 41647 5797 41659 5831
rect 41601 5791 41659 5797
rect 36541 5723 36599 5729
rect 36648 5732 37780 5760
rect 34149 5695 34207 5701
rect 34149 5692 34161 5695
rect 33836 5664 34161 5692
rect 33836 5652 33842 5664
rect 34149 5661 34161 5664
rect 34195 5661 34207 5695
rect 34149 5655 34207 5661
rect 34790 5652 34796 5704
rect 34848 5692 34854 5704
rect 34977 5695 35035 5701
rect 34977 5692 34989 5695
rect 34848 5664 34989 5692
rect 34848 5652 34854 5664
rect 34977 5661 34989 5664
rect 35023 5661 35035 5695
rect 34977 5655 35035 5661
rect 35434 5652 35440 5704
rect 35492 5692 35498 5704
rect 35713 5695 35771 5701
rect 35713 5692 35725 5695
rect 35492 5664 35725 5692
rect 35492 5652 35498 5664
rect 35713 5661 35725 5664
rect 35759 5692 35771 5695
rect 36449 5695 36507 5701
rect 36449 5692 36461 5695
rect 35759 5664 36461 5692
rect 35759 5661 35771 5664
rect 35713 5655 35771 5661
rect 36449 5661 36461 5664
rect 36495 5692 36507 5695
rect 36648 5692 36676 5732
rect 36495 5664 36676 5692
rect 36495 5661 36507 5664
rect 36449 5655 36507 5661
rect 37366 5652 37372 5704
rect 37424 5692 37430 5704
rect 37461 5695 37519 5701
rect 37461 5692 37473 5695
rect 37424 5664 37473 5692
rect 37424 5652 37430 5664
rect 37461 5661 37473 5664
rect 37507 5661 37519 5695
rect 37461 5655 37519 5661
rect 37645 5695 37703 5701
rect 37645 5661 37657 5695
rect 37691 5692 37703 5695
rect 37734 5692 37740 5704
rect 37691 5664 37740 5692
rect 37691 5661 37703 5664
rect 37645 5655 37703 5661
rect 37734 5652 37740 5664
rect 37792 5652 37798 5704
rect 38396 5692 38424 5788
rect 38562 5720 38568 5772
rect 38620 5760 38626 5772
rect 39301 5763 39359 5769
rect 39301 5760 39313 5763
rect 38620 5732 39313 5760
rect 38620 5720 38626 5732
rect 39301 5729 39313 5732
rect 39347 5729 39359 5763
rect 57974 5760 57980 5772
rect 39301 5723 39359 5729
rect 56980 5732 57980 5760
rect 55858 5692 55864 5704
rect 38396 5664 55864 5692
rect 31938 5624 31944 5636
rect 29840 5596 31944 5624
rect 29733 5587 29791 5593
rect 26510 5556 26516 5568
rect 23584 5528 26516 5556
rect 23385 5519 23443 5525
rect 26510 5516 26516 5528
rect 26568 5516 26574 5568
rect 27614 5516 27620 5568
rect 27672 5556 27678 5568
rect 29748 5556 29776 5587
rect 31938 5584 31944 5596
rect 31996 5584 32002 5636
rect 33597 5627 33655 5633
rect 33597 5593 33609 5627
rect 33643 5624 33655 5627
rect 34054 5624 34060 5636
rect 33643 5596 34060 5624
rect 33643 5593 33655 5596
rect 33597 5587 33655 5593
rect 34054 5584 34060 5596
rect 34112 5584 34118 5636
rect 35161 5627 35219 5633
rect 35161 5593 35173 5627
rect 35207 5624 35219 5627
rect 38010 5624 38016 5636
rect 35207 5596 38016 5624
rect 35207 5593 35219 5596
rect 35161 5587 35219 5593
rect 38010 5584 38016 5596
rect 38068 5584 38074 5636
rect 38838 5584 38844 5636
rect 38896 5624 38902 5636
rect 39224 5633 39252 5664
rect 55858 5652 55864 5664
rect 55916 5652 55922 5704
rect 56980 5701 57008 5732
rect 57974 5720 57980 5732
rect 58032 5720 58038 5772
rect 58158 5760 58164 5772
rect 58119 5732 58164 5760
rect 58158 5720 58164 5732
rect 58216 5720 58222 5772
rect 56965 5695 57023 5701
rect 56965 5661 56977 5695
rect 57011 5661 57023 5695
rect 56965 5655 57023 5661
rect 57790 5652 57796 5704
rect 57848 5692 57854 5704
rect 57885 5695 57943 5701
rect 57885 5692 57897 5695
rect 57848 5664 57897 5692
rect 57848 5652 57854 5664
rect 57885 5661 57897 5664
rect 57931 5661 57943 5695
rect 57885 5655 57943 5661
rect 39117 5627 39175 5633
rect 39117 5624 39129 5627
rect 38896 5596 39129 5624
rect 38896 5584 38902 5596
rect 39117 5593 39129 5596
rect 39163 5593 39175 5627
rect 39117 5587 39175 5593
rect 39209 5627 39267 5633
rect 39209 5593 39221 5627
rect 39255 5593 39267 5627
rect 39209 5587 39267 5593
rect 27672 5528 29776 5556
rect 27672 5516 27678 5528
rect 31570 5516 31576 5568
rect 31628 5556 31634 5568
rect 31846 5556 31852 5568
rect 31628 5528 31852 5556
rect 31628 5516 31634 5528
rect 31846 5516 31852 5528
rect 31904 5556 31910 5568
rect 32585 5559 32643 5565
rect 32585 5556 32597 5559
rect 31904 5528 32597 5556
rect 31904 5516 31910 5528
rect 32585 5525 32597 5528
rect 32631 5525 32643 5559
rect 34238 5556 34244 5568
rect 34199 5528 34244 5556
rect 32585 5519 32643 5525
rect 34238 5516 34244 5528
rect 34296 5516 34302 5568
rect 36354 5556 36360 5568
rect 36315 5528 36360 5556
rect 36354 5516 36360 5528
rect 36412 5516 36418 5568
rect 37550 5516 37556 5568
rect 37608 5556 37614 5568
rect 37829 5559 37887 5565
rect 37829 5556 37841 5559
rect 37608 5528 37841 5556
rect 37608 5516 37614 5528
rect 37829 5525 37841 5528
rect 37875 5525 37887 5559
rect 37829 5519 37887 5525
rect 38749 5559 38807 5565
rect 38749 5525 38761 5559
rect 38795 5556 38807 5559
rect 38930 5556 38936 5568
rect 38795 5528 38936 5556
rect 38795 5525 38807 5528
rect 38749 5519 38807 5525
rect 38930 5516 38936 5528
rect 38988 5516 38994 5568
rect 39132 5556 39160 5587
rect 40034 5584 40040 5636
rect 40092 5624 40098 5636
rect 40129 5627 40187 5633
rect 40129 5624 40141 5627
rect 40092 5596 40141 5624
rect 40092 5584 40098 5596
rect 40129 5593 40141 5596
rect 40175 5593 40187 5627
rect 40129 5587 40187 5593
rect 41414 5584 41420 5636
rect 41472 5624 41478 5636
rect 57238 5624 57244 5636
rect 41472 5596 41517 5624
rect 57199 5596 57244 5624
rect 41472 5584 41478 5596
rect 57238 5584 57244 5596
rect 57296 5584 57302 5636
rect 39942 5556 39948 5568
rect 39132 5528 39948 5556
rect 39942 5516 39948 5528
rect 40000 5516 40006 5568
rect 1104 5466 58880 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 58880 5466
rect 1104 5392 58880 5414
rect 9401 5355 9459 5361
rect 9401 5321 9413 5355
rect 9447 5352 9459 5355
rect 9582 5352 9588 5364
rect 9447 5324 9588 5352
rect 9447 5321 9459 5324
rect 9401 5315 9459 5321
rect 9582 5312 9588 5324
rect 9640 5312 9646 5364
rect 10134 5352 10140 5364
rect 10095 5324 10140 5352
rect 10134 5312 10140 5324
rect 10192 5312 10198 5364
rect 14185 5355 14243 5361
rect 14185 5352 14197 5355
rect 12912 5324 14197 5352
rect 8938 5284 8944 5296
rect 8899 5256 8944 5284
rect 8938 5244 8944 5256
rect 8996 5244 9002 5296
rect 12912 5293 12940 5324
rect 14185 5321 14197 5324
rect 14231 5352 14243 5355
rect 14274 5352 14280 5364
rect 14231 5324 14280 5352
rect 14231 5321 14243 5324
rect 14185 5315 14243 5321
rect 14274 5312 14280 5324
rect 14332 5312 14338 5364
rect 18598 5352 18604 5364
rect 14660 5324 18604 5352
rect 12897 5287 12955 5293
rect 12897 5253 12909 5287
rect 12943 5253 12955 5287
rect 14660 5284 14688 5324
rect 18598 5312 18604 5324
rect 18656 5312 18662 5364
rect 19245 5355 19303 5361
rect 19245 5321 19257 5355
rect 19291 5352 19303 5355
rect 19334 5352 19340 5364
rect 19291 5324 19340 5352
rect 19291 5321 19303 5324
rect 19245 5315 19303 5321
rect 19334 5312 19340 5324
rect 19392 5312 19398 5364
rect 19705 5355 19763 5361
rect 19705 5321 19717 5355
rect 19751 5352 19763 5355
rect 20625 5355 20683 5361
rect 20625 5352 20637 5355
rect 19751 5324 20637 5352
rect 19751 5321 19763 5324
rect 19705 5315 19763 5321
rect 20625 5321 20637 5324
rect 20671 5321 20683 5355
rect 20625 5315 20683 5321
rect 25869 5355 25927 5361
rect 25869 5321 25881 5355
rect 25915 5352 25927 5355
rect 26050 5352 26056 5364
rect 25915 5324 26056 5352
rect 25915 5321 25927 5324
rect 25869 5315 25927 5321
rect 26050 5312 26056 5324
rect 26108 5312 26114 5364
rect 31110 5352 31116 5364
rect 26344 5324 30972 5352
rect 31071 5324 31116 5352
rect 12897 5247 12955 5253
rect 13648 5256 14688 5284
rect 1578 5216 1584 5228
rect 1539 5188 1584 5216
rect 1578 5176 1584 5188
rect 1636 5176 1642 5228
rect 8110 5176 8116 5228
rect 8168 5216 8174 5228
rect 8297 5219 8355 5225
rect 8297 5216 8309 5219
rect 8168 5188 8309 5216
rect 8168 5176 8174 5188
rect 8297 5185 8309 5188
rect 8343 5185 8355 5219
rect 8956 5216 8984 5244
rect 9582 5216 9588 5228
rect 8956 5188 9588 5216
rect 8297 5179 8355 5185
rect 9582 5176 9588 5188
rect 9640 5176 9646 5228
rect 10042 5176 10048 5228
rect 10100 5216 10106 5228
rect 10321 5219 10379 5225
rect 10321 5216 10333 5219
rect 10100 5188 10333 5216
rect 10100 5176 10106 5188
rect 10321 5185 10333 5188
rect 10367 5185 10379 5219
rect 10502 5216 10508 5228
rect 10463 5188 10508 5216
rect 10321 5179 10379 5185
rect 10502 5176 10508 5188
rect 10560 5176 10566 5228
rect 11974 5176 11980 5228
rect 12032 5216 12038 5228
rect 12161 5219 12219 5225
rect 12161 5216 12173 5219
rect 12032 5188 12173 5216
rect 12032 5176 12038 5188
rect 12161 5185 12173 5188
rect 12207 5185 12219 5219
rect 13648 5216 13676 5256
rect 14734 5244 14740 5296
rect 14792 5284 14798 5296
rect 20898 5284 20904 5296
rect 14792 5256 20904 5284
rect 14792 5244 14798 5256
rect 20898 5244 20904 5256
rect 20956 5244 20962 5296
rect 21085 5287 21143 5293
rect 21085 5253 21097 5287
rect 21131 5284 21143 5287
rect 26344 5284 26372 5324
rect 21131 5256 26372 5284
rect 21131 5253 21143 5256
rect 21085 5247 21143 5253
rect 26418 5244 26424 5296
rect 26476 5284 26482 5296
rect 27982 5284 27988 5296
rect 26476 5256 27988 5284
rect 26476 5244 26482 5256
rect 27982 5244 27988 5256
rect 28040 5244 28046 5296
rect 28442 5284 28448 5296
rect 28403 5256 28448 5284
rect 28442 5244 28448 5256
rect 28500 5284 28506 5296
rect 30834 5284 30840 5296
rect 28500 5256 30696 5284
rect 30795 5256 30840 5284
rect 28500 5244 28506 5256
rect 12161 5179 12219 5185
rect 12268 5188 13676 5216
rect 1762 5148 1768 5160
rect 1723 5120 1768 5148
rect 1762 5108 1768 5120
rect 1820 5108 1826 5160
rect 10413 5151 10471 5157
rect 10413 5117 10425 5151
rect 10459 5117 10471 5151
rect 10413 5111 10471 5117
rect 8481 5083 8539 5089
rect 8481 5049 8493 5083
rect 8527 5080 8539 5083
rect 8754 5080 8760 5092
rect 8527 5052 8760 5080
rect 8527 5049 8539 5052
rect 8481 5043 8539 5049
rect 8754 5040 8760 5052
rect 8812 5040 8818 5092
rect 9217 5083 9275 5089
rect 9217 5049 9229 5083
rect 9263 5049 9275 5083
rect 10428 5080 10456 5111
rect 10594 5108 10600 5160
rect 10652 5148 10658 5160
rect 10652 5120 10697 5148
rect 10652 5108 10658 5120
rect 12268 5080 12296 5188
rect 13722 5176 13728 5228
rect 13780 5216 13786 5228
rect 14001 5219 14059 5225
rect 14001 5216 14013 5219
rect 13780 5188 14013 5216
rect 13780 5176 13786 5188
rect 14001 5185 14013 5188
rect 14047 5185 14059 5219
rect 14001 5179 14059 5185
rect 17037 5219 17095 5225
rect 17037 5185 17049 5219
rect 17083 5185 17095 5219
rect 17037 5179 17095 5185
rect 17313 5219 17371 5225
rect 17313 5185 17325 5219
rect 17359 5216 17371 5219
rect 17402 5216 17408 5228
rect 17359 5188 17408 5216
rect 17359 5185 17371 5188
rect 17313 5179 17371 5185
rect 13357 5151 13415 5157
rect 13357 5117 13369 5151
rect 13403 5148 13415 5151
rect 13814 5148 13820 5160
rect 13403 5120 13820 5148
rect 13403 5117 13415 5120
rect 13357 5111 13415 5117
rect 13814 5108 13820 5120
rect 13872 5108 13878 5160
rect 10428 5052 12296 5080
rect 12345 5083 12403 5089
rect 9217 5043 9275 5049
rect 12345 5049 12357 5083
rect 12391 5080 12403 5083
rect 13173 5083 13231 5089
rect 13173 5080 13185 5083
rect 12391 5052 13185 5080
rect 12391 5049 12403 5052
rect 12345 5043 12403 5049
rect 13173 5049 13185 5052
rect 13219 5049 13231 5083
rect 17052 5080 17080 5179
rect 17402 5176 17408 5188
rect 17460 5176 17466 5228
rect 18046 5216 18052 5228
rect 18007 5188 18052 5216
rect 18046 5176 18052 5188
rect 18104 5176 18110 5228
rect 19334 5176 19340 5228
rect 19392 5216 19398 5228
rect 19613 5219 19671 5225
rect 19613 5216 19625 5219
rect 19392 5188 19625 5216
rect 19392 5176 19398 5188
rect 19613 5185 19625 5188
rect 19659 5216 19671 5219
rect 20254 5216 20260 5228
rect 19659 5188 20260 5216
rect 19659 5185 19671 5188
rect 19613 5179 19671 5185
rect 20254 5176 20260 5188
rect 20312 5176 20318 5228
rect 20622 5176 20628 5228
rect 20680 5216 20686 5228
rect 20993 5219 21051 5225
rect 20993 5216 21005 5219
rect 20680 5188 21005 5216
rect 20680 5176 20686 5188
rect 20993 5185 21005 5188
rect 21039 5185 21051 5219
rect 20993 5179 21051 5185
rect 22557 5219 22615 5225
rect 22557 5185 22569 5219
rect 22603 5216 22615 5219
rect 23382 5216 23388 5228
rect 22603 5188 23388 5216
rect 22603 5185 22615 5188
rect 22557 5179 22615 5185
rect 23382 5176 23388 5188
rect 23440 5176 23446 5228
rect 24946 5216 24952 5228
rect 23952 5188 24952 5216
rect 17126 5108 17132 5160
rect 17184 5148 17190 5160
rect 18325 5151 18383 5157
rect 18325 5148 18337 5151
rect 17184 5120 18337 5148
rect 17184 5108 17190 5120
rect 18325 5117 18337 5120
rect 18371 5117 18383 5151
rect 19886 5148 19892 5160
rect 19847 5120 19892 5148
rect 18325 5111 18383 5117
rect 19886 5108 19892 5120
rect 19944 5108 19950 5160
rect 21269 5151 21327 5157
rect 21269 5117 21281 5151
rect 21315 5148 21327 5151
rect 21358 5148 21364 5160
rect 21315 5120 21364 5148
rect 21315 5117 21327 5120
rect 21269 5111 21327 5117
rect 21358 5108 21364 5120
rect 21416 5108 21422 5160
rect 22462 5108 22468 5160
rect 22520 5148 22526 5160
rect 22741 5151 22799 5157
rect 22741 5148 22753 5151
rect 22520 5120 22753 5148
rect 22520 5108 22526 5120
rect 22741 5117 22753 5120
rect 22787 5117 22799 5151
rect 22741 5111 22799 5117
rect 23952 5080 23980 5188
rect 24946 5176 24952 5188
rect 25004 5176 25010 5228
rect 25130 5216 25136 5228
rect 25091 5188 25136 5216
rect 25130 5176 25136 5188
rect 25188 5176 25194 5228
rect 26237 5219 26295 5225
rect 26237 5216 26249 5219
rect 25240 5188 26249 5216
rect 24210 5108 24216 5160
rect 24268 5148 24274 5160
rect 25240 5148 25268 5188
rect 26237 5185 26249 5188
rect 26283 5185 26295 5219
rect 27154 5216 27160 5228
rect 27115 5188 27160 5216
rect 26237 5179 26295 5185
rect 27154 5176 27160 5188
rect 27212 5176 27218 5228
rect 27246 5176 27252 5228
rect 27304 5216 27310 5228
rect 28534 5216 28540 5228
rect 27304 5188 27349 5216
rect 28495 5188 28540 5216
rect 27304 5176 27310 5188
rect 28534 5176 28540 5188
rect 28592 5176 28598 5228
rect 29730 5216 29736 5228
rect 28644 5188 28994 5216
rect 29691 5188 29736 5216
rect 26326 5148 26332 5160
rect 24268 5120 25268 5148
rect 26287 5120 26332 5148
rect 24268 5108 24274 5120
rect 26326 5108 26332 5120
rect 26384 5108 26390 5160
rect 26510 5148 26516 5160
rect 26471 5120 26516 5148
rect 26510 5108 26516 5120
rect 26568 5148 26574 5160
rect 26878 5148 26884 5160
rect 26568 5120 26884 5148
rect 26568 5108 26574 5120
rect 26878 5108 26884 5120
rect 26936 5108 26942 5160
rect 28074 5108 28080 5160
rect 28132 5148 28138 5160
rect 28644 5148 28672 5188
rect 28132 5120 28672 5148
rect 28721 5151 28779 5157
rect 28132 5108 28138 5120
rect 28721 5117 28733 5151
rect 28767 5117 28779 5151
rect 28966 5148 28994 5188
rect 29730 5176 29736 5188
rect 29788 5176 29794 5228
rect 29917 5219 29975 5225
rect 29917 5185 29929 5219
rect 29963 5185 29975 5219
rect 29917 5179 29975 5185
rect 30009 5219 30067 5225
rect 30009 5185 30021 5219
rect 30055 5185 30067 5219
rect 30009 5179 30067 5185
rect 30153 5219 30211 5225
rect 30153 5185 30165 5219
rect 30199 5216 30211 5219
rect 30558 5216 30564 5228
rect 30199 5188 30564 5216
rect 30199 5185 30211 5188
rect 30153 5179 30211 5185
rect 29932 5148 29960 5179
rect 28966 5120 29960 5148
rect 30024 5148 30052 5179
rect 30558 5176 30564 5188
rect 30616 5176 30622 5228
rect 30668 5216 30696 5256
rect 30834 5244 30840 5256
rect 30892 5244 30898 5296
rect 30944 5284 30972 5324
rect 31110 5312 31116 5324
rect 31168 5312 31174 5364
rect 31205 5355 31263 5361
rect 31205 5321 31217 5355
rect 31251 5352 31263 5355
rect 31386 5352 31392 5364
rect 31251 5324 31392 5352
rect 31251 5321 31263 5324
rect 31205 5315 31263 5321
rect 31386 5312 31392 5324
rect 31444 5312 31450 5364
rect 35618 5312 35624 5364
rect 35676 5352 35682 5364
rect 35676 5324 40632 5352
rect 35676 5312 35682 5324
rect 32582 5284 32588 5296
rect 30944 5256 32588 5284
rect 32582 5244 32588 5256
rect 32640 5244 32646 5296
rect 32861 5287 32919 5293
rect 32861 5253 32873 5287
rect 32907 5284 32919 5287
rect 33597 5287 33655 5293
rect 33597 5284 33609 5287
rect 32907 5256 33609 5284
rect 32907 5253 32919 5256
rect 32861 5247 32919 5253
rect 33597 5253 33609 5256
rect 33643 5284 33655 5287
rect 33778 5284 33784 5296
rect 33643 5256 33784 5284
rect 33643 5253 33655 5256
rect 33597 5247 33655 5253
rect 33778 5244 33784 5256
rect 33836 5284 33842 5296
rect 34333 5287 34391 5293
rect 34333 5284 34345 5287
rect 33836 5256 34345 5284
rect 33836 5244 33842 5256
rect 34333 5253 34345 5256
rect 34379 5253 34391 5287
rect 34333 5247 34391 5253
rect 34790 5244 34796 5296
rect 34848 5284 34854 5296
rect 34848 5256 36400 5284
rect 34848 5244 34854 5256
rect 30668 5188 30972 5216
rect 30944 5148 30972 5188
rect 31018 5176 31024 5228
rect 31076 5216 31082 5228
rect 31076 5188 31121 5216
rect 31076 5176 31082 5188
rect 31294 5176 31300 5228
rect 31352 5216 31358 5228
rect 31389 5219 31447 5225
rect 31389 5216 31401 5219
rect 31352 5188 31401 5216
rect 31352 5176 31358 5188
rect 31389 5185 31401 5188
rect 31435 5185 31447 5219
rect 31389 5179 31447 5185
rect 34977 5219 35035 5225
rect 34977 5185 34989 5219
rect 35023 5216 35035 5219
rect 35342 5216 35348 5228
rect 35023 5188 35348 5216
rect 35023 5185 35035 5188
rect 34977 5179 35035 5185
rect 35342 5176 35348 5188
rect 35400 5176 35406 5228
rect 35894 5216 35900 5228
rect 35855 5188 35900 5216
rect 35894 5176 35900 5188
rect 35952 5176 35958 5228
rect 36372 5216 36400 5256
rect 36446 5244 36452 5296
rect 36504 5284 36510 5296
rect 40218 5284 40224 5296
rect 36504 5256 40224 5284
rect 36504 5244 36510 5256
rect 40218 5244 40224 5256
rect 40276 5244 40282 5296
rect 40604 5284 40632 5324
rect 40678 5312 40684 5364
rect 40736 5352 40742 5364
rect 41969 5355 42027 5361
rect 41969 5352 41981 5355
rect 40736 5324 41981 5352
rect 40736 5312 40742 5324
rect 41969 5321 41981 5324
rect 42015 5321 42027 5355
rect 42794 5352 42800 5364
rect 42755 5324 42800 5352
rect 41969 5315 42027 5321
rect 42794 5312 42800 5324
rect 42852 5312 42858 5364
rect 43162 5312 43168 5364
rect 43220 5352 43226 5364
rect 43533 5355 43591 5361
rect 43533 5352 43545 5355
rect 43220 5324 43545 5352
rect 43220 5312 43226 5324
rect 43533 5321 43545 5324
rect 43579 5321 43591 5355
rect 58253 5355 58311 5361
rect 58253 5352 58265 5355
rect 43533 5315 43591 5321
rect 55186 5324 58265 5352
rect 55186 5284 55214 5324
rect 58253 5321 58265 5324
rect 58299 5321 58311 5355
rect 58253 5315 58311 5321
rect 40604 5256 55214 5284
rect 37182 5216 37188 5228
rect 36372 5188 37188 5216
rect 37182 5176 37188 5188
rect 37240 5176 37246 5228
rect 37366 5176 37372 5228
rect 37424 5216 37430 5228
rect 37461 5219 37519 5225
rect 37461 5216 37473 5219
rect 37424 5188 37473 5216
rect 37424 5176 37430 5188
rect 37461 5185 37473 5188
rect 37507 5185 37519 5219
rect 37642 5216 37648 5228
rect 37603 5188 37648 5216
rect 37461 5179 37519 5185
rect 33226 5148 33232 5160
rect 30024 5120 30788 5148
rect 30944 5120 33232 5148
rect 28721 5111 28779 5117
rect 13173 5043 13231 5049
rect 13280 5052 16804 5080
rect 17052 5052 23980 5080
rect 24029 5083 24087 5089
rect 7098 4972 7104 5024
rect 7156 5012 7162 5024
rect 9232 5012 9260 5043
rect 7156 4984 9260 5012
rect 7156 4972 7162 4984
rect 9674 4972 9680 5024
rect 9732 5012 9738 5024
rect 13280 5012 13308 5052
rect 9732 4984 13308 5012
rect 16301 5015 16359 5021
rect 9732 4972 9738 4984
rect 16301 4981 16313 5015
rect 16347 5012 16359 5015
rect 16666 5012 16672 5024
rect 16347 4984 16672 5012
rect 16347 4981 16359 4984
rect 16301 4975 16359 4981
rect 16666 4972 16672 4984
rect 16724 4972 16730 5024
rect 16776 5012 16804 5052
rect 24029 5049 24041 5083
rect 24075 5080 24087 5083
rect 24075 5052 25728 5080
rect 24075 5049 24087 5052
rect 24029 5043 24087 5049
rect 20257 5015 20315 5021
rect 20257 5012 20269 5015
rect 16776 4984 20269 5012
rect 20257 4981 20269 4984
rect 20303 5012 20315 5015
rect 20622 5012 20628 5024
rect 20303 4984 20628 5012
rect 20303 4981 20315 4984
rect 20257 4975 20315 4981
rect 20622 4972 20628 4984
rect 20680 4972 20686 5024
rect 24670 5012 24676 5024
rect 24631 4984 24676 5012
rect 24670 4972 24676 4984
rect 24728 4972 24734 5024
rect 24946 4972 24952 5024
rect 25004 5012 25010 5024
rect 25317 5015 25375 5021
rect 25317 5012 25329 5015
rect 25004 4984 25329 5012
rect 25004 4972 25010 4984
rect 25317 4981 25329 4984
rect 25363 4981 25375 5015
rect 25700 5012 25728 5052
rect 28626 5040 28632 5092
rect 28684 5080 28690 5092
rect 28736 5080 28764 5111
rect 28684 5052 28764 5080
rect 28684 5040 28690 5052
rect 28810 5040 28816 5092
rect 28868 5080 28874 5092
rect 30190 5080 30196 5092
rect 28868 5052 30196 5080
rect 28868 5040 28874 5052
rect 30190 5040 30196 5052
rect 30248 5040 30254 5092
rect 25774 5012 25780 5024
rect 25700 4984 25780 5012
rect 25317 4975 25375 4981
rect 25774 4972 25780 4984
rect 25832 4972 25838 5024
rect 25866 4972 25872 5024
rect 25924 5012 25930 5024
rect 27157 5015 27215 5021
rect 27157 5012 27169 5015
rect 25924 4984 27169 5012
rect 25924 4972 25930 4984
rect 27157 4981 27169 4984
rect 27203 4981 27215 5015
rect 27522 5012 27528 5024
rect 27483 4984 27528 5012
rect 27157 4975 27215 4981
rect 27522 4972 27528 4984
rect 27580 4972 27586 5024
rect 28074 5012 28080 5024
rect 28035 4984 28080 5012
rect 28074 4972 28080 4984
rect 28132 4972 28138 5024
rect 30006 4972 30012 5024
rect 30064 5012 30070 5024
rect 30285 5015 30343 5021
rect 30285 5012 30297 5015
rect 30064 4984 30297 5012
rect 30064 4972 30070 4984
rect 30285 4981 30297 4984
rect 30331 4981 30343 5015
rect 30760 5012 30788 5120
rect 33226 5108 33232 5120
rect 33284 5108 33290 5160
rect 34790 5108 34796 5160
rect 34848 5148 34854 5160
rect 35161 5151 35219 5157
rect 35161 5148 35173 5151
rect 34848 5120 35173 5148
rect 34848 5108 34854 5120
rect 35161 5117 35173 5120
rect 35207 5117 35219 5151
rect 35161 5111 35219 5117
rect 35434 5108 35440 5160
rect 35492 5148 35498 5160
rect 36081 5151 36139 5157
rect 36081 5148 36093 5151
rect 35492 5120 36093 5148
rect 35492 5108 35498 5120
rect 36081 5117 36093 5120
rect 36127 5117 36139 5151
rect 37476 5148 37504 5179
rect 37642 5176 37648 5188
rect 37700 5176 37706 5228
rect 38930 5216 38936 5228
rect 38891 5188 38936 5216
rect 38930 5176 38936 5188
rect 38988 5176 38994 5228
rect 39666 5216 39672 5228
rect 39627 5188 39672 5216
rect 39666 5176 39672 5188
rect 39724 5176 39730 5228
rect 40313 5219 40371 5225
rect 40313 5216 40325 5219
rect 39776 5188 40325 5216
rect 38749 5151 38807 5157
rect 38749 5148 38761 5151
rect 37476 5120 38761 5148
rect 36081 5111 36139 5117
rect 38749 5117 38761 5120
rect 38795 5117 38807 5151
rect 38749 5111 38807 5117
rect 33042 5080 33048 5092
rect 33003 5052 33048 5080
rect 33042 5040 33048 5052
rect 33100 5040 33106 5092
rect 33781 5083 33839 5089
rect 33781 5049 33793 5083
rect 33827 5080 33839 5083
rect 33827 5052 34652 5080
rect 33827 5049 33839 5052
rect 33781 5043 33839 5049
rect 34146 5012 34152 5024
rect 30760 4984 34152 5012
rect 30285 4975 30343 4981
rect 34146 4972 34152 4984
rect 34204 4972 34210 5024
rect 34422 5012 34428 5024
rect 34383 4984 34428 5012
rect 34422 4972 34428 4984
rect 34480 4972 34486 5024
rect 34624 5012 34652 5052
rect 38470 5040 38476 5092
rect 38528 5080 38534 5092
rect 39776 5080 39804 5188
rect 40313 5185 40325 5188
rect 40359 5185 40371 5219
rect 40313 5179 40371 5185
rect 40494 5176 40500 5228
rect 40552 5216 40558 5228
rect 41141 5219 41199 5225
rect 41141 5216 41153 5219
rect 40552 5188 41153 5216
rect 40552 5176 40558 5188
rect 41141 5185 41153 5188
rect 41187 5185 41199 5219
rect 41141 5179 41199 5185
rect 41598 5176 41604 5228
rect 41656 5216 41662 5228
rect 41785 5219 41843 5225
rect 41785 5216 41797 5219
rect 41656 5188 41797 5216
rect 41656 5176 41662 5188
rect 41785 5185 41797 5188
rect 41831 5185 41843 5219
rect 41785 5179 41843 5185
rect 41874 5176 41880 5228
rect 41932 5216 41938 5228
rect 42705 5219 42763 5225
rect 42705 5216 42717 5219
rect 41932 5188 42717 5216
rect 41932 5176 41938 5188
rect 42705 5185 42717 5188
rect 42751 5185 42763 5219
rect 42705 5179 42763 5185
rect 42886 5176 42892 5228
rect 42944 5216 42950 5228
rect 43441 5219 43499 5225
rect 43441 5216 43453 5219
rect 42944 5188 43453 5216
rect 42944 5176 42950 5188
rect 43441 5185 43453 5188
rect 43487 5185 43499 5219
rect 44174 5216 44180 5228
rect 44135 5188 44180 5216
rect 43441 5179 43499 5185
rect 44174 5176 44180 5188
rect 44232 5176 44238 5228
rect 44542 5176 44548 5228
rect 44600 5216 44606 5228
rect 44913 5219 44971 5225
rect 44913 5216 44925 5219
rect 44600 5188 44925 5216
rect 44600 5176 44606 5188
rect 44913 5185 44925 5188
rect 44959 5185 44971 5219
rect 44913 5179 44971 5185
rect 45646 5176 45652 5228
rect 45704 5216 45710 5228
rect 45833 5219 45891 5225
rect 45833 5216 45845 5219
rect 45704 5188 45845 5216
rect 45704 5176 45710 5188
rect 45833 5185 45845 5188
rect 45879 5185 45891 5219
rect 48774 5216 48780 5228
rect 48735 5188 48780 5216
rect 45833 5179 45891 5185
rect 48774 5176 48780 5188
rect 48832 5176 48838 5228
rect 49033 5219 49091 5225
rect 49033 5216 49045 5219
rect 48884 5188 49045 5216
rect 46017 5151 46075 5157
rect 46017 5148 46029 5151
rect 40512 5120 46029 5148
rect 38528 5052 39804 5080
rect 38528 5040 38534 5052
rect 40218 5040 40224 5092
rect 40276 5080 40282 5092
rect 40512 5080 40540 5120
rect 46017 5117 46029 5120
rect 46063 5117 46075 5151
rect 46017 5111 46075 5117
rect 46750 5108 46756 5160
rect 46808 5148 46814 5160
rect 48884 5148 48912 5188
rect 49033 5185 49045 5188
rect 49079 5185 49091 5219
rect 58066 5216 58072 5228
rect 58027 5188 58072 5216
rect 49033 5179 49091 5185
rect 58066 5176 58072 5188
rect 58124 5176 58130 5228
rect 46808 5120 48912 5148
rect 46808 5108 46814 5120
rect 40276 5052 40540 5080
rect 44361 5083 44419 5089
rect 40276 5040 40282 5052
rect 44361 5049 44373 5083
rect 44407 5080 44419 5083
rect 44450 5080 44456 5092
rect 44407 5052 44456 5080
rect 44407 5049 44419 5052
rect 44361 5043 44419 5049
rect 44450 5040 44456 5052
rect 44508 5040 44514 5092
rect 44634 5040 44640 5092
rect 44692 5080 44698 5092
rect 45186 5080 45192 5092
rect 44692 5052 45192 5080
rect 44692 5040 44698 5052
rect 45186 5040 45192 5052
rect 45244 5040 45250 5092
rect 34698 5012 34704 5024
rect 34624 4984 34704 5012
rect 34698 4972 34704 4984
rect 34756 4972 34762 5024
rect 37826 5012 37832 5024
rect 37787 4984 37832 5012
rect 37826 4972 37832 4984
rect 37884 4972 37890 5024
rect 38838 4972 38844 5024
rect 38896 5012 38902 5024
rect 39117 5015 39175 5021
rect 39117 5012 39129 5015
rect 38896 4984 39129 5012
rect 38896 4972 38902 4984
rect 39117 4981 39129 4984
rect 39163 4981 39175 5015
rect 39117 4975 39175 4981
rect 39206 4972 39212 5024
rect 39264 5012 39270 5024
rect 39761 5015 39819 5021
rect 39761 5012 39773 5015
rect 39264 4984 39773 5012
rect 39264 4972 39270 4984
rect 39761 4981 39773 4984
rect 39807 4981 39819 5015
rect 39761 4975 39819 4981
rect 40497 5015 40555 5021
rect 40497 4981 40509 5015
rect 40543 5012 40555 5015
rect 40678 5012 40684 5024
rect 40543 4984 40684 5012
rect 40543 4981 40555 4984
rect 40497 4975 40555 4981
rect 40678 4972 40684 4984
rect 40736 4972 40742 5024
rect 41138 4972 41144 5024
rect 41196 5012 41202 5024
rect 41233 5015 41291 5021
rect 41233 5012 41245 5015
rect 41196 4984 41245 5012
rect 41196 4972 41202 4984
rect 41233 4981 41245 4984
rect 41279 4981 41291 5015
rect 41233 4975 41291 4981
rect 41690 4972 41696 5024
rect 41748 5012 41754 5024
rect 44266 5012 44272 5024
rect 41748 4984 44272 5012
rect 41748 4972 41754 4984
rect 44266 4972 44272 4984
rect 44324 4972 44330 5024
rect 45002 5012 45008 5024
rect 44963 4984 45008 5012
rect 45002 4972 45008 4984
rect 45060 4972 45066 5024
rect 50157 5015 50215 5021
rect 50157 4981 50169 5015
rect 50203 5012 50215 5015
rect 51442 5012 51448 5024
rect 50203 4984 51448 5012
rect 50203 4981 50215 4984
rect 50157 4975 50215 4981
rect 51442 4972 51448 4984
rect 51500 4972 51506 5024
rect 1104 4922 58880 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 58880 4922
rect 1104 4848 58880 4870
rect 9858 4808 9864 4820
rect 9646 4780 9864 4808
rect 1578 4700 1584 4752
rect 1636 4740 1642 4752
rect 8573 4743 8631 4749
rect 1636 4712 2774 4740
rect 1636 4700 1642 4712
rect 2746 4672 2774 4712
rect 8573 4709 8585 4743
rect 8619 4740 8631 4743
rect 9646 4740 9674 4780
rect 9858 4768 9864 4780
rect 9916 4768 9922 4820
rect 11057 4811 11115 4817
rect 11057 4777 11069 4811
rect 11103 4808 11115 4811
rect 11238 4808 11244 4820
rect 11103 4780 11244 4808
rect 11103 4777 11115 4780
rect 11057 4771 11115 4777
rect 11238 4768 11244 4780
rect 11296 4768 11302 4820
rect 13722 4768 13728 4820
rect 13780 4808 13786 4820
rect 15381 4811 15439 4817
rect 15381 4808 15393 4811
rect 13780 4780 15393 4808
rect 13780 4768 13786 4780
rect 15381 4777 15393 4780
rect 15427 4777 15439 4811
rect 15381 4771 15439 4777
rect 17494 4768 17500 4820
rect 17552 4808 17558 4820
rect 21821 4811 21879 4817
rect 21821 4808 21833 4811
rect 17552 4780 21833 4808
rect 17552 4768 17558 4780
rect 21821 4777 21833 4780
rect 21867 4777 21879 4811
rect 21821 4771 21879 4777
rect 24670 4768 24676 4820
rect 24728 4808 24734 4820
rect 25590 4808 25596 4820
rect 24728 4780 25596 4808
rect 24728 4768 24734 4780
rect 25590 4768 25596 4780
rect 25648 4768 25654 4820
rect 27525 4811 27583 4817
rect 27525 4808 27537 4811
rect 26252 4780 27537 4808
rect 8619 4712 9674 4740
rect 8619 4709 8631 4712
rect 8573 4703 8631 4709
rect 10042 4700 10048 4752
rect 10100 4740 10106 4752
rect 10873 4743 10931 4749
rect 10873 4740 10885 4743
rect 10100 4712 10885 4740
rect 10100 4700 10106 4712
rect 10873 4709 10885 4712
rect 10919 4709 10931 4743
rect 10873 4703 10931 4709
rect 12066 4700 12072 4752
rect 12124 4740 12130 4752
rect 13541 4743 13599 4749
rect 13541 4740 13553 4743
rect 12124 4712 13553 4740
rect 12124 4700 12130 4712
rect 13541 4709 13553 4712
rect 13587 4709 13599 4743
rect 14553 4743 14611 4749
rect 14553 4740 14565 4743
rect 13541 4703 13599 4709
rect 13648 4712 14565 4740
rect 9585 4675 9643 4681
rect 9585 4672 9597 4675
rect 2746 4644 9597 4672
rect 9585 4641 9597 4644
rect 9631 4641 9643 4675
rect 9585 4635 9643 4641
rect 9674 4632 9680 4684
rect 9732 4632 9738 4684
rect 9766 4632 9772 4684
rect 9824 4672 9830 4684
rect 9824 4644 9869 4672
rect 9824 4632 9830 4644
rect 9950 4632 9956 4684
rect 10008 4672 10014 4684
rect 10410 4672 10416 4684
rect 10008 4644 10416 4672
rect 10008 4632 10014 4644
rect 10410 4632 10416 4644
rect 10468 4672 10474 4684
rect 10597 4675 10655 4681
rect 10597 4672 10609 4675
rect 10468 4644 10609 4672
rect 10468 4632 10474 4644
rect 10597 4641 10609 4644
rect 10643 4641 10655 4675
rect 10597 4635 10655 4641
rect 12805 4675 12863 4681
rect 12805 4641 12817 4675
rect 12851 4672 12863 4675
rect 13648 4672 13676 4712
rect 14553 4709 14565 4712
rect 14599 4709 14611 4743
rect 14734 4740 14740 4752
rect 14695 4712 14740 4740
rect 14553 4703 14611 4709
rect 14734 4700 14740 4712
rect 14792 4700 14798 4752
rect 15194 4700 15200 4752
rect 15252 4740 15258 4752
rect 15654 4740 15660 4752
rect 15252 4712 15660 4740
rect 15252 4700 15258 4712
rect 15654 4700 15660 4712
rect 15712 4740 15718 4752
rect 17310 4740 17316 4752
rect 15712 4712 17316 4740
rect 15712 4700 15718 4712
rect 17310 4700 17316 4712
rect 17368 4700 17374 4752
rect 19886 4700 19892 4752
rect 19944 4740 19950 4752
rect 23750 4740 23756 4752
rect 19944 4712 23756 4740
rect 19944 4700 19950 4712
rect 23750 4700 23756 4712
rect 23808 4740 23814 4752
rect 23808 4712 23888 4740
rect 23808 4700 23814 4712
rect 12851 4644 13676 4672
rect 17773 4675 17831 4681
rect 12851 4641 12863 4644
rect 12805 4635 12863 4641
rect 17773 4641 17785 4675
rect 17819 4672 17831 4675
rect 18874 4672 18880 4684
rect 17819 4644 18880 4672
rect 17819 4641 17831 4644
rect 17773 4635 17831 4641
rect 18874 4632 18880 4644
rect 18932 4632 18938 4684
rect 18966 4632 18972 4684
rect 19024 4672 19030 4684
rect 20993 4675 21051 4681
rect 20993 4672 21005 4675
rect 19024 4644 21005 4672
rect 19024 4632 19030 4644
rect 20993 4641 21005 4644
rect 21039 4641 21051 4675
rect 21174 4672 21180 4684
rect 21135 4644 21180 4672
rect 20993 4635 21051 4641
rect 4614 4564 4620 4616
rect 4672 4604 4678 4616
rect 9692 4604 9720 4632
rect 4672 4576 9720 4604
rect 4672 4564 4678 4576
rect 9858 4564 9864 4616
rect 9916 4604 9922 4616
rect 10045 4607 10103 4613
rect 9916 4576 9961 4604
rect 9916 4564 9922 4576
rect 10045 4573 10057 4607
rect 10091 4604 10103 4607
rect 12069 4607 12127 4613
rect 10091 4576 10180 4604
rect 10091 4573 10103 4576
rect 10045 4567 10103 4573
rect 6914 4536 6920 4548
rect 6875 4508 6920 4536
rect 6914 4496 6920 4508
rect 6972 4496 6978 4548
rect 7653 4539 7711 4545
rect 7653 4505 7665 4539
rect 7699 4536 7711 4539
rect 8294 4536 8300 4548
rect 7699 4508 8300 4536
rect 7699 4505 7711 4508
rect 7653 4499 7711 4505
rect 8294 4496 8300 4508
rect 8352 4496 8358 4548
rect 8389 4539 8447 4545
rect 8389 4505 8401 4539
rect 8435 4505 8447 4539
rect 8389 4499 8447 4505
rect 7006 4468 7012 4480
rect 6967 4440 7012 4468
rect 7006 4428 7012 4440
rect 7064 4428 7070 4480
rect 7558 4428 7564 4480
rect 7616 4468 7622 4480
rect 7745 4471 7803 4477
rect 7745 4468 7757 4471
rect 7616 4440 7757 4468
rect 7616 4428 7622 4440
rect 7745 4437 7757 4440
rect 7791 4437 7803 4471
rect 8404 4468 8432 4499
rect 8846 4496 8852 4548
rect 8904 4536 8910 4548
rect 8904 4508 9904 4536
rect 8904 4496 8910 4508
rect 9766 4468 9772 4480
rect 8404 4440 9772 4468
rect 7745 4431 7803 4437
rect 9766 4428 9772 4440
rect 9824 4428 9830 4480
rect 9876 4468 9904 4508
rect 10152 4468 10180 4576
rect 12069 4573 12081 4607
rect 12115 4604 12127 4607
rect 12986 4604 12992 4616
rect 12115 4576 12992 4604
rect 12115 4573 12127 4576
rect 12069 4567 12127 4573
rect 12986 4564 12992 4576
rect 13044 4564 13050 4616
rect 13265 4607 13323 4613
rect 13265 4573 13277 4607
rect 13311 4604 13323 4607
rect 14274 4604 14280 4616
rect 13311 4576 14280 4604
rect 13311 4573 13323 4576
rect 13265 4567 13323 4573
rect 14274 4564 14280 4576
rect 14332 4564 14338 4616
rect 14734 4564 14740 4616
rect 14792 4604 14798 4616
rect 15289 4607 15347 4613
rect 15289 4604 15301 4607
rect 14792 4576 15301 4604
rect 14792 4564 14798 4576
rect 15289 4573 15301 4576
rect 15335 4573 15347 4607
rect 15289 4567 15347 4573
rect 16117 4607 16175 4613
rect 16117 4573 16129 4607
rect 16163 4604 16175 4607
rect 16390 4604 16396 4616
rect 16163 4576 16396 4604
rect 16163 4573 16175 4576
rect 16117 4567 16175 4573
rect 16390 4564 16396 4576
rect 16448 4564 16454 4616
rect 16574 4604 16580 4616
rect 16535 4576 16580 4604
rect 16574 4564 16580 4576
rect 16632 4564 16638 4616
rect 17497 4607 17555 4613
rect 17497 4573 17509 4607
rect 17543 4604 17555 4607
rect 17862 4604 17868 4616
rect 17543 4576 17868 4604
rect 17543 4573 17555 4576
rect 17497 4567 17555 4573
rect 17862 4564 17868 4576
rect 17920 4564 17926 4616
rect 18322 4564 18328 4616
rect 18380 4604 18386 4616
rect 18417 4607 18475 4613
rect 18417 4604 18429 4607
rect 18380 4576 18429 4604
rect 18380 4564 18386 4576
rect 18417 4573 18429 4576
rect 18463 4573 18475 4607
rect 19426 4604 19432 4616
rect 18417 4567 18475 4573
rect 19306 4576 19432 4604
rect 11790 4496 11796 4548
rect 11848 4536 11854 4548
rect 11885 4539 11943 4545
rect 11885 4536 11897 4539
rect 11848 4508 11897 4536
rect 11848 4496 11854 4508
rect 11885 4505 11897 4508
rect 11931 4505 11943 4539
rect 11885 4499 11943 4505
rect 12621 4539 12679 4545
rect 12621 4505 12633 4539
rect 12667 4536 12679 4539
rect 13078 4536 13084 4548
rect 12667 4508 13084 4536
rect 12667 4505 12679 4508
rect 12621 4499 12679 4505
rect 13078 4496 13084 4508
rect 13136 4496 13142 4548
rect 16853 4539 16911 4545
rect 16853 4505 16865 4539
rect 16899 4536 16911 4539
rect 18046 4536 18052 4548
rect 16899 4508 18052 4536
rect 16899 4505 16911 4508
rect 16853 4499 16911 4505
rect 18046 4496 18052 4508
rect 18104 4496 18110 4548
rect 18693 4539 18751 4545
rect 18693 4505 18705 4539
rect 18739 4536 18751 4539
rect 19306 4536 19334 4576
rect 19426 4564 19432 4576
rect 19484 4564 19490 4616
rect 19613 4607 19671 4613
rect 19613 4573 19625 4607
rect 19659 4604 19671 4607
rect 20070 4604 20076 4616
rect 19659 4576 20076 4604
rect 19659 4573 19671 4576
rect 19613 4567 19671 4573
rect 20070 4564 20076 4576
rect 20128 4564 20134 4616
rect 21008 4604 21036 4635
rect 21174 4632 21180 4644
rect 21232 4632 21238 4684
rect 23860 4681 23888 4712
rect 25222 4700 25228 4752
rect 25280 4740 25286 4752
rect 25866 4740 25872 4752
rect 25280 4712 25872 4740
rect 25280 4700 25286 4712
rect 25866 4700 25872 4712
rect 25924 4700 25930 4752
rect 25958 4700 25964 4752
rect 26016 4740 26022 4752
rect 26252 4740 26280 4780
rect 27525 4777 27537 4780
rect 27571 4777 27583 4811
rect 27706 4808 27712 4820
rect 27667 4780 27712 4808
rect 27525 4771 27583 4777
rect 27706 4768 27712 4780
rect 27764 4768 27770 4820
rect 30469 4811 30527 4817
rect 30469 4777 30481 4811
rect 30515 4808 30527 4811
rect 31754 4808 31760 4820
rect 30515 4780 31760 4808
rect 30515 4777 30527 4780
rect 30469 4771 30527 4777
rect 31754 4768 31760 4780
rect 31812 4768 31818 4820
rect 35342 4768 35348 4820
rect 35400 4808 35406 4820
rect 37645 4811 37703 4817
rect 37645 4808 37657 4811
rect 35400 4780 37657 4808
rect 35400 4768 35406 4780
rect 37645 4777 37657 4780
rect 37691 4777 37703 4811
rect 40770 4808 40776 4820
rect 37645 4771 37703 4777
rect 37752 4780 40776 4808
rect 26016 4712 26280 4740
rect 26016 4700 26022 4712
rect 26326 4700 26332 4752
rect 26384 4740 26390 4752
rect 31846 4740 31852 4752
rect 26384 4712 31852 4740
rect 26384 4700 26390 4712
rect 31846 4700 31852 4712
rect 31904 4700 31910 4752
rect 32125 4743 32183 4749
rect 32125 4709 32137 4743
rect 32171 4740 32183 4743
rect 32171 4712 33548 4740
rect 32171 4709 32183 4712
rect 32125 4703 32183 4709
rect 23845 4675 23903 4681
rect 23845 4641 23857 4675
rect 23891 4641 23903 4675
rect 23845 4635 23903 4641
rect 24946 4632 24952 4684
rect 25004 4672 25010 4684
rect 26697 4675 26755 4681
rect 25004 4644 26648 4672
rect 25004 4632 25010 4644
rect 21358 4604 21364 4616
rect 21008 4576 21364 4604
rect 21358 4564 21364 4576
rect 21416 4564 21422 4616
rect 21729 4607 21787 4613
rect 21729 4573 21741 4607
rect 21775 4604 21787 4607
rect 22002 4604 22008 4616
rect 21775 4576 22008 4604
rect 21775 4573 21787 4576
rect 21729 4567 21787 4573
rect 22002 4564 22008 4576
rect 22060 4564 22066 4616
rect 22370 4604 22376 4616
rect 22331 4576 22376 4604
rect 22370 4564 22376 4576
rect 22428 4564 22434 4616
rect 24486 4604 24492 4616
rect 22572 4576 24492 4604
rect 19886 4536 19892 4548
rect 18739 4508 19334 4536
rect 19847 4508 19892 4536
rect 18739 4505 18751 4508
rect 18693 4499 18751 4505
rect 19886 4496 19892 4508
rect 19944 4496 19950 4548
rect 20901 4539 20959 4545
rect 20364 4508 20668 4536
rect 9876 4440 10180 4468
rect 13725 4471 13783 4477
rect 13725 4437 13737 4471
rect 13771 4468 13783 4471
rect 17218 4468 17224 4480
rect 13771 4440 17224 4468
rect 13771 4437 13783 4440
rect 13725 4431 13783 4437
rect 17218 4428 17224 4440
rect 17276 4428 17282 4480
rect 17310 4428 17316 4480
rect 17368 4468 17374 4480
rect 20364 4468 20392 4508
rect 20530 4468 20536 4480
rect 17368 4440 20392 4468
rect 20491 4440 20536 4468
rect 17368 4428 17374 4440
rect 20530 4428 20536 4440
rect 20588 4428 20594 4480
rect 20640 4468 20668 4508
rect 20901 4505 20913 4539
rect 20947 4536 20959 4539
rect 22572 4536 22600 4576
rect 24486 4564 24492 4576
rect 24544 4564 24550 4616
rect 24670 4604 24676 4616
rect 24631 4576 24676 4604
rect 24670 4564 24676 4576
rect 24728 4564 24734 4616
rect 25406 4564 25412 4616
rect 25464 4604 25470 4616
rect 25958 4604 25964 4616
rect 25464 4576 25964 4604
rect 25464 4564 25470 4576
rect 25958 4564 25964 4576
rect 26016 4564 26022 4616
rect 26418 4604 26424 4616
rect 26379 4576 26424 4604
rect 26418 4564 26424 4576
rect 26476 4564 26482 4616
rect 26513 4607 26571 4613
rect 26513 4573 26525 4607
rect 26559 4573 26571 4607
rect 26620 4604 26648 4644
rect 26697 4641 26709 4675
rect 26743 4672 26755 4675
rect 28350 4672 28356 4684
rect 26743 4644 28356 4672
rect 26743 4641 26755 4644
rect 26697 4635 26755 4641
rect 28350 4632 28356 4644
rect 28408 4632 28414 4684
rect 31938 4672 31944 4684
rect 28552 4644 31944 4672
rect 28552 4613 28580 4644
rect 31938 4632 31944 4644
rect 31996 4632 32002 4684
rect 32030 4632 32036 4684
rect 32088 4672 32094 4684
rect 32677 4675 32735 4681
rect 32677 4672 32689 4675
rect 32088 4644 32689 4672
rect 32088 4632 32094 4644
rect 32677 4641 32689 4644
rect 32723 4672 32735 4675
rect 32858 4672 32864 4684
rect 32723 4644 32864 4672
rect 32723 4641 32735 4644
rect 32677 4635 32735 4641
rect 32858 4632 32864 4644
rect 32916 4632 32922 4684
rect 27157 4607 27215 4613
rect 27157 4604 27169 4607
rect 26620 4576 27169 4604
rect 26513 4567 26571 4573
rect 27157 4573 27169 4576
rect 27203 4573 27215 4607
rect 27157 4567 27215 4573
rect 28537 4607 28595 4613
rect 28537 4573 28549 4607
rect 28583 4573 28595 4607
rect 28537 4567 28595 4573
rect 20947 4508 22600 4536
rect 22649 4539 22707 4545
rect 20947 4505 20959 4508
rect 20901 4499 20959 4505
rect 22649 4505 22661 4539
rect 22695 4536 22707 4539
rect 22738 4536 22744 4548
rect 22695 4508 22744 4536
rect 22695 4505 22707 4508
rect 22649 4499 22707 4505
rect 22738 4496 22744 4508
rect 22796 4496 22802 4548
rect 23661 4539 23719 4545
rect 23661 4505 23673 4539
rect 23707 4536 23719 4539
rect 25041 4539 25099 4545
rect 25041 4536 25053 4539
rect 23707 4508 25053 4536
rect 23707 4505 23719 4508
rect 23661 4499 23719 4505
rect 25041 4505 25053 4508
rect 25087 4536 25099 4539
rect 25498 4536 25504 4548
rect 25087 4508 25504 4536
rect 25087 4505 25099 4508
rect 25041 4499 25099 4505
rect 25498 4496 25504 4508
rect 25556 4496 25562 4548
rect 25590 4496 25596 4548
rect 25648 4536 25654 4548
rect 26234 4536 26240 4548
rect 25648 4508 26240 4536
rect 25648 4496 25654 4508
rect 26234 4496 26240 4508
rect 26292 4496 26298 4548
rect 26528 4536 26556 4567
rect 28718 4564 28724 4616
rect 28776 4604 28782 4616
rect 29825 4607 29883 4613
rect 29825 4604 29837 4607
rect 28776 4576 29837 4604
rect 28776 4564 28782 4576
rect 29825 4573 29837 4576
rect 29871 4604 29883 4607
rect 30469 4607 30527 4613
rect 30469 4604 30481 4607
rect 29871 4576 30481 4604
rect 29871 4573 29883 4576
rect 29825 4567 29883 4573
rect 30469 4573 30481 4576
rect 30515 4604 30527 4607
rect 30558 4604 30564 4616
rect 30515 4576 30564 4604
rect 30515 4573 30527 4576
rect 30469 4567 30527 4573
rect 30558 4564 30564 4576
rect 30616 4564 30622 4616
rect 30653 4607 30711 4613
rect 30653 4573 30665 4607
rect 30699 4573 30711 4607
rect 30653 4567 30711 4573
rect 27062 4536 27068 4548
rect 26528 4508 27068 4536
rect 27062 4496 27068 4508
rect 27120 4496 27126 4548
rect 27614 4545 27620 4548
rect 27571 4539 27620 4545
rect 27571 4505 27583 4539
rect 27617 4505 27620 4539
rect 27571 4499 27620 4505
rect 27614 4496 27620 4499
rect 27672 4496 27678 4548
rect 28626 4496 28632 4548
rect 28684 4536 28690 4548
rect 28905 4539 28963 4545
rect 28905 4536 28917 4539
rect 28684 4508 28917 4536
rect 28684 4496 28690 4508
rect 28905 4505 28917 4508
rect 28951 4505 28963 4539
rect 28905 4499 28963 4505
rect 21450 4468 21456 4480
rect 20640 4440 21456 4468
rect 21450 4428 21456 4440
rect 21508 4428 21514 4480
rect 23293 4471 23351 4477
rect 23293 4437 23305 4471
rect 23339 4468 23351 4471
rect 23566 4468 23572 4480
rect 23339 4440 23572 4468
rect 23339 4437 23351 4440
rect 23293 4431 23351 4437
rect 23566 4428 23572 4440
rect 23624 4428 23630 4480
rect 23750 4428 23756 4480
rect 23808 4468 23814 4480
rect 23808 4440 23853 4468
rect 23808 4428 23814 4440
rect 23934 4428 23940 4480
rect 23992 4468 23998 4480
rect 28644 4468 28672 4496
rect 23992 4440 28672 4468
rect 23992 4428 23998 4440
rect 28810 4428 28816 4480
rect 28868 4468 28874 4480
rect 29917 4471 29975 4477
rect 29917 4468 29929 4471
rect 28868 4440 29929 4468
rect 28868 4428 28874 4440
rect 29917 4437 29929 4440
rect 29963 4437 29975 4471
rect 29917 4431 29975 4437
rect 30006 4428 30012 4480
rect 30064 4468 30070 4480
rect 30668 4468 30696 4567
rect 32214 4564 32220 4616
rect 32272 4604 32278 4616
rect 32585 4607 32643 4613
rect 32585 4604 32597 4607
rect 32272 4576 32597 4604
rect 32272 4564 32278 4576
rect 32585 4573 32597 4576
rect 32631 4573 32643 4607
rect 32585 4567 32643 4573
rect 33134 4564 33140 4616
rect 33192 4604 33198 4616
rect 33520 4613 33548 4712
rect 36538 4700 36544 4752
rect 36596 4740 36602 4752
rect 36814 4740 36820 4752
rect 36596 4712 36820 4740
rect 36596 4700 36602 4712
rect 36814 4700 36820 4712
rect 36872 4740 36878 4752
rect 37752 4740 37780 4780
rect 40770 4768 40776 4780
rect 40828 4768 40834 4820
rect 42444 4780 43576 4808
rect 40310 4740 40316 4752
rect 36872 4712 37780 4740
rect 38304 4712 40316 4740
rect 36872 4700 36878 4712
rect 37366 4632 37372 4684
rect 37424 4672 37430 4684
rect 37918 4672 37924 4684
rect 37424 4644 37924 4672
rect 37424 4632 37430 4644
rect 37918 4632 37924 4644
rect 37976 4632 37982 4684
rect 33321 4607 33379 4613
rect 33321 4604 33333 4607
rect 33192 4576 33333 4604
rect 33192 4564 33198 4576
rect 33321 4573 33333 4576
rect 33367 4573 33379 4607
rect 33321 4567 33379 4573
rect 33505 4607 33563 4613
rect 33505 4573 33517 4607
rect 33551 4573 33563 4607
rect 33505 4567 33563 4573
rect 35529 4607 35587 4613
rect 35529 4573 35541 4607
rect 35575 4604 35587 4607
rect 35618 4604 35624 4616
rect 35575 4576 35624 4604
rect 35575 4573 35587 4576
rect 35529 4567 35587 4573
rect 35618 4564 35624 4576
rect 35676 4564 35682 4616
rect 35796 4607 35854 4613
rect 35796 4573 35808 4607
rect 35842 4604 35854 4607
rect 37826 4604 37832 4616
rect 35842 4576 37832 4604
rect 35842 4573 35854 4576
rect 35796 4567 35854 4573
rect 37826 4564 37832 4576
rect 37884 4564 37890 4616
rect 38304 4613 38332 4712
rect 40310 4700 40316 4712
rect 40368 4700 40374 4752
rect 38841 4675 38899 4681
rect 38841 4641 38853 4675
rect 38887 4672 38899 4675
rect 39022 4672 39028 4684
rect 38887 4644 39028 4672
rect 38887 4641 38899 4644
rect 38841 4635 38899 4641
rect 39022 4632 39028 4644
rect 39080 4632 39086 4684
rect 39482 4632 39488 4684
rect 39540 4672 39546 4684
rect 42444 4681 42472 4780
rect 43346 4740 43352 4752
rect 42536 4712 43352 4740
rect 41693 4675 41751 4681
rect 41693 4672 41705 4675
rect 39540 4644 41705 4672
rect 39540 4632 39546 4644
rect 41693 4641 41705 4644
rect 41739 4641 41751 4675
rect 41693 4635 41751 4641
rect 42429 4675 42487 4681
rect 42429 4641 42441 4675
rect 42475 4641 42487 4675
rect 42429 4635 42487 4641
rect 38289 4607 38347 4613
rect 38289 4573 38301 4607
rect 38335 4573 38347 4607
rect 40865 4607 40923 4613
rect 40865 4604 40877 4607
rect 38289 4567 38347 4573
rect 38396 4576 40877 4604
rect 31110 4496 31116 4548
rect 31168 4536 31174 4548
rect 31168 4508 32444 4536
rect 31168 4496 31174 4508
rect 30064 4440 30696 4468
rect 30064 4428 30070 4440
rect 31570 4428 31576 4480
rect 31628 4468 31634 4480
rect 32214 4468 32220 4480
rect 31628 4440 32220 4468
rect 31628 4428 31634 4440
rect 32214 4428 32220 4440
rect 32272 4428 32278 4480
rect 32416 4468 32444 4508
rect 32490 4496 32496 4548
rect 32548 4536 32554 4548
rect 34514 4536 34520 4548
rect 32548 4508 34520 4536
rect 32548 4496 32554 4508
rect 34514 4496 34520 4508
rect 34572 4496 34578 4548
rect 37182 4496 37188 4548
rect 37240 4536 37246 4548
rect 37553 4539 37611 4545
rect 37553 4536 37565 4539
rect 37240 4508 37565 4536
rect 37240 4496 37246 4508
rect 37553 4505 37565 4508
rect 37599 4505 37611 4539
rect 37553 4499 37611 4505
rect 38194 4496 38200 4548
rect 38252 4536 38258 4548
rect 38396 4536 38424 4576
rect 40865 4573 40877 4576
rect 40911 4573 40923 4607
rect 40865 4567 40923 4573
rect 40954 4564 40960 4616
rect 41012 4604 41018 4616
rect 42337 4607 42395 4613
rect 42337 4604 42349 4607
rect 41012 4576 42349 4604
rect 41012 4564 41018 4576
rect 42337 4573 42349 4576
rect 42383 4604 42395 4607
rect 42536 4604 42564 4712
rect 43346 4700 43352 4712
rect 43404 4700 43410 4752
rect 43548 4740 43576 4780
rect 43622 4768 43628 4820
rect 43680 4808 43686 4820
rect 44177 4811 44235 4817
rect 44177 4808 44189 4811
rect 43680 4780 44189 4808
rect 43680 4768 43686 4780
rect 44177 4777 44189 4780
rect 44223 4777 44235 4811
rect 44177 4771 44235 4777
rect 44266 4768 44272 4820
rect 44324 4808 44330 4820
rect 45373 4811 45431 4817
rect 45373 4808 45385 4811
rect 44324 4780 45385 4808
rect 44324 4768 44330 4780
rect 45373 4777 45385 4780
rect 45419 4777 45431 4811
rect 45373 4771 45431 4777
rect 56502 4768 56508 4820
rect 56560 4808 56566 4820
rect 58253 4811 58311 4817
rect 58253 4808 58265 4811
rect 56560 4780 58265 4808
rect 56560 4768 56566 4780
rect 58253 4777 58265 4780
rect 58299 4777 58311 4811
rect 58253 4771 58311 4777
rect 50706 4740 50712 4752
rect 43548 4712 50712 4740
rect 50706 4700 50712 4712
rect 50764 4700 50770 4752
rect 42613 4675 42671 4681
rect 42613 4641 42625 4675
rect 42659 4641 42671 4675
rect 42613 4635 42671 4641
rect 42383 4576 42564 4604
rect 42383 4573 42395 4576
rect 42337 4567 42395 4573
rect 38252 4508 38424 4536
rect 38252 4496 38258 4508
rect 38746 4496 38752 4548
rect 38804 4536 38810 4548
rect 40126 4536 40132 4548
rect 38804 4508 39344 4536
rect 40087 4508 40132 4536
rect 38804 4496 38810 4508
rect 33410 4468 33416 4480
rect 32416 4440 33416 4468
rect 33410 4428 33416 4440
rect 33468 4428 33474 4480
rect 33502 4428 33508 4480
rect 33560 4468 33566 4480
rect 33689 4471 33747 4477
rect 33689 4468 33701 4471
rect 33560 4440 33701 4468
rect 33560 4428 33566 4440
rect 33689 4437 33701 4440
rect 33735 4437 33747 4471
rect 33689 4431 33747 4437
rect 36354 4428 36360 4480
rect 36412 4468 36418 4480
rect 36909 4471 36967 4477
rect 36909 4468 36921 4471
rect 36412 4440 36921 4468
rect 36412 4428 36418 4440
rect 36909 4437 36921 4440
rect 36955 4437 36967 4471
rect 36909 4431 36967 4437
rect 37458 4428 37464 4480
rect 37516 4468 37522 4480
rect 39206 4468 39212 4480
rect 37516 4440 39212 4468
rect 37516 4428 37522 4440
rect 39206 4428 39212 4440
rect 39264 4428 39270 4480
rect 39316 4468 39344 4508
rect 40126 4496 40132 4508
rect 40184 4496 40190 4548
rect 40770 4496 40776 4548
rect 40828 4536 40834 4548
rect 42518 4536 42524 4548
rect 40828 4508 42524 4536
rect 40828 4496 40834 4508
rect 42518 4496 42524 4508
rect 42576 4536 42582 4548
rect 42628 4536 42656 4635
rect 42978 4632 42984 4684
rect 43036 4672 43042 4684
rect 43036 4644 43852 4672
rect 43036 4632 43042 4644
rect 42705 4607 42763 4613
rect 42705 4573 42717 4607
rect 42751 4573 42763 4607
rect 43622 4604 43628 4616
rect 43583 4576 43628 4604
rect 42705 4567 42763 4573
rect 42576 4508 42656 4536
rect 42576 4496 42582 4508
rect 40221 4471 40279 4477
rect 40221 4468 40233 4471
rect 39316 4440 40233 4468
rect 40221 4437 40233 4440
rect 40267 4437 40279 4471
rect 40221 4431 40279 4437
rect 40310 4428 40316 4480
rect 40368 4468 40374 4480
rect 40957 4471 41015 4477
rect 40957 4468 40969 4471
rect 40368 4440 40969 4468
rect 40368 4428 40374 4440
rect 40957 4437 40969 4440
rect 41003 4437 41015 4471
rect 42720 4468 42748 4567
rect 43622 4564 43628 4576
rect 43680 4564 43686 4616
rect 43824 4613 43852 4644
rect 43898 4632 43904 4684
rect 43956 4672 43962 4684
rect 53098 4672 53104 4684
rect 43956 4644 53104 4672
rect 43956 4632 43962 4644
rect 53098 4632 53104 4644
rect 53156 4632 53162 4684
rect 43809 4607 43867 4613
rect 43809 4573 43821 4607
rect 43855 4573 43867 4607
rect 43809 4567 43867 4573
rect 43990 4564 43996 4616
rect 44048 4613 44054 4616
rect 44048 4604 44056 4613
rect 46201 4607 46259 4613
rect 46201 4604 46213 4607
rect 44048 4576 44093 4604
rect 45020 4576 46213 4604
rect 44048 4567 44056 4576
rect 44048 4564 44054 4567
rect 43901 4539 43959 4545
rect 43901 4505 43913 4539
rect 43947 4536 43959 4539
rect 45020 4536 45048 4576
rect 46201 4573 46213 4576
rect 46247 4573 46259 4607
rect 51258 4604 51264 4616
rect 51219 4576 51264 4604
rect 46201 4567 46259 4573
rect 51258 4564 51264 4576
rect 51316 4564 51322 4616
rect 51442 4604 51448 4616
rect 51403 4576 51448 4604
rect 51442 4564 51448 4576
rect 51500 4564 51506 4616
rect 57790 4564 57796 4616
rect 57848 4604 57854 4616
rect 58069 4607 58127 4613
rect 58069 4604 58081 4607
rect 57848 4576 58081 4604
rect 57848 4564 57854 4576
rect 58069 4573 58081 4576
rect 58115 4573 58127 4607
rect 58069 4567 58127 4573
rect 43947 4508 45048 4536
rect 43947 4505 43959 4508
rect 43901 4499 43959 4505
rect 45094 4496 45100 4548
rect 45152 4536 45158 4548
rect 45281 4539 45339 4545
rect 45281 4536 45293 4539
rect 45152 4508 45293 4536
rect 45152 4496 45158 4508
rect 45281 4505 45293 4508
rect 45327 4505 45339 4539
rect 46014 4536 46020 4548
rect 45975 4508 46020 4536
rect 45281 4499 45339 4505
rect 46014 4496 46020 4508
rect 46072 4496 46078 4548
rect 44358 4468 44364 4480
rect 42720 4440 44364 4468
rect 40957 4431 41015 4437
rect 44358 4428 44364 4440
rect 44416 4428 44422 4480
rect 51629 4471 51687 4477
rect 51629 4437 51641 4471
rect 51675 4468 51687 4471
rect 53558 4468 53564 4480
rect 51675 4440 53564 4468
rect 51675 4437 51687 4440
rect 51629 4431 51687 4437
rect 53558 4428 53564 4440
rect 53616 4428 53622 4480
rect 1104 4378 58880 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 58880 4378
rect 1104 4304 58880 4326
rect 7006 4224 7012 4276
rect 7064 4264 7070 4276
rect 7064 4236 14504 4264
rect 7064 4224 7070 4236
rect 5813 4199 5871 4205
rect 5813 4165 5825 4199
rect 5859 4196 5871 4199
rect 6454 4196 6460 4208
rect 5859 4168 6460 4196
rect 5859 4165 5871 4168
rect 5813 4159 5871 4165
rect 6454 4156 6460 4168
rect 6512 4156 6518 4208
rect 6641 4199 6699 4205
rect 6641 4165 6653 4199
rect 6687 4196 6699 4199
rect 7282 4196 7288 4208
rect 6687 4168 7288 4196
rect 6687 4165 6699 4168
rect 6641 4159 6699 4165
rect 7282 4156 7288 4168
rect 7340 4156 7346 4208
rect 7377 4199 7435 4205
rect 7377 4165 7389 4199
rect 7423 4196 7435 4199
rect 8478 4196 8484 4208
rect 7423 4168 8484 4196
rect 7423 4165 7435 4168
rect 7377 4159 7435 4165
rect 8478 4156 8484 4168
rect 8536 4156 8542 4208
rect 9582 4196 9588 4208
rect 8588 4168 9588 4196
rect 1581 4131 1639 4137
rect 1581 4097 1593 4131
rect 1627 4128 1639 4131
rect 5902 4128 5908 4140
rect 1627 4100 5908 4128
rect 1627 4097 1639 4100
rect 1581 4091 1639 4097
rect 5902 4088 5908 4100
rect 5960 4088 5966 4140
rect 6822 4128 6828 4140
rect 6783 4100 6828 4128
rect 6822 4088 6828 4100
rect 6880 4088 6886 4140
rect 8021 4131 8079 4137
rect 8021 4097 8033 4131
rect 8067 4128 8079 4131
rect 8202 4128 8208 4140
rect 8067 4100 8208 4128
rect 8067 4097 8079 4100
rect 8021 4091 8079 4097
rect 8202 4088 8208 4100
rect 8260 4128 8266 4140
rect 8588 4128 8616 4168
rect 9324 4137 9352 4168
rect 9582 4156 9588 4168
rect 9640 4156 9646 4208
rect 10965 4199 11023 4205
rect 10965 4165 10977 4199
rect 11011 4196 11023 4199
rect 11698 4196 11704 4208
rect 11011 4168 11704 4196
rect 11011 4165 11023 4168
rect 10965 4159 11023 4165
rect 11698 4156 11704 4168
rect 11756 4156 11762 4208
rect 11793 4199 11851 4205
rect 11793 4165 11805 4199
rect 11839 4196 11851 4199
rect 12434 4196 12440 4208
rect 11839 4168 12440 4196
rect 11839 4165 11851 4168
rect 11793 4159 11851 4165
rect 12434 4156 12440 4168
rect 12492 4156 12498 4208
rect 13357 4199 13415 4205
rect 13357 4196 13369 4199
rect 12636 4168 13369 4196
rect 8260 4100 8616 4128
rect 9309 4131 9367 4137
rect 8260 4088 8266 4100
rect 9309 4097 9321 4131
rect 9355 4097 9367 4131
rect 9309 4091 9367 4097
rect 9490 4088 9496 4140
rect 9548 4128 9554 4140
rect 11146 4128 11152 4140
rect 9548 4100 10456 4128
rect 11107 4100 11152 4128
rect 9548 4088 9554 4100
rect 1762 4060 1768 4072
rect 1723 4032 1768 4060
rect 1762 4020 1768 4032
rect 1820 4020 1826 4072
rect 8481 4063 8539 4069
rect 8481 4029 8493 4063
rect 8527 4060 8539 4063
rect 8527 4032 8892 4060
rect 8527 4029 8539 4032
rect 8481 4023 8539 4029
rect 5997 3995 6055 4001
rect 5997 3961 6009 3995
rect 6043 3992 6055 3995
rect 6638 3992 6644 4004
rect 6043 3964 6644 3992
rect 6043 3961 6055 3964
rect 5997 3955 6055 3961
rect 6638 3952 6644 3964
rect 6696 3952 6702 4004
rect 8389 3995 8447 4001
rect 8389 3961 8401 3995
rect 8435 3992 8447 3995
rect 8662 3992 8668 4004
rect 8435 3964 8668 3992
rect 8435 3961 8447 3964
rect 8389 3955 8447 3961
rect 8662 3952 8668 3964
rect 8720 3952 8726 4004
rect 8864 3992 8892 4032
rect 8938 4020 8944 4072
rect 8996 4060 9002 4072
rect 9125 4063 9183 4069
rect 9125 4060 9137 4063
rect 8996 4032 9137 4060
rect 8996 4020 9002 4032
rect 9125 4029 9137 4032
rect 9171 4029 9183 4063
rect 9125 4023 9183 4029
rect 9214 4020 9220 4072
rect 9272 4060 9278 4072
rect 9272 4032 9317 4060
rect 9272 4020 9278 4032
rect 9398 4020 9404 4072
rect 9456 4060 9462 4072
rect 9456 4032 9501 4060
rect 9456 4020 9462 4032
rect 9582 4020 9588 4072
rect 9640 4060 9646 4072
rect 9953 4063 10011 4069
rect 9953 4060 9965 4063
rect 9640 4032 9965 4060
rect 9640 4020 9646 4032
rect 9953 4029 9965 4032
rect 9999 4060 10011 4063
rect 10318 4060 10324 4072
rect 9999 4032 10324 4060
rect 9999 4029 10011 4032
rect 9953 4023 10011 4029
rect 10318 4020 10324 4032
rect 10376 4020 10382 4072
rect 10428 4069 10456 4100
rect 11146 4088 11152 4100
rect 11204 4088 11210 4140
rect 11977 4131 12035 4137
rect 11977 4097 11989 4131
rect 12023 4128 12035 4131
rect 12066 4128 12072 4140
rect 12023 4100 12072 4128
rect 12023 4097 12035 4100
rect 11977 4091 12035 4097
rect 12066 4088 12072 4100
rect 12124 4088 12130 4140
rect 12636 4128 12664 4168
rect 13357 4165 13369 4168
rect 13403 4196 13415 4199
rect 14274 4196 14280 4208
rect 13403 4168 14280 4196
rect 13403 4165 13415 4168
rect 13357 4159 13415 4165
rect 14274 4156 14280 4168
rect 14332 4156 14338 4208
rect 14476 4196 14504 4236
rect 16574 4224 16580 4276
rect 16632 4264 16638 4276
rect 19334 4264 19340 4276
rect 16632 4236 19340 4264
rect 16632 4224 16638 4236
rect 19334 4224 19340 4236
rect 19392 4224 19398 4276
rect 22370 4224 22376 4276
rect 22428 4264 22434 4276
rect 24118 4264 24124 4276
rect 22428 4236 24124 4264
rect 22428 4224 22434 4236
rect 24118 4224 24124 4236
rect 24176 4224 24182 4276
rect 24670 4264 24676 4276
rect 24631 4236 24676 4264
rect 24670 4224 24676 4236
rect 24728 4224 24734 4276
rect 26421 4267 26479 4273
rect 26421 4233 26433 4267
rect 26467 4264 26479 4267
rect 27798 4264 27804 4276
rect 26467 4236 27804 4264
rect 26467 4233 26479 4236
rect 26421 4227 26479 4233
rect 27798 4224 27804 4236
rect 27856 4224 27862 4276
rect 27982 4224 27988 4276
rect 28040 4264 28046 4276
rect 31570 4264 31576 4276
rect 28040 4236 31576 4264
rect 28040 4224 28046 4236
rect 31570 4224 31576 4236
rect 31628 4224 31634 4276
rect 32677 4267 32735 4273
rect 32677 4233 32689 4267
rect 32723 4264 32735 4267
rect 33318 4264 33324 4276
rect 32723 4236 33324 4264
rect 32723 4233 32735 4236
rect 32677 4227 32735 4233
rect 33318 4224 33324 4236
rect 33376 4264 33382 4276
rect 33686 4264 33692 4276
rect 33376 4236 33692 4264
rect 33376 4224 33382 4236
rect 33686 4224 33692 4236
rect 33744 4224 33750 4276
rect 34146 4224 34152 4276
rect 34204 4264 34210 4276
rect 52454 4264 52460 4276
rect 34204 4236 52460 4264
rect 34204 4224 34210 4236
rect 52454 4224 52460 4236
rect 52512 4224 52518 4276
rect 53098 4264 53104 4276
rect 53059 4236 53104 4264
rect 53098 4224 53104 4236
rect 53156 4224 53162 4276
rect 19518 4196 19524 4208
rect 14476 4168 19524 4196
rect 19518 4156 19524 4168
rect 19576 4156 19582 4208
rect 20248 4199 20306 4205
rect 20248 4165 20260 4199
rect 20294 4196 20306 4199
rect 20530 4196 20536 4208
rect 20294 4168 20536 4196
rect 20294 4165 20306 4168
rect 20248 4159 20306 4165
rect 20530 4156 20536 4168
rect 20588 4156 20594 4208
rect 24854 4196 24860 4208
rect 21284 4168 24860 4196
rect 15841 4131 15899 4137
rect 12452 4100 12664 4128
rect 12728 4100 13676 4128
rect 10413 4063 10471 4069
rect 10413 4029 10425 4063
rect 10459 4029 10471 4063
rect 10413 4023 10471 4029
rect 12342 4020 12348 4072
rect 12400 4060 12406 4072
rect 12452 4069 12480 4100
rect 12437 4063 12495 4069
rect 12437 4060 12449 4063
rect 12400 4032 12449 4060
rect 12400 4020 12406 4032
rect 12437 4029 12449 4032
rect 12483 4029 12495 4063
rect 12437 4023 12495 4029
rect 10042 3992 10048 4004
rect 8864 3964 10048 3992
rect 10042 3952 10048 3964
rect 10100 3952 10106 4004
rect 10229 3995 10287 4001
rect 10229 3961 10241 3995
rect 10275 3961 10287 3995
rect 10229 3955 10287 3961
rect 7466 3924 7472 3936
rect 7427 3896 7472 3924
rect 7466 3884 7472 3896
rect 7524 3884 7530 3936
rect 8570 3884 8576 3936
rect 8628 3924 8634 3936
rect 8941 3927 8999 3933
rect 8941 3924 8953 3927
rect 8628 3896 8953 3924
rect 8628 3884 8634 3896
rect 8941 3893 8953 3896
rect 8987 3893 8999 3927
rect 8941 3887 8999 3893
rect 9030 3884 9036 3936
rect 9088 3924 9094 3936
rect 10244 3924 10272 3955
rect 11238 3952 11244 4004
rect 11296 3992 11302 4004
rect 12728 3992 12756 4100
rect 12894 4060 12900 4072
rect 12855 4032 12900 4060
rect 12894 4020 12900 4032
rect 12952 4020 12958 4072
rect 11296 3964 12756 3992
rect 12805 3995 12863 4001
rect 11296 3952 11302 3964
rect 12805 3961 12817 3995
rect 12851 3992 12863 3995
rect 12986 3992 12992 4004
rect 12851 3964 12992 3992
rect 12851 3961 12863 3964
rect 12805 3955 12863 3961
rect 12986 3952 12992 3964
rect 13044 3952 13050 4004
rect 13648 4001 13676 4100
rect 15841 4097 15853 4131
rect 15887 4097 15899 4131
rect 16942 4128 16948 4140
rect 16903 4100 16948 4128
rect 15841 4091 15899 4097
rect 14737 4063 14795 4069
rect 14737 4029 14749 4063
rect 14783 4060 14795 4063
rect 14826 4060 14832 4072
rect 14783 4032 14832 4060
rect 14783 4029 14795 4032
rect 14737 4023 14795 4029
rect 14826 4020 14832 4032
rect 14884 4020 14890 4072
rect 13633 3995 13691 4001
rect 13633 3961 13645 3995
rect 13679 3961 13691 3995
rect 14553 3995 14611 4001
rect 14553 3992 14565 3995
rect 13633 3955 13691 3961
rect 13740 3964 14565 3992
rect 9088 3896 10272 3924
rect 9088 3884 9094 3896
rect 11146 3884 11152 3936
rect 11204 3924 11210 3936
rect 13740 3924 13768 3964
rect 14553 3961 14565 3964
rect 14599 3961 14611 3995
rect 15856 3992 15884 4091
rect 16942 4088 16948 4100
rect 17000 4088 17006 4140
rect 17586 4088 17592 4140
rect 17644 4128 17650 4140
rect 17865 4131 17923 4137
rect 17865 4128 17877 4131
rect 17644 4100 17877 4128
rect 17644 4088 17650 4100
rect 17865 4097 17877 4100
rect 17911 4097 17923 4131
rect 18598 4128 18604 4140
rect 17865 4091 17923 4097
rect 17972 4100 18604 4128
rect 16114 4060 16120 4072
rect 16075 4032 16120 4060
rect 16114 4020 16120 4032
rect 16172 4020 16178 4072
rect 17221 4063 17279 4069
rect 17221 4029 17233 4063
rect 17267 4060 17279 4063
rect 17972 4060 18000 4100
rect 18598 4088 18604 4100
rect 18656 4088 18662 4140
rect 19058 4088 19064 4140
rect 19116 4128 19122 4140
rect 19153 4131 19211 4137
rect 19153 4128 19165 4131
rect 19116 4100 19165 4128
rect 19116 4088 19122 4100
rect 19153 4097 19165 4100
rect 19199 4097 19211 4131
rect 19610 4128 19616 4140
rect 19153 4091 19211 4097
rect 19260 4100 19616 4128
rect 17267 4032 18000 4060
rect 18141 4063 18199 4069
rect 17267 4029 17279 4032
rect 17221 4023 17279 4029
rect 18141 4029 18153 4063
rect 18187 4060 18199 4063
rect 18506 4060 18512 4072
rect 18187 4032 18512 4060
rect 18187 4029 18199 4032
rect 18141 4023 18199 4029
rect 18506 4020 18512 4032
rect 18564 4020 18570 4072
rect 19260 4069 19288 4100
rect 19610 4088 19616 4100
rect 19668 4088 19674 4140
rect 19794 4088 19800 4140
rect 19852 4128 19858 4140
rect 20990 4128 20996 4140
rect 19852 4100 20996 4128
rect 19852 4088 19858 4100
rect 20990 4088 20996 4100
rect 21048 4088 21054 4140
rect 19245 4063 19303 4069
rect 19245 4060 19257 4063
rect 19155 4032 19257 4060
rect 19245 4029 19257 4032
rect 19291 4029 19303 4063
rect 19245 4023 19303 4029
rect 19337 4063 19395 4069
rect 19337 4029 19349 4063
rect 19383 4060 19395 4063
rect 19426 4060 19432 4072
rect 19383 4032 19432 4060
rect 19383 4029 19395 4032
rect 19337 4023 19395 4029
rect 15856 3964 18920 3992
rect 14553 3955 14611 3961
rect 11204 3896 13768 3924
rect 13817 3927 13875 3933
rect 11204 3884 11210 3896
rect 13817 3893 13829 3927
rect 13863 3924 13875 3927
rect 16758 3924 16764 3936
rect 13863 3896 16764 3924
rect 13863 3893 13875 3896
rect 13817 3887 13875 3893
rect 16758 3884 16764 3896
rect 16816 3884 16822 3936
rect 18138 3884 18144 3936
rect 18196 3924 18202 3936
rect 18414 3924 18420 3936
rect 18196 3896 18420 3924
rect 18196 3884 18202 3896
rect 18414 3884 18420 3896
rect 18472 3884 18478 3936
rect 18782 3924 18788 3936
rect 18743 3896 18788 3924
rect 18782 3884 18788 3896
rect 18840 3884 18846 3936
rect 18892 3924 18920 3964
rect 18966 3952 18972 4004
rect 19024 3992 19030 4004
rect 19260 3992 19288 4023
rect 19426 4020 19432 4032
rect 19484 4020 19490 4072
rect 19978 4060 19984 4072
rect 19939 4032 19984 4060
rect 19978 4020 19984 4032
rect 20036 4020 20042 4072
rect 19024 3964 19288 3992
rect 19024 3952 19030 3964
rect 19426 3924 19432 3936
rect 18892 3896 19432 3924
rect 19426 3884 19432 3896
rect 19484 3884 19490 3936
rect 19610 3884 19616 3936
rect 19668 3924 19674 3936
rect 21284 3924 21312 4168
rect 24854 4156 24860 4168
rect 24912 4156 24918 4208
rect 27608 4199 27666 4205
rect 27608 4165 27620 4199
rect 27654 4196 27666 4199
rect 28074 4196 28080 4208
rect 27654 4168 28080 4196
rect 27654 4165 27666 4168
rect 27608 4159 27666 4165
rect 28074 4156 28080 4168
rect 28132 4156 28138 4208
rect 28166 4156 28172 4208
rect 28224 4196 28230 4208
rect 28224 4168 28580 4196
rect 28224 4156 28230 4168
rect 22370 4128 22376 4140
rect 22331 4100 22376 4128
rect 22370 4088 22376 4100
rect 22428 4088 22434 4140
rect 23566 4137 23572 4140
rect 23560 4128 23572 4137
rect 23527 4100 23572 4128
rect 23560 4091 23572 4100
rect 23566 4088 23572 4091
rect 23624 4088 23630 4140
rect 25133 4131 25191 4137
rect 25133 4097 25145 4131
rect 25179 4128 25191 4131
rect 28442 4128 28448 4140
rect 25179 4100 28448 4128
rect 25179 4097 25191 4100
rect 25133 4091 25191 4097
rect 28442 4088 28448 4100
rect 28500 4088 28506 4140
rect 28552 4128 28580 4168
rect 29564 4168 29868 4196
rect 29564 4128 29592 4168
rect 29730 4128 29736 4140
rect 28552 4100 29592 4128
rect 29691 4100 29736 4128
rect 29730 4088 29736 4100
rect 29788 4088 29794 4140
rect 29840 4128 29868 4168
rect 30466 4156 30472 4208
rect 30524 4196 30530 4208
rect 30745 4199 30803 4205
rect 30745 4196 30757 4199
rect 30524 4168 30757 4196
rect 30524 4156 30530 4168
rect 30745 4165 30757 4168
rect 30791 4196 30803 4199
rect 30926 4196 30932 4208
rect 30791 4168 30932 4196
rect 30791 4165 30803 4168
rect 30745 4159 30803 4165
rect 30926 4156 30932 4168
rect 30984 4156 30990 4208
rect 33410 4156 33416 4208
rect 33468 4196 33474 4208
rect 37366 4196 37372 4208
rect 33468 4168 37372 4196
rect 33468 4156 33474 4168
rect 37366 4156 37372 4168
rect 37424 4156 37430 4208
rect 37642 4156 37648 4208
rect 37700 4196 37706 4208
rect 41325 4199 41383 4205
rect 41325 4196 41337 4199
rect 37700 4168 41337 4196
rect 37700 4156 37706 4168
rect 41325 4165 41337 4168
rect 41371 4165 41383 4199
rect 41325 4159 41383 4165
rect 42058 4156 42064 4208
rect 42116 4196 42122 4208
rect 44453 4199 44511 4205
rect 44453 4196 44465 4199
rect 42116 4168 44465 4196
rect 42116 4156 42122 4168
rect 44453 4165 44465 4168
rect 44499 4165 44511 4199
rect 44453 4159 44511 4165
rect 45370 4156 45376 4208
rect 45428 4156 45434 4208
rect 46106 4156 46112 4208
rect 46164 4196 46170 4208
rect 46845 4199 46903 4205
rect 46845 4196 46857 4199
rect 46164 4168 46857 4196
rect 46164 4156 46170 4168
rect 46845 4165 46857 4168
rect 46891 4165 46903 4199
rect 46845 4159 46903 4165
rect 51994 4156 52000 4208
rect 52052 4196 52058 4208
rect 52181 4199 52239 4205
rect 52181 4196 52193 4199
rect 52052 4168 52193 4196
rect 52052 4156 52058 4168
rect 52181 4165 52193 4168
rect 52227 4165 52239 4199
rect 52181 4159 52239 4165
rect 52822 4156 52828 4208
rect 52880 4196 52886 4208
rect 53009 4199 53067 4205
rect 53009 4196 53021 4199
rect 52880 4168 53021 4196
rect 52880 4156 52886 4168
rect 53009 4165 53021 4168
rect 53055 4165 53067 4199
rect 53009 4159 53067 4165
rect 53374 4156 53380 4208
rect 53432 4196 53438 4208
rect 53745 4199 53803 4205
rect 53745 4196 53757 4199
rect 53432 4168 53757 4196
rect 53432 4156 53438 4168
rect 53745 4165 53757 4168
rect 53791 4165 53803 4199
rect 53745 4159 53803 4165
rect 57882 4156 57888 4208
rect 57940 4196 57946 4208
rect 58161 4199 58219 4205
rect 58161 4196 58173 4199
rect 57940 4168 58173 4196
rect 57940 4156 57946 4168
rect 58161 4165 58173 4168
rect 58207 4165 58219 4199
rect 58161 4159 58219 4165
rect 31202 4128 31208 4140
rect 29840 4100 31208 4128
rect 31202 4088 31208 4100
rect 31260 4088 31266 4140
rect 31478 4088 31484 4140
rect 31536 4128 31542 4140
rect 31573 4131 31631 4137
rect 31573 4128 31585 4131
rect 31536 4100 31585 4128
rect 31536 4088 31542 4100
rect 31573 4097 31585 4100
rect 31619 4128 31631 4131
rect 33505 4131 33563 4137
rect 33505 4128 33517 4131
rect 31619 4100 33517 4128
rect 31619 4097 31631 4100
rect 31573 4091 31631 4097
rect 33505 4097 33517 4100
rect 33551 4097 33563 4131
rect 34422 4128 34428 4140
rect 34383 4100 34428 4128
rect 33505 4091 33563 4097
rect 34422 4088 34428 4100
rect 34480 4088 34486 4140
rect 35345 4131 35403 4137
rect 35345 4128 35357 4131
rect 34532 4100 35357 4128
rect 22649 4063 22707 4069
rect 22649 4029 22661 4063
rect 22695 4060 22707 4063
rect 23014 4060 23020 4072
rect 22695 4032 23020 4060
rect 22695 4029 22707 4032
rect 22649 4023 22707 4029
rect 23014 4020 23020 4032
rect 23072 4020 23078 4072
rect 23290 4060 23296 4072
rect 23251 4032 23296 4060
rect 23290 4020 23296 4032
rect 23348 4020 23354 4072
rect 24670 4020 24676 4072
rect 24728 4060 24734 4072
rect 25317 4063 25375 4069
rect 25317 4060 25329 4063
rect 24728 4032 25329 4060
rect 24728 4020 24734 4032
rect 25317 4029 25329 4032
rect 25363 4029 25375 4063
rect 25317 4023 25375 4029
rect 27341 4063 27399 4069
rect 27341 4029 27353 4063
rect 27387 4029 27399 4063
rect 27341 4023 27399 4029
rect 24486 3952 24492 4004
rect 24544 3992 24550 4004
rect 27246 3992 27252 4004
rect 24544 3964 27252 3992
rect 24544 3952 24550 3964
rect 27246 3952 27252 3964
rect 27304 3952 27310 4004
rect 19668 3896 21312 3924
rect 19668 3884 19674 3896
rect 21358 3884 21364 3936
rect 21416 3924 21422 3936
rect 21416 3896 21461 3924
rect 21416 3884 21422 3896
rect 23198 3884 23204 3936
rect 23256 3924 23262 3936
rect 25958 3924 25964 3936
rect 23256 3896 25964 3924
rect 23256 3884 23262 3896
rect 25958 3884 25964 3896
rect 26016 3884 26022 3936
rect 27356 3924 27384 4023
rect 29638 4020 29644 4072
rect 29696 4060 29702 4072
rect 29917 4063 29975 4069
rect 29917 4060 29929 4063
rect 29696 4032 29929 4060
rect 29696 4020 29702 4032
rect 29917 4029 29929 4032
rect 29963 4029 29975 4063
rect 32766 4060 32772 4072
rect 32727 4032 32772 4060
rect 29917 4023 29975 4029
rect 32766 4020 32772 4032
rect 32824 4020 32830 4072
rect 32858 4020 32864 4072
rect 32916 4060 32922 4072
rect 33689 4063 33747 4069
rect 32916 4032 32961 4060
rect 32916 4020 32922 4032
rect 33689 4029 33701 4063
rect 33735 4029 33747 4063
rect 33689 4023 33747 4029
rect 28994 3992 29000 4004
rect 28276 3964 29000 3992
rect 28276 3924 28304 3964
rect 28994 3952 29000 3964
rect 29052 3992 29058 4004
rect 30098 3992 30104 4004
rect 29052 3964 30104 3992
rect 29052 3952 29058 3964
rect 30098 3952 30104 3964
rect 30156 3952 30162 4004
rect 31757 3995 31815 4001
rect 31757 3961 31769 3995
rect 31803 3992 31815 3995
rect 31803 3964 32628 3992
rect 31803 3961 31815 3964
rect 31757 3955 31815 3961
rect 28718 3924 28724 3936
rect 27356 3896 28304 3924
rect 28679 3896 28724 3924
rect 28718 3884 28724 3896
rect 28776 3884 28782 3936
rect 30834 3924 30840 3936
rect 30795 3896 30840 3924
rect 30834 3884 30840 3896
rect 30892 3884 30898 3936
rect 32030 3884 32036 3936
rect 32088 3924 32094 3936
rect 32309 3927 32367 3933
rect 32309 3924 32321 3927
rect 32088 3896 32321 3924
rect 32088 3884 32094 3896
rect 32309 3893 32321 3896
rect 32355 3893 32367 3927
rect 32600 3924 32628 3964
rect 32674 3952 32680 4004
rect 32732 3992 32738 4004
rect 33704 3992 33732 4023
rect 34054 4020 34060 4072
rect 34112 4060 34118 4072
rect 34532 4060 34560 4100
rect 35345 4097 35357 4100
rect 35391 4097 35403 4131
rect 36262 4128 36268 4140
rect 36223 4100 36268 4128
rect 35345 4091 35403 4097
rect 36262 4088 36268 4100
rect 36320 4088 36326 4140
rect 37182 4088 37188 4140
rect 37240 4128 37246 4140
rect 38838 4137 38844 4140
rect 37461 4131 37519 4137
rect 37461 4128 37473 4131
rect 37240 4100 37473 4128
rect 37240 4088 37246 4100
rect 37461 4097 37473 4100
rect 37507 4097 37519 4131
rect 37461 4091 37519 4097
rect 38832 4091 38844 4137
rect 38896 4128 38902 4140
rect 40126 4128 40132 4140
rect 38896 4100 38932 4128
rect 39592 4100 40132 4128
rect 38838 4088 38844 4091
rect 38896 4088 38902 4100
rect 34112 4032 34560 4060
rect 34609 4063 34667 4069
rect 34112 4020 34118 4032
rect 34609 4029 34621 4063
rect 34655 4029 34667 4063
rect 34609 4023 34667 4029
rect 35529 4063 35587 4069
rect 35529 4029 35541 4063
rect 35575 4029 35587 4063
rect 35529 4023 35587 4029
rect 32732 3964 33732 3992
rect 32732 3952 32738 3964
rect 33410 3924 33416 3936
rect 32600 3896 33416 3924
rect 32309 3887 32367 3893
rect 33410 3884 33416 3896
rect 33468 3884 33474 3936
rect 33594 3884 33600 3936
rect 33652 3924 33658 3936
rect 34624 3924 34652 4023
rect 33652 3896 34652 3924
rect 33652 3884 33658 3896
rect 35434 3884 35440 3936
rect 35492 3924 35498 3936
rect 35544 3924 35572 4023
rect 35710 4020 35716 4072
rect 35768 4060 35774 4072
rect 36449 4063 36507 4069
rect 36449 4060 36461 4063
rect 35768 4032 36461 4060
rect 35768 4020 35774 4032
rect 36449 4029 36461 4032
rect 36495 4029 36507 4063
rect 36449 4023 36507 4029
rect 36722 4020 36728 4072
rect 36780 4060 36786 4072
rect 37645 4063 37703 4069
rect 37645 4060 37657 4063
rect 36780 4032 37657 4060
rect 36780 4020 36786 4032
rect 37645 4029 37657 4032
rect 37691 4029 37703 4063
rect 37645 4023 37703 4029
rect 38565 4063 38623 4069
rect 38565 4029 38577 4063
rect 38611 4029 38623 4063
rect 38565 4023 38623 4029
rect 35618 3952 35624 4004
rect 35676 3992 35682 4004
rect 38580 3992 38608 4023
rect 35676 3964 38608 3992
rect 35676 3952 35682 3964
rect 35492 3896 35572 3924
rect 35492 3884 35498 3896
rect 37826 3884 37832 3936
rect 37884 3924 37890 3936
rect 39592 3924 39620 4100
rect 40126 4088 40132 4100
rect 40184 4088 40190 4140
rect 40586 4128 40592 4140
rect 40547 4100 40592 4128
rect 40586 4088 40592 4100
rect 40644 4088 40650 4140
rect 41506 4128 41512 4140
rect 41467 4100 41512 4128
rect 41506 4088 41512 4100
rect 41564 4088 41570 4140
rect 43346 4128 43352 4140
rect 43307 4100 43352 4128
rect 43346 4088 43352 4100
rect 43404 4088 43410 4140
rect 43717 4131 43775 4137
rect 43717 4097 43729 4131
rect 43763 4097 43775 4131
rect 43717 4091 43775 4097
rect 39850 4020 39856 4072
rect 39908 4060 39914 4072
rect 40773 4063 40831 4069
rect 40773 4060 40785 4063
rect 39908 4032 40785 4060
rect 39908 4020 39914 4032
rect 40773 4029 40785 4032
rect 40819 4029 40831 4063
rect 43438 4060 43444 4072
rect 43399 4032 43444 4060
rect 40773 4023 40831 4029
rect 43438 4020 43444 4032
rect 43496 4020 43502 4072
rect 43625 4063 43683 4069
rect 43625 4029 43637 4063
rect 43671 4029 43683 4063
rect 43625 4023 43683 4029
rect 39942 3992 39948 4004
rect 39903 3964 39948 3992
rect 39942 3952 39948 3964
rect 40000 3952 40006 4004
rect 42981 3995 43039 4001
rect 42981 3961 42993 3995
rect 43027 3992 43039 3995
rect 43530 3992 43536 4004
rect 43027 3964 43536 3992
rect 43027 3961 43039 3964
rect 42981 3955 43039 3961
rect 43530 3952 43536 3964
rect 43588 3952 43594 4004
rect 43640 3936 43668 4023
rect 43732 3992 43760 4091
rect 44358 4088 44364 4140
rect 44416 4128 44422 4140
rect 45189 4131 45247 4137
rect 44416 4100 44588 4128
rect 44416 4088 44422 4100
rect 44560 4060 44588 4100
rect 45189 4097 45201 4131
rect 45235 4128 45247 4131
rect 45388 4128 45416 4156
rect 45922 4128 45928 4140
rect 45235 4100 45416 4128
rect 45883 4100 45928 4128
rect 45235 4097 45247 4100
rect 45189 4091 45247 4097
rect 45922 4088 45928 4100
rect 45980 4088 45986 4140
rect 46661 4131 46719 4137
rect 46661 4097 46673 4131
rect 46707 4097 46719 4131
rect 46661 4091 46719 4097
rect 44637 4063 44695 4069
rect 44637 4060 44649 4063
rect 44560 4032 44649 4060
rect 44637 4029 44649 4032
rect 44683 4029 44695 4063
rect 44637 4023 44695 4029
rect 44726 4020 44732 4072
rect 44784 4060 44790 4072
rect 45373 4063 45431 4069
rect 45373 4060 45385 4063
rect 44784 4032 45385 4060
rect 44784 4020 44790 4032
rect 45373 4029 45385 4032
rect 45419 4029 45431 4063
rect 45373 4023 45431 4029
rect 45462 4020 45468 4072
rect 45520 4060 45526 4072
rect 46109 4063 46167 4069
rect 46109 4060 46121 4063
rect 45520 4032 46121 4060
rect 45520 4020 45526 4032
rect 46109 4029 46121 4032
rect 46155 4029 46167 4063
rect 46109 4023 46167 4029
rect 44358 3992 44364 4004
rect 43732 3964 44364 3992
rect 44358 3952 44364 3964
rect 44416 3952 44422 4004
rect 44818 3952 44824 4004
rect 44876 3992 44882 4004
rect 46676 3992 46704 4091
rect 48130 4088 48136 4140
rect 48188 4128 48194 4140
rect 48225 4131 48283 4137
rect 48225 4128 48237 4131
rect 48188 4100 48237 4128
rect 48188 4088 48194 4100
rect 48225 4097 48237 4100
rect 48271 4097 48283 4131
rect 48225 4091 48283 4097
rect 51718 4088 51724 4140
rect 51776 4128 51782 4140
rect 53929 4131 53987 4137
rect 53929 4128 53941 4131
rect 51776 4100 53941 4128
rect 51776 4088 51782 4100
rect 53929 4097 53941 4100
rect 53975 4097 53987 4131
rect 53929 4091 53987 4097
rect 54478 4088 54484 4140
rect 54536 4128 54542 4140
rect 54573 4131 54631 4137
rect 54573 4128 54585 4131
rect 54536 4100 54585 4128
rect 54536 4088 54542 4100
rect 54573 4097 54585 4100
rect 54619 4097 54631 4131
rect 58342 4128 58348 4140
rect 58303 4100 58348 4128
rect 54573 4091 54631 4097
rect 58342 4088 58348 4100
rect 58400 4088 58406 4140
rect 46842 4020 46848 4072
rect 46900 4060 46906 4072
rect 53466 4060 53472 4072
rect 46900 4032 53472 4060
rect 46900 4020 46906 4032
rect 53466 4020 53472 4032
rect 53524 4020 53530 4072
rect 48406 3992 48412 4004
rect 44876 3964 46704 3992
rect 48367 3964 48412 3992
rect 44876 3952 44882 3964
rect 48406 3952 48412 3964
rect 48464 3952 48470 4004
rect 53650 3952 53656 4004
rect 53708 3992 53714 4004
rect 54757 3995 54815 4001
rect 54757 3992 54769 3995
rect 53708 3964 54769 3992
rect 53708 3952 53714 3964
rect 54757 3961 54769 3964
rect 54803 3961 54815 3995
rect 54757 3955 54815 3961
rect 37884 3896 39620 3924
rect 37884 3884 37890 3896
rect 42518 3884 42524 3936
rect 42576 3924 42582 3936
rect 43622 3924 43628 3936
rect 42576 3896 43628 3924
rect 42576 3884 42582 3896
rect 43622 3884 43628 3896
rect 43680 3884 43686 3936
rect 43990 3884 43996 3936
rect 44048 3924 44054 3936
rect 45922 3924 45928 3936
rect 44048 3896 45928 3924
rect 44048 3884 44054 3896
rect 45922 3884 45928 3896
rect 45980 3884 45986 3936
rect 47026 3884 47032 3936
rect 47084 3924 47090 3936
rect 47302 3924 47308 3936
rect 47084 3896 47308 3924
rect 47084 3884 47090 3896
rect 47302 3884 47308 3896
rect 47360 3884 47366 3936
rect 47486 3884 47492 3936
rect 47544 3924 47550 3936
rect 52273 3927 52331 3933
rect 52273 3924 52285 3927
rect 47544 3896 52285 3924
rect 47544 3884 47550 3896
rect 52273 3893 52285 3896
rect 52319 3893 52331 3927
rect 52273 3887 52331 3893
rect 1104 3834 58880 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 58880 3834
rect 1104 3760 58880 3782
rect 5169 3723 5227 3729
rect 5169 3689 5181 3723
rect 5215 3720 5227 3723
rect 7006 3720 7012 3732
rect 5215 3692 7012 3720
rect 5215 3689 5227 3692
rect 5169 3683 5227 3689
rect 7006 3680 7012 3692
rect 7064 3680 7070 3732
rect 7466 3680 7472 3732
rect 7524 3720 7530 3732
rect 7524 3692 9168 3720
rect 7524 3680 7530 3692
rect 5994 3652 6000 3664
rect 5955 3624 6000 3652
rect 5994 3612 6000 3624
rect 6052 3612 6058 3664
rect 7558 3652 7564 3664
rect 7519 3624 7564 3652
rect 7558 3612 7564 3624
rect 7616 3612 7622 3664
rect 7650 3612 7656 3664
rect 7708 3652 7714 3664
rect 8389 3655 8447 3661
rect 7708 3624 7753 3652
rect 7708 3612 7714 3624
rect 8389 3621 8401 3655
rect 8435 3621 8447 3655
rect 8389 3615 8447 3621
rect 8573 3655 8631 3661
rect 8573 3621 8585 3655
rect 8619 3652 8631 3655
rect 8846 3652 8852 3664
rect 8619 3624 8852 3652
rect 8619 3621 8631 3624
rect 8573 3615 8631 3621
rect 6733 3587 6791 3593
rect 2746 3556 6316 3584
rect 1581 3519 1639 3525
rect 1581 3485 1593 3519
rect 1627 3516 1639 3519
rect 2746 3516 2774 3556
rect 1627 3488 2774 3516
rect 5077 3519 5135 3525
rect 1627 3485 1639 3488
rect 1581 3479 1639 3485
rect 5077 3485 5089 3519
rect 5123 3516 5135 3519
rect 6178 3516 6184 3528
rect 5123 3488 6184 3516
rect 5123 3485 5135 3488
rect 5077 3479 5135 3485
rect 6178 3476 6184 3488
rect 6236 3476 6242 3528
rect 6288 3516 6316 3556
rect 6733 3553 6745 3587
rect 6779 3584 6791 3587
rect 8404 3584 8432 3615
rect 8846 3612 8852 3624
rect 8904 3612 8910 3664
rect 9140 3652 9168 3692
rect 10594 3680 10600 3732
rect 10652 3720 10658 3732
rect 10873 3723 10931 3729
rect 10873 3720 10885 3723
rect 10652 3692 10885 3720
rect 10652 3680 10658 3692
rect 10873 3689 10885 3692
rect 10919 3689 10931 3723
rect 12805 3723 12863 3729
rect 10873 3683 10931 3689
rect 12452 3692 12756 3720
rect 10689 3655 10747 3661
rect 10689 3652 10701 3655
rect 9140 3624 10701 3652
rect 10689 3621 10701 3624
rect 10735 3621 10747 3655
rect 11882 3652 11888 3664
rect 11843 3624 11888 3652
rect 10689 3615 10747 3621
rect 11882 3612 11888 3624
rect 11940 3612 11946 3664
rect 6779 3556 8432 3584
rect 9401 3587 9459 3593
rect 6779 3553 6791 3556
rect 6733 3547 6791 3553
rect 9401 3553 9413 3587
rect 9447 3553 9459 3587
rect 9401 3547 9459 3553
rect 9677 3587 9735 3593
rect 9677 3553 9689 3587
rect 9723 3584 9735 3587
rect 12452 3584 12480 3692
rect 12618 3652 12624 3664
rect 12579 3624 12624 3652
rect 12618 3612 12624 3624
rect 12676 3612 12682 3664
rect 12728 3652 12756 3692
rect 12805 3689 12817 3723
rect 12851 3720 12863 3723
rect 12894 3720 12900 3732
rect 12851 3692 12900 3720
rect 12851 3689 12863 3692
rect 12805 3683 12863 3689
rect 12894 3680 12900 3692
rect 12952 3680 12958 3732
rect 13725 3723 13783 3729
rect 13725 3689 13737 3723
rect 13771 3720 13783 3723
rect 14642 3720 14648 3732
rect 13771 3692 14648 3720
rect 13771 3689 13783 3692
rect 13725 3683 13783 3689
rect 14642 3680 14648 3692
rect 14700 3680 14706 3732
rect 16117 3723 16175 3729
rect 16117 3689 16129 3723
rect 16163 3720 16175 3723
rect 17954 3720 17960 3732
rect 16163 3692 17960 3720
rect 16163 3689 16175 3692
rect 16117 3683 16175 3689
rect 17954 3680 17960 3692
rect 18012 3680 18018 3732
rect 18506 3680 18512 3732
rect 18564 3720 18570 3732
rect 19242 3720 19248 3732
rect 18564 3692 19248 3720
rect 18564 3680 18570 3692
rect 19242 3680 19248 3692
rect 19300 3680 19306 3732
rect 20346 3720 20352 3732
rect 19628 3692 20352 3720
rect 13538 3652 13544 3664
rect 12728 3624 13544 3652
rect 13538 3612 13544 3624
rect 13596 3612 13602 3664
rect 13633 3655 13691 3661
rect 13633 3621 13645 3655
rect 13679 3652 13691 3655
rect 13814 3652 13820 3664
rect 13679 3624 13820 3652
rect 13679 3621 13691 3624
rect 13633 3615 13691 3621
rect 13814 3612 13820 3624
rect 13872 3612 13878 3664
rect 15930 3652 15936 3664
rect 15891 3624 15936 3652
rect 15930 3612 15936 3624
rect 15988 3612 15994 3664
rect 19628 3652 19656 3692
rect 20346 3680 20352 3692
rect 20404 3680 20410 3732
rect 20714 3680 20720 3732
rect 20772 3720 20778 3732
rect 20772 3692 23704 3720
rect 20772 3680 20778 3692
rect 20990 3652 20996 3664
rect 17788 3624 19656 3652
rect 20951 3624 20996 3652
rect 9723 3556 12480 3584
rect 9723 3553 9735 3556
rect 9677 3547 9735 3553
rect 9416 3516 9444 3547
rect 12526 3544 12532 3596
rect 12584 3584 12590 3596
rect 17788 3593 17816 3624
rect 20990 3612 20996 3624
rect 21048 3612 21054 3664
rect 17773 3587 17831 3593
rect 12584 3556 17724 3584
rect 12584 3544 12590 3556
rect 9582 3516 9588 3528
rect 6288 3488 9444 3516
rect 9543 3488 9588 3516
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 9769 3519 9827 3525
rect 9769 3485 9781 3519
rect 9815 3485 9827 3519
rect 9769 3479 9827 3485
rect 1854 3448 1860 3460
rect 1815 3420 1860 3448
rect 1854 3408 1860 3420
rect 1912 3408 1918 3460
rect 5813 3451 5871 3457
rect 5813 3417 5825 3451
rect 5859 3448 5871 3451
rect 6549 3451 6607 3457
rect 5859 3420 6500 3448
rect 5859 3417 5871 3420
rect 5813 3411 5871 3417
rect 6472 3380 6500 3420
rect 6549 3417 6561 3451
rect 6595 3448 6607 3451
rect 7193 3451 7251 3457
rect 6595 3420 7144 3448
rect 6595 3417 6607 3420
rect 6549 3411 6607 3417
rect 7006 3380 7012 3392
rect 6472 3352 7012 3380
rect 7006 3340 7012 3352
rect 7064 3340 7070 3392
rect 7116 3380 7144 3420
rect 7193 3417 7205 3451
rect 7239 3448 7251 3451
rect 8113 3451 8171 3457
rect 8113 3448 8125 3451
rect 7239 3420 8125 3448
rect 7239 3417 7251 3420
rect 7193 3411 7251 3417
rect 8113 3417 8125 3420
rect 8159 3448 8171 3451
rect 8202 3448 8208 3460
rect 8159 3420 8208 3448
rect 8159 3417 8171 3420
rect 8113 3411 8171 3417
rect 8202 3408 8208 3420
rect 8260 3448 8266 3460
rect 8386 3448 8392 3460
rect 8260 3420 8392 3448
rect 8260 3408 8266 3420
rect 8386 3408 8392 3420
rect 8444 3408 8450 3460
rect 8478 3408 8484 3460
rect 8536 3448 8542 3460
rect 8846 3448 8852 3460
rect 8536 3420 8852 3448
rect 8536 3408 8542 3420
rect 8846 3408 8852 3420
rect 8904 3408 8910 3460
rect 9784 3448 9812 3479
rect 9858 3476 9864 3528
rect 9916 3516 9922 3528
rect 9916 3488 9961 3516
rect 9916 3476 9922 3488
rect 10318 3476 10324 3528
rect 10376 3516 10382 3528
rect 10413 3519 10471 3525
rect 10413 3516 10425 3519
rect 10376 3488 10425 3516
rect 10376 3476 10382 3488
rect 10413 3485 10425 3488
rect 10459 3485 10471 3519
rect 10413 3479 10471 3485
rect 11701 3519 11759 3525
rect 11701 3485 11713 3519
rect 11747 3516 11759 3519
rect 13354 3516 13360 3528
rect 11747 3488 13360 3516
rect 11747 3485 11759 3488
rect 11701 3479 11759 3485
rect 13354 3476 13360 3488
rect 13412 3476 13418 3528
rect 14737 3519 14795 3525
rect 14737 3485 14749 3519
rect 14783 3516 14795 3519
rect 15102 3516 15108 3528
rect 14783 3488 15108 3516
rect 14783 3485 14795 3488
rect 14737 3479 14795 3485
rect 15102 3476 15108 3488
rect 15160 3476 15166 3528
rect 15654 3516 15660 3528
rect 15615 3488 15660 3516
rect 15654 3476 15660 3488
rect 15712 3476 15718 3528
rect 17037 3519 17095 3525
rect 17037 3485 17049 3519
rect 17083 3516 17095 3519
rect 17218 3516 17224 3528
rect 17083 3488 17224 3516
rect 17083 3485 17095 3488
rect 17037 3479 17095 3485
rect 17218 3476 17224 3488
rect 17276 3476 17282 3528
rect 17494 3516 17500 3528
rect 17455 3488 17500 3516
rect 17494 3476 17500 3488
rect 17552 3476 17558 3528
rect 17696 3516 17724 3556
rect 17773 3553 17785 3587
rect 17819 3553 17831 3587
rect 18966 3584 18972 3596
rect 17773 3547 17831 3553
rect 18340 3556 18972 3584
rect 18340 3516 18368 3556
rect 18966 3544 18972 3556
rect 19024 3544 19030 3596
rect 19518 3584 19524 3596
rect 19352 3556 19524 3584
rect 17696 3488 18368 3516
rect 18414 3476 18420 3528
rect 18472 3516 18478 3528
rect 19352 3516 19380 3556
rect 19518 3544 19524 3556
rect 19576 3544 19582 3596
rect 21174 3544 21180 3596
rect 21232 3584 21238 3596
rect 22097 3587 22155 3593
rect 22097 3584 22109 3587
rect 21232 3556 22109 3584
rect 21232 3544 21238 3556
rect 22097 3553 22109 3556
rect 22143 3584 22155 3587
rect 22370 3584 22376 3596
rect 22143 3556 22376 3584
rect 22143 3553 22155 3556
rect 22097 3547 22155 3553
rect 22370 3544 22376 3556
rect 22428 3544 22434 3596
rect 18472 3488 18517 3516
rect 18616 3488 19380 3516
rect 19613 3519 19671 3525
rect 18472 3476 18478 3488
rect 9950 3448 9956 3460
rect 9784 3420 9956 3448
rect 9950 3408 9956 3420
rect 10008 3408 10014 3460
rect 12342 3448 12348 3460
rect 12255 3420 12348 3448
rect 12342 3408 12348 3420
rect 12400 3448 12406 3460
rect 13265 3451 13323 3457
rect 13265 3448 13277 3451
rect 12400 3420 13277 3448
rect 12400 3408 12406 3420
rect 13265 3417 13277 3420
rect 13311 3417 13323 3451
rect 14182 3448 14188 3460
rect 13265 3411 13323 3417
rect 13372 3420 14188 3448
rect 8570 3380 8576 3392
rect 7116 3352 8576 3380
rect 8570 3340 8576 3352
rect 8628 3340 8634 3392
rect 9214 3340 9220 3392
rect 9272 3380 9278 3392
rect 12526 3380 12532 3392
rect 9272 3352 12532 3380
rect 9272 3340 9278 3352
rect 12526 3340 12532 3352
rect 12584 3340 12590 3392
rect 12802 3340 12808 3392
rect 12860 3380 12866 3392
rect 13372 3380 13400 3420
rect 14182 3408 14188 3420
rect 14240 3408 14246 3460
rect 15013 3451 15071 3457
rect 15013 3417 15025 3451
rect 15059 3448 15071 3451
rect 15562 3448 15568 3460
rect 15059 3420 15568 3448
rect 15059 3417 15071 3420
rect 15013 3411 15071 3417
rect 15562 3408 15568 3420
rect 15620 3408 15626 3460
rect 16574 3408 16580 3460
rect 16632 3448 16638 3460
rect 17770 3448 17776 3460
rect 16632 3420 17776 3448
rect 16632 3408 16638 3420
rect 17770 3408 17776 3420
rect 17828 3408 17834 3460
rect 12860 3352 13400 3380
rect 12860 3340 12866 3352
rect 13538 3340 13544 3392
rect 13596 3380 13602 3392
rect 18616 3380 18644 3488
rect 19613 3485 19625 3519
rect 19659 3516 19671 3519
rect 22649 3519 22707 3525
rect 22649 3516 22661 3519
rect 19659 3488 22661 3516
rect 19659 3485 19671 3488
rect 19613 3479 19671 3485
rect 20088 3460 20116 3488
rect 22649 3485 22661 3488
rect 22695 3516 22707 3519
rect 23290 3516 23296 3528
rect 22695 3488 23296 3516
rect 22695 3485 22707 3488
rect 22649 3479 22707 3485
rect 23290 3476 23296 3488
rect 23348 3476 23354 3528
rect 23676 3516 23704 3692
rect 23750 3680 23756 3732
rect 23808 3720 23814 3732
rect 24581 3723 24639 3729
rect 24581 3720 24593 3723
rect 23808 3692 24593 3720
rect 23808 3680 23814 3692
rect 24581 3689 24593 3692
rect 24627 3689 24639 3723
rect 27706 3720 27712 3732
rect 27667 3692 27712 3720
rect 24581 3683 24639 3689
rect 27706 3680 27712 3692
rect 27764 3680 27770 3732
rect 33686 3720 33692 3732
rect 27816 3692 33272 3720
rect 33647 3692 33692 3720
rect 27816 3652 27844 3692
rect 25056 3624 27844 3652
rect 25056 3593 25084 3624
rect 28258 3612 28264 3664
rect 28316 3652 28322 3664
rect 29730 3652 29736 3664
rect 28316 3624 29736 3652
rect 28316 3612 28322 3624
rect 29730 3612 29736 3624
rect 29788 3612 29794 3664
rect 33244 3652 33272 3692
rect 33686 3680 33692 3692
rect 33744 3680 33750 3732
rect 37182 3680 37188 3732
rect 37240 3720 37246 3732
rect 39666 3720 39672 3732
rect 37240 3692 39672 3720
rect 37240 3680 37246 3692
rect 39666 3680 39672 3692
rect 39724 3680 39730 3732
rect 42426 3680 42432 3732
rect 42484 3720 42490 3732
rect 42889 3723 42947 3729
rect 42889 3720 42901 3723
rect 42484 3692 42901 3720
rect 42484 3680 42490 3692
rect 42889 3689 42901 3692
rect 42935 3689 42947 3723
rect 42889 3683 42947 3689
rect 43714 3680 43720 3732
rect 43772 3720 43778 3732
rect 44174 3720 44180 3732
rect 43772 3692 44180 3720
rect 43772 3680 43778 3692
rect 44174 3680 44180 3692
rect 44232 3680 44238 3732
rect 44358 3680 44364 3732
rect 44416 3720 44422 3732
rect 46109 3723 46167 3729
rect 46109 3720 46121 3723
rect 44416 3692 46121 3720
rect 44416 3680 44422 3692
rect 46109 3689 46121 3692
rect 46155 3689 46167 3723
rect 47026 3720 47032 3732
rect 46987 3692 47032 3720
rect 46109 3683 46167 3689
rect 47026 3680 47032 3692
rect 47084 3680 47090 3732
rect 47854 3680 47860 3732
rect 47912 3720 47918 3732
rect 47949 3723 48007 3729
rect 47949 3720 47961 3723
rect 47912 3692 47961 3720
rect 47912 3680 47918 3692
rect 47949 3689 47961 3692
rect 47995 3689 48007 3723
rect 47949 3683 48007 3689
rect 48590 3680 48596 3732
rect 48648 3720 48654 3732
rect 48685 3723 48743 3729
rect 48685 3720 48697 3723
rect 48648 3692 48697 3720
rect 48648 3680 48654 3692
rect 48685 3689 48697 3692
rect 48731 3689 48743 3723
rect 49418 3720 49424 3732
rect 49379 3692 49424 3720
rect 48685 3683 48743 3689
rect 49418 3680 49424 3692
rect 49476 3680 49482 3732
rect 52454 3680 52460 3732
rect 52512 3720 52518 3732
rect 53469 3723 53527 3729
rect 53469 3720 53481 3723
rect 52512 3692 53481 3720
rect 52512 3680 52518 3692
rect 53469 3689 53481 3692
rect 53515 3689 53527 3723
rect 54202 3720 54208 3732
rect 54163 3692 54208 3720
rect 53469 3683 53527 3689
rect 54202 3680 54208 3692
rect 54260 3680 54266 3732
rect 55030 3680 55036 3732
rect 55088 3720 55094 3732
rect 55677 3723 55735 3729
rect 55677 3720 55689 3723
rect 55088 3692 55689 3720
rect 55088 3680 55094 3692
rect 55677 3689 55689 3692
rect 55723 3689 55735 3723
rect 55677 3683 55735 3689
rect 33244 3624 37228 3652
rect 25041 3587 25099 3593
rect 25041 3553 25053 3587
rect 25087 3553 25099 3587
rect 25041 3547 25099 3553
rect 25225 3587 25283 3593
rect 25225 3553 25237 3587
rect 25271 3584 25283 3587
rect 27430 3584 27436 3596
rect 25271 3556 26832 3584
rect 25271 3553 25283 3556
rect 25225 3547 25283 3553
rect 24949 3519 25007 3525
rect 24949 3516 24961 3519
rect 23676 3488 24961 3516
rect 24949 3485 24961 3488
rect 24995 3485 25007 3519
rect 24949 3479 25007 3485
rect 25777 3519 25835 3525
rect 25777 3485 25789 3519
rect 25823 3516 25835 3519
rect 26510 3516 26516 3528
rect 25823 3488 26516 3516
rect 25823 3485 25835 3488
rect 25777 3479 25835 3485
rect 26510 3476 26516 3488
rect 26568 3476 26574 3528
rect 18693 3451 18751 3457
rect 18693 3417 18705 3451
rect 18739 3417 18751 3451
rect 18693 3411 18751 3417
rect 13596 3352 18644 3380
rect 18708 3380 18736 3411
rect 18782 3408 18788 3460
rect 18840 3448 18846 3460
rect 19869 3451 19927 3457
rect 18840 3420 19656 3448
rect 18840 3408 18846 3420
rect 19518 3380 19524 3392
rect 18708 3352 19524 3380
rect 13596 3340 13602 3352
rect 19518 3340 19524 3352
rect 19576 3340 19582 3392
rect 19628 3380 19656 3420
rect 19869 3417 19881 3451
rect 19915 3417 19927 3451
rect 19869 3411 19927 3417
rect 19884 3380 19912 3411
rect 19978 3408 19984 3460
rect 20036 3408 20042 3460
rect 20070 3408 20076 3460
rect 20128 3408 20134 3460
rect 20898 3408 20904 3460
rect 20956 3448 20962 3460
rect 21818 3448 21824 3460
rect 20956 3420 21588 3448
rect 21779 3420 21824 3448
rect 20956 3408 20962 3420
rect 19628 3352 19912 3380
rect 19996 3380 20024 3408
rect 21082 3380 21088 3392
rect 19996 3352 21088 3380
rect 21082 3340 21088 3352
rect 21140 3340 21146 3392
rect 21450 3380 21456 3392
rect 21411 3352 21456 3380
rect 21450 3340 21456 3352
rect 21508 3340 21514 3392
rect 21560 3380 21588 3420
rect 21818 3408 21824 3420
rect 21876 3408 21882 3460
rect 22916 3451 22974 3457
rect 22916 3417 22928 3451
rect 22962 3448 22974 3451
rect 23198 3448 23204 3460
rect 22962 3420 23204 3448
rect 22962 3417 22974 3420
rect 22916 3411 22974 3417
rect 23198 3408 23204 3420
rect 23256 3408 23262 3460
rect 24118 3408 24124 3460
rect 24176 3448 24182 3460
rect 26053 3451 26111 3457
rect 26053 3448 26065 3451
rect 24176 3420 26065 3448
rect 24176 3408 24182 3420
rect 26053 3417 26065 3420
rect 26099 3417 26111 3451
rect 26694 3448 26700 3460
rect 26655 3420 26700 3448
rect 26053 3411 26111 3417
rect 26694 3408 26700 3420
rect 26752 3408 26758 3460
rect 26804 3448 26832 3556
rect 26896 3556 27436 3584
rect 26896 3525 26924 3556
rect 27430 3544 27436 3556
rect 27488 3544 27494 3596
rect 28353 3587 28411 3593
rect 28353 3553 28365 3587
rect 28399 3584 28411 3587
rect 29362 3584 29368 3596
rect 28399 3556 29368 3584
rect 28399 3553 28411 3556
rect 28353 3547 28411 3553
rect 29362 3544 29368 3556
rect 29420 3544 29426 3596
rect 30098 3544 30104 3596
rect 30156 3584 30162 3596
rect 32214 3584 32220 3596
rect 30156 3556 32220 3584
rect 30156 3544 30162 3556
rect 32214 3544 32220 3556
rect 32272 3584 32278 3596
rect 32309 3587 32367 3593
rect 32309 3584 32321 3587
rect 32272 3556 32321 3584
rect 32272 3544 32278 3556
rect 32309 3553 32321 3556
rect 32355 3553 32367 3587
rect 32585 3587 32643 3593
rect 32585 3584 32597 3587
rect 32309 3547 32367 3553
rect 32416 3556 32597 3584
rect 26881 3519 26939 3525
rect 26881 3485 26893 3519
rect 26927 3485 26939 3519
rect 26881 3479 26939 3485
rect 26993 3519 27051 3525
rect 26993 3485 27005 3519
rect 27039 3516 27051 3519
rect 28718 3516 28724 3528
rect 27039 3488 28724 3516
rect 27039 3485 27051 3488
rect 26993 3479 27051 3485
rect 28718 3476 28724 3488
rect 28776 3476 28782 3528
rect 29086 3516 29092 3528
rect 28828 3488 29092 3516
rect 27083 3451 27141 3457
rect 27083 3448 27095 3451
rect 26804 3420 27095 3448
rect 26896 3392 26924 3420
rect 27083 3417 27095 3420
rect 27129 3417 27141 3451
rect 27246 3448 27252 3460
rect 27207 3420 27252 3448
rect 27083 3411 27141 3417
rect 27246 3408 27252 3420
rect 27304 3408 27310 3460
rect 27338 3408 27344 3460
rect 27396 3448 27402 3460
rect 28169 3451 28227 3457
rect 28169 3448 28181 3451
rect 27396 3420 28181 3448
rect 27396 3408 27402 3420
rect 28169 3417 28181 3420
rect 28215 3448 28227 3451
rect 28828 3448 28856 3488
rect 29086 3476 29092 3488
rect 29144 3476 29150 3528
rect 29181 3519 29239 3525
rect 29181 3485 29193 3519
rect 29227 3516 29239 3519
rect 30285 3519 30343 3525
rect 30285 3516 30297 3519
rect 29227 3488 30297 3516
rect 29227 3485 29239 3488
rect 29181 3479 29239 3485
rect 30285 3485 30297 3488
rect 30331 3485 30343 3519
rect 31570 3516 31576 3528
rect 31531 3488 31576 3516
rect 30285 3479 30343 3485
rect 31570 3476 31576 3488
rect 31628 3476 31634 3528
rect 31665 3519 31723 3525
rect 31665 3485 31677 3519
rect 31711 3516 31723 3519
rect 32030 3516 32036 3528
rect 31711 3488 32036 3516
rect 31711 3485 31723 3488
rect 31665 3479 31723 3485
rect 32030 3476 32036 3488
rect 32088 3476 32094 3528
rect 28215 3420 28856 3448
rect 28997 3451 29055 3457
rect 28215 3417 28227 3420
rect 28169 3411 28227 3417
rect 28997 3417 29009 3451
rect 29043 3448 29055 3451
rect 29270 3448 29276 3460
rect 29043 3420 29276 3448
rect 29043 3417 29055 3420
rect 28997 3411 29055 3417
rect 29270 3408 29276 3420
rect 29328 3408 29334 3460
rect 30190 3408 30196 3460
rect 30248 3448 30254 3460
rect 30561 3451 30619 3457
rect 30561 3448 30573 3451
rect 30248 3420 30573 3448
rect 30248 3408 30254 3420
rect 30561 3417 30573 3420
rect 30607 3417 30619 3451
rect 30561 3411 30619 3417
rect 31849 3451 31907 3457
rect 31849 3417 31861 3451
rect 31895 3448 31907 3451
rect 32416 3448 32444 3556
rect 32585 3553 32597 3556
rect 32631 3553 32643 3587
rect 32585 3547 32643 3553
rect 33226 3544 33232 3596
rect 33284 3584 33290 3596
rect 35069 3587 35127 3593
rect 35069 3584 35081 3587
rect 33284 3556 35081 3584
rect 33284 3544 33290 3556
rect 35069 3553 35081 3556
rect 35115 3553 35127 3587
rect 35069 3547 35127 3553
rect 36078 3544 36084 3596
rect 36136 3584 36142 3596
rect 36814 3584 36820 3596
rect 36136 3556 36820 3584
rect 36136 3544 36142 3556
rect 36814 3544 36820 3556
rect 36872 3544 36878 3596
rect 32858 3476 32864 3528
rect 32916 3516 32922 3528
rect 33318 3516 33324 3528
rect 32916 3488 33324 3516
rect 32916 3476 32922 3488
rect 33318 3476 33324 3488
rect 33376 3476 33382 3528
rect 33410 3476 33416 3528
rect 33468 3516 33474 3528
rect 33962 3516 33968 3528
rect 33468 3488 33968 3516
rect 33468 3476 33474 3488
rect 33962 3476 33968 3488
rect 34020 3476 34026 3528
rect 34698 3476 34704 3528
rect 34756 3516 34762 3528
rect 34885 3519 34943 3525
rect 34885 3516 34897 3519
rect 34756 3488 34897 3516
rect 34756 3476 34762 3488
rect 34885 3485 34897 3488
rect 34931 3485 34943 3519
rect 36170 3516 36176 3528
rect 36131 3488 36176 3516
rect 34885 3479 34943 3485
rect 36170 3476 36176 3488
rect 36228 3476 36234 3528
rect 37200 3516 37228 3624
rect 38286 3612 38292 3664
rect 38344 3652 38350 3664
rect 38657 3655 38715 3661
rect 38657 3652 38669 3655
rect 38344 3624 38669 3652
rect 38344 3612 38350 3624
rect 38657 3621 38669 3624
rect 38703 3621 38715 3655
rect 38657 3615 38715 3621
rect 40770 3612 40776 3664
rect 40828 3652 40834 3664
rect 41966 3652 41972 3664
rect 40828 3624 41092 3652
rect 41927 3624 41972 3652
rect 40828 3612 40834 3624
rect 37277 3587 37335 3593
rect 37277 3553 37289 3587
rect 37323 3584 37335 3587
rect 39114 3584 39120 3596
rect 37323 3556 39120 3584
rect 37323 3553 37335 3556
rect 37277 3547 37335 3553
rect 39114 3544 39120 3556
rect 39172 3544 39178 3596
rect 40126 3584 40132 3596
rect 40087 3556 40132 3584
rect 40126 3544 40132 3556
rect 40184 3544 40190 3596
rect 40862 3584 40868 3596
rect 40823 3556 40868 3584
rect 40862 3544 40868 3556
rect 40920 3544 40926 3596
rect 41064 3593 41092 3624
rect 41966 3612 41972 3624
rect 42024 3612 42030 3664
rect 42702 3612 42708 3664
rect 42760 3652 42766 3664
rect 42760 3624 44772 3652
rect 42760 3612 42766 3624
rect 41049 3587 41107 3593
rect 41049 3553 41061 3587
rect 41095 3553 41107 3587
rect 41049 3547 41107 3553
rect 43346 3544 43352 3596
rect 43404 3544 43410 3596
rect 43806 3544 43812 3596
rect 43864 3544 43870 3596
rect 44082 3584 44088 3596
rect 44013 3556 44088 3584
rect 37366 3516 37372 3528
rect 37200 3488 37372 3516
rect 37366 3476 37372 3488
rect 37424 3476 37430 3528
rect 37550 3516 37556 3528
rect 37511 3488 37556 3516
rect 37550 3476 37556 3488
rect 37608 3476 37614 3528
rect 40773 3519 40831 3525
rect 40773 3516 40785 3519
rect 38212 3488 40785 3516
rect 34330 3448 34336 3460
rect 31895 3420 32444 3448
rect 33244 3420 34336 3448
rect 31895 3417 31907 3420
rect 31849 3411 31907 3417
rect 21913 3383 21971 3389
rect 21913 3380 21925 3383
rect 21560 3352 21925 3380
rect 21913 3349 21925 3352
rect 21959 3349 21971 3383
rect 21913 3343 21971 3349
rect 23658 3340 23664 3392
rect 23716 3380 23722 3392
rect 24029 3383 24087 3389
rect 24029 3380 24041 3383
rect 23716 3352 24041 3380
rect 23716 3340 23722 3352
rect 24029 3349 24041 3352
rect 24075 3349 24087 3383
rect 24029 3343 24087 3349
rect 26878 3340 26884 3392
rect 26936 3340 26942 3392
rect 28074 3380 28080 3392
rect 28035 3352 28080 3380
rect 28074 3340 28080 3352
rect 28132 3340 28138 3392
rect 28442 3340 28448 3392
rect 28500 3380 28506 3392
rect 32858 3380 32864 3392
rect 28500 3352 32864 3380
rect 28500 3340 28506 3352
rect 32858 3340 32864 3352
rect 32916 3340 32922 3392
rect 32950 3340 32956 3392
rect 33008 3380 33014 3392
rect 33244 3380 33272 3420
rect 34330 3408 34336 3420
rect 34388 3408 34394 3460
rect 34606 3408 34612 3460
rect 34664 3448 34670 3460
rect 35710 3448 35716 3460
rect 34664 3420 35716 3448
rect 34664 3408 34670 3420
rect 35710 3408 35716 3420
rect 35768 3408 35774 3460
rect 36725 3451 36783 3457
rect 36725 3417 36737 3451
rect 36771 3417 36783 3451
rect 36725 3411 36783 3417
rect 33008 3352 33272 3380
rect 33008 3340 33014 3352
rect 33318 3340 33324 3392
rect 33376 3380 33382 3392
rect 33870 3380 33876 3392
rect 33376 3352 33876 3380
rect 33376 3340 33382 3352
rect 33870 3340 33876 3352
rect 33928 3340 33934 3392
rect 34054 3340 34060 3392
rect 34112 3380 34118 3392
rect 35434 3380 35440 3392
rect 34112 3352 35440 3380
rect 34112 3340 34118 3352
rect 35434 3340 35440 3352
rect 35492 3340 35498 3392
rect 36538 3340 36544 3392
rect 36596 3380 36602 3392
rect 36740 3380 36768 3411
rect 38212 3380 38240 3488
rect 40773 3485 40785 3488
rect 40819 3516 40831 3519
rect 40954 3516 40960 3528
rect 40819 3488 40960 3516
rect 40819 3485 40831 3488
rect 40773 3479 40831 3485
rect 40954 3476 40960 3488
rect 41012 3476 41018 3528
rect 41138 3516 41144 3528
rect 41099 3488 41144 3516
rect 41138 3476 41144 3488
rect 41196 3476 41202 3528
rect 41785 3519 41843 3525
rect 41785 3485 41797 3519
rect 41831 3485 41843 3519
rect 41785 3479 41843 3485
rect 38286 3408 38292 3460
rect 38344 3448 38350 3460
rect 41800 3448 41828 3479
rect 42518 3476 42524 3528
rect 42576 3516 42582 3528
rect 43245 3519 43303 3525
rect 43245 3516 43257 3519
rect 42576 3488 43257 3516
rect 42576 3476 42582 3488
rect 43245 3485 43257 3488
rect 43291 3485 43303 3519
rect 43364 3516 43392 3544
rect 43533 3519 43591 3525
rect 43364 3514 43484 3516
rect 43533 3514 43545 3519
rect 43364 3488 43545 3514
rect 43456 3486 43545 3488
rect 43245 3479 43303 3485
rect 43533 3485 43545 3486
rect 43579 3485 43591 3519
rect 43646 3519 43704 3525
rect 43646 3516 43658 3519
rect 43640 3486 43658 3516
rect 43533 3479 43591 3485
rect 43646 3485 43658 3486
rect 43692 3514 43704 3519
rect 43824 3516 43852 3544
rect 43732 3514 43852 3516
rect 43692 3488 43852 3514
rect 43901 3519 43959 3525
rect 43692 3486 43760 3488
rect 43692 3485 43704 3486
rect 43646 3479 43704 3485
rect 43901 3485 43913 3519
rect 43947 3514 43959 3519
rect 44013 3514 44041 3556
rect 44082 3544 44088 3556
rect 44140 3544 44146 3596
rect 44744 3584 44772 3624
rect 45094 3612 45100 3664
rect 45152 3652 45158 3664
rect 46014 3652 46020 3664
rect 45152 3624 46020 3652
rect 45152 3612 45158 3624
rect 46014 3612 46020 3624
rect 46072 3612 46078 3664
rect 47394 3612 47400 3664
rect 47452 3652 47458 3664
rect 50617 3655 50675 3661
rect 50617 3652 50629 3655
rect 47452 3624 50629 3652
rect 47452 3612 47458 3624
rect 50617 3621 50629 3624
rect 50663 3621 50675 3655
rect 50617 3615 50675 3621
rect 44744 3556 45324 3584
rect 44174 3516 44180 3528
rect 43947 3486 44041 3514
rect 44135 3488 44180 3516
rect 43947 3485 43959 3486
rect 43901 3479 43959 3485
rect 44174 3476 44180 3488
rect 44232 3476 44238 3528
rect 45296 3525 45324 3556
rect 46842 3544 46848 3596
rect 46900 3584 46906 3596
rect 51353 3587 51411 3593
rect 51353 3584 51365 3587
rect 46900 3556 51365 3584
rect 46900 3544 46906 3556
rect 51353 3553 51365 3556
rect 51399 3553 51411 3587
rect 52825 3587 52883 3593
rect 52825 3584 52837 3587
rect 51353 3547 51411 3553
rect 51460 3556 52837 3584
rect 45281 3519 45339 3525
rect 45281 3485 45293 3519
rect 45327 3485 45339 3519
rect 45281 3479 45339 3485
rect 47578 3476 47584 3528
rect 47636 3516 47642 3528
rect 48501 3519 48559 3525
rect 48501 3516 48513 3519
rect 47636 3488 48513 3516
rect 47636 3476 47642 3488
rect 48501 3485 48513 3488
rect 48547 3485 48559 3519
rect 48501 3479 48559 3485
rect 48774 3476 48780 3528
rect 48832 3516 48838 3528
rect 49237 3519 49295 3525
rect 49237 3516 49249 3519
rect 48832 3488 49249 3516
rect 48832 3476 48838 3488
rect 49237 3485 49249 3488
rect 49283 3485 49295 3519
rect 49237 3479 49295 3485
rect 49326 3476 49332 3528
rect 49384 3516 49390 3528
rect 51460 3516 51488 3556
rect 52825 3553 52837 3556
rect 52871 3553 52883 3587
rect 56870 3584 56876 3596
rect 56831 3556 56876 3584
rect 52825 3547 52883 3553
rect 56870 3544 56876 3556
rect 56928 3544 56934 3596
rect 49384 3488 51488 3516
rect 49384 3476 49390 3488
rect 51718 3476 51724 3528
rect 51776 3516 51782 3528
rect 52641 3519 52699 3525
rect 52641 3516 52653 3519
rect 51776 3488 52653 3516
rect 51776 3476 51782 3488
rect 52641 3485 52653 3488
rect 52687 3485 52699 3519
rect 52641 3479 52699 3485
rect 53190 3476 53196 3528
rect 53248 3516 53254 3528
rect 54113 3519 54171 3525
rect 54113 3516 54125 3519
rect 53248 3488 54125 3516
rect 53248 3476 53254 3488
rect 54113 3485 54125 3488
rect 54159 3485 54171 3519
rect 54113 3479 54171 3485
rect 54754 3476 54760 3528
rect 54812 3516 54818 3528
rect 55493 3519 55551 3525
rect 55493 3516 55505 3519
rect 54812 3488 55505 3516
rect 54812 3476 54818 3488
rect 55493 3485 55505 3488
rect 55539 3485 55551 3519
rect 55493 3479 55551 3485
rect 46017 3451 46075 3457
rect 46017 3448 46029 3451
rect 38344 3420 41828 3448
rect 43548 3420 46029 3448
rect 38344 3408 38350 3420
rect 36596 3352 38240 3380
rect 36596 3340 36602 3352
rect 38562 3340 38568 3392
rect 38620 3380 38626 3392
rect 40586 3380 40592 3392
rect 38620 3352 40592 3380
rect 38620 3340 38626 3352
rect 40586 3340 40592 3352
rect 40644 3340 40650 3392
rect 43254 3340 43260 3392
rect 43312 3380 43318 3392
rect 43548 3380 43576 3420
rect 46017 3417 46029 3420
rect 46063 3417 46075 3451
rect 46017 3411 46075 3417
rect 46750 3408 46756 3460
rect 46808 3448 46814 3460
rect 46937 3451 46995 3457
rect 46937 3448 46949 3451
rect 46808 3420 46949 3448
rect 46808 3408 46814 3420
rect 46937 3417 46949 3420
rect 46983 3417 46995 3451
rect 46937 3411 46995 3417
rect 47857 3451 47915 3457
rect 47857 3417 47869 3451
rect 47903 3417 47915 3451
rect 47857 3411 47915 3417
rect 43312 3352 43576 3380
rect 43312 3340 43318 3352
rect 43622 3340 43628 3392
rect 43680 3380 43686 3392
rect 45373 3383 45431 3389
rect 45373 3380 45385 3383
rect 43680 3352 45385 3380
rect 43680 3340 43686 3352
rect 45373 3349 45385 3352
rect 45419 3349 45431 3383
rect 45373 3343 45431 3349
rect 45462 3340 45468 3392
rect 45520 3380 45526 3392
rect 47872 3380 47900 3411
rect 49878 3408 49884 3460
rect 49936 3448 49942 3460
rect 50433 3451 50491 3457
rect 50433 3448 50445 3451
rect 49936 3420 50445 3448
rect 49936 3408 49942 3420
rect 50433 3417 50445 3420
rect 50479 3417 50491 3451
rect 50433 3411 50491 3417
rect 50614 3408 50620 3460
rect 50672 3448 50678 3460
rect 51169 3451 51227 3457
rect 51169 3448 51181 3451
rect 50672 3420 51181 3448
rect 50672 3408 50678 3420
rect 51169 3417 51181 3420
rect 51215 3417 51227 3451
rect 51169 3411 51227 3417
rect 51258 3408 51264 3460
rect 51316 3448 51322 3460
rect 51905 3451 51963 3457
rect 51905 3448 51917 3451
rect 51316 3420 51917 3448
rect 51316 3408 51322 3420
rect 51905 3417 51917 3420
rect 51951 3417 51963 3451
rect 51905 3411 51963 3417
rect 52270 3408 52276 3460
rect 52328 3448 52334 3460
rect 53377 3451 53435 3457
rect 53377 3448 53389 3451
rect 52328 3420 53389 3448
rect 52328 3408 52334 3420
rect 53377 3417 53389 3420
rect 53423 3417 53435 3451
rect 53377 3411 53435 3417
rect 53558 3408 53564 3460
rect 53616 3448 53622 3460
rect 57118 3451 57176 3457
rect 57118 3448 57130 3451
rect 53616 3420 57130 3448
rect 53616 3408 53622 3420
rect 57118 3417 57130 3420
rect 57164 3417 57176 3451
rect 57118 3411 57176 3417
rect 45520 3352 47900 3380
rect 45520 3340 45526 3352
rect 50798 3340 50804 3392
rect 50856 3380 50862 3392
rect 51997 3383 52055 3389
rect 51997 3380 52009 3383
rect 50856 3352 52009 3380
rect 50856 3340 50862 3352
rect 51997 3349 52009 3352
rect 52043 3349 52055 3383
rect 51997 3343 52055 3349
rect 57238 3340 57244 3392
rect 57296 3380 57302 3392
rect 58253 3383 58311 3389
rect 58253 3380 58265 3383
rect 57296 3352 58265 3380
rect 57296 3340 57302 3352
rect 58253 3349 58265 3352
rect 58299 3349 58311 3383
rect 58253 3343 58311 3349
rect 1104 3290 58880 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 58880 3290
rect 1104 3216 58880 3238
rect 8018 3176 8024 3188
rect 2746 3148 8024 3176
rect 1581 3043 1639 3049
rect 1581 3009 1593 3043
rect 1627 3040 1639 3043
rect 2746 3040 2774 3148
rect 8018 3136 8024 3148
rect 8076 3136 8082 3188
rect 8941 3179 8999 3185
rect 8941 3145 8953 3179
rect 8987 3176 8999 3179
rect 9858 3176 9864 3188
rect 8987 3148 9864 3176
rect 8987 3145 8999 3148
rect 8941 3139 8999 3145
rect 9858 3136 9864 3148
rect 9916 3136 9922 3188
rect 10873 3179 10931 3185
rect 10873 3145 10885 3179
rect 10919 3176 10931 3179
rect 12894 3176 12900 3188
rect 10919 3148 12900 3176
rect 10919 3145 10931 3148
rect 10873 3139 10931 3145
rect 12894 3136 12900 3148
rect 12952 3136 12958 3188
rect 12989 3179 13047 3185
rect 12989 3145 13001 3179
rect 13035 3176 13047 3179
rect 15930 3176 15936 3188
rect 13035 3148 15936 3176
rect 13035 3145 13047 3148
rect 12989 3139 13047 3145
rect 15930 3136 15936 3148
rect 15988 3136 15994 3188
rect 23198 3176 23204 3188
rect 16040 3148 23060 3176
rect 23159 3148 23204 3176
rect 4341 3111 4399 3117
rect 4341 3077 4353 3111
rect 4387 3108 4399 3111
rect 5902 3108 5908 3120
rect 4387 3080 5908 3108
rect 4387 3077 4399 3080
rect 4341 3071 4399 3077
rect 5902 3068 5908 3080
rect 5960 3068 5966 3120
rect 9122 3108 9128 3120
rect 7024 3080 9128 3108
rect 1627 3012 2774 3040
rect 4525 3043 4583 3049
rect 1627 3009 1639 3012
rect 1581 3003 1639 3009
rect 4525 3009 4537 3043
rect 4571 3040 4583 3043
rect 4614 3040 4620 3052
rect 4571 3012 4620 3040
rect 4571 3009 4583 3012
rect 4525 3003 4583 3009
rect 4614 3000 4620 3012
rect 4672 3000 4678 3052
rect 5077 3043 5135 3049
rect 5077 3009 5089 3043
rect 5123 3009 5135 3043
rect 5077 3003 5135 3009
rect 5813 3043 5871 3049
rect 5813 3009 5825 3043
rect 5859 3040 5871 3043
rect 7024 3040 7052 3080
rect 9122 3068 9128 3080
rect 9180 3068 9186 3120
rect 9784 3080 10272 3108
rect 5859 3012 7052 3040
rect 7101 3043 7159 3049
rect 5859 3009 5871 3012
rect 5813 3003 5871 3009
rect 7101 3009 7113 3043
rect 7147 3040 7159 3043
rect 7837 3043 7895 3049
rect 7147 3012 7788 3040
rect 7147 3009 7159 3012
rect 7101 3003 7159 3009
rect 1762 2972 1768 2984
rect 1723 2944 1768 2972
rect 1762 2932 1768 2944
rect 1820 2932 1826 2984
rect 5092 2972 5120 3003
rect 7558 2972 7564 2984
rect 5092 2944 7564 2972
rect 7558 2932 7564 2944
rect 7616 2932 7622 2984
rect 7760 2972 7788 3012
rect 7837 3009 7849 3043
rect 7883 3040 7895 3043
rect 9214 3040 9220 3052
rect 7883 3012 9220 3040
rect 7883 3009 7895 3012
rect 7837 3003 7895 3009
rect 9214 3000 9220 3012
rect 9272 3000 9278 3052
rect 9582 3040 9588 3052
rect 9543 3012 9588 3040
rect 9582 3000 9588 3012
rect 9640 3000 9646 3052
rect 9677 3043 9735 3049
rect 9677 3009 9689 3043
rect 9723 3040 9735 3043
rect 9784 3040 9812 3080
rect 9723 3012 9812 3040
rect 9861 3043 9919 3049
rect 9723 3009 9735 3012
rect 9677 3003 9735 3009
rect 9861 3009 9873 3043
rect 9907 3040 9919 3043
rect 10042 3040 10048 3052
rect 9907 3012 10048 3040
rect 9907 3009 9919 3012
rect 9861 3003 9919 3009
rect 10042 3000 10048 3012
rect 10100 3000 10106 3052
rect 10244 3040 10272 3080
rect 10318 3068 10324 3120
rect 10376 3108 10382 3120
rect 10413 3111 10471 3117
rect 10413 3108 10425 3111
rect 10376 3080 10425 3108
rect 10376 3068 10382 3080
rect 10413 3077 10425 3080
rect 10459 3077 10471 3111
rect 16040 3108 16068 3148
rect 18138 3108 18144 3120
rect 10413 3071 10471 3077
rect 12084 3080 16068 3108
rect 17696 3080 18144 3108
rect 12084 3040 12112 3080
rect 10244 3012 12112 3040
rect 12161 3043 12219 3049
rect 12161 3009 12173 3043
rect 12207 3040 12219 3043
rect 12802 3040 12808 3052
rect 12207 3012 12808 3040
rect 12207 3009 12219 3012
rect 12161 3003 12219 3009
rect 12802 3000 12808 3012
rect 12860 3000 12866 3052
rect 12897 3043 12955 3049
rect 12897 3009 12909 3043
rect 12943 3009 12955 3043
rect 12897 3003 12955 3009
rect 13541 3043 13599 3049
rect 13541 3009 13553 3043
rect 13587 3040 13599 3043
rect 13630 3040 13636 3052
rect 13587 3012 13636 3040
rect 13587 3009 13599 3012
rect 13541 3003 13599 3009
rect 8202 2972 8208 2984
rect 7760 2944 8208 2972
rect 8202 2932 8208 2944
rect 8260 2932 8266 2984
rect 8386 2932 8392 2984
rect 8444 2972 8450 2984
rect 8481 2975 8539 2981
rect 8481 2972 8493 2975
rect 8444 2944 8493 2972
rect 8444 2932 8450 2944
rect 8481 2941 8493 2944
rect 8527 2941 8539 2975
rect 9760 2975 9818 2981
rect 8481 2935 8539 2941
rect 8588 2944 9536 2972
rect 5261 2907 5319 2913
rect 5261 2873 5273 2907
rect 5307 2904 5319 2907
rect 8588 2904 8616 2944
rect 8754 2904 8760 2916
rect 5307 2876 8616 2904
rect 8715 2876 8760 2904
rect 5307 2873 5319 2876
rect 5261 2867 5319 2873
rect 8754 2864 8760 2876
rect 8812 2864 8818 2916
rect 5905 2839 5963 2845
rect 5905 2805 5917 2839
rect 5951 2836 5963 2839
rect 7098 2836 7104 2848
rect 5951 2808 7104 2836
rect 5951 2805 5963 2808
rect 5905 2799 5963 2805
rect 7098 2796 7104 2808
rect 7156 2796 7162 2848
rect 7193 2839 7251 2845
rect 7193 2805 7205 2839
rect 7239 2836 7251 2839
rect 7374 2836 7380 2848
rect 7239 2808 7380 2836
rect 7239 2805 7251 2808
rect 7193 2799 7251 2805
rect 7374 2796 7380 2808
rect 7432 2796 7438 2848
rect 7926 2836 7932 2848
rect 7887 2808 7932 2836
rect 7926 2796 7932 2808
rect 7984 2796 7990 2848
rect 8018 2796 8024 2848
rect 8076 2836 8082 2848
rect 9401 2839 9459 2845
rect 9401 2836 9413 2839
rect 8076 2808 9413 2836
rect 8076 2796 8082 2808
rect 9401 2805 9413 2808
rect 9447 2805 9459 2839
rect 9508 2836 9536 2944
rect 9760 2941 9772 2975
rect 9806 2972 9818 2975
rect 9950 2972 9956 2984
rect 9806 2944 9956 2972
rect 9806 2941 9818 2944
rect 9760 2935 9818 2941
rect 9950 2932 9956 2944
rect 10008 2932 10014 2984
rect 11790 2932 11796 2984
rect 11848 2972 11854 2984
rect 12250 2972 12256 2984
rect 11848 2944 12256 2972
rect 11848 2932 11854 2944
rect 12250 2932 12256 2944
rect 12308 2932 12314 2984
rect 12912 2972 12940 3003
rect 13630 3000 13636 3012
rect 13688 3000 13694 3052
rect 14366 3040 14372 3052
rect 13740 3012 14372 3040
rect 13740 2972 13768 3012
rect 14366 3000 14372 3012
rect 14424 3000 14430 3052
rect 14458 3000 14464 3052
rect 14516 3040 14522 3052
rect 15286 3040 15292 3052
rect 14516 3012 14561 3040
rect 14660 3012 15292 3040
rect 14516 3000 14522 3012
rect 12912 2944 13768 2972
rect 13817 2975 13875 2981
rect 13817 2941 13829 2975
rect 13863 2972 13875 2975
rect 14660 2972 14688 3012
rect 15286 3000 15292 3012
rect 15344 3000 15350 3052
rect 15381 3043 15439 3049
rect 15381 3009 15393 3043
rect 15427 3040 15439 3043
rect 15654 3040 15660 3052
rect 15427 3012 15660 3040
rect 15427 3009 15439 3012
rect 15381 3003 15439 3009
rect 15654 3000 15660 3012
rect 15712 3000 15718 3052
rect 16853 3043 16911 3049
rect 16853 3009 16865 3043
rect 16899 3040 16911 3043
rect 17696 3040 17724 3080
rect 18138 3068 18144 3080
rect 18196 3068 18202 3120
rect 18230 3068 18236 3120
rect 18288 3108 18294 3120
rect 18969 3111 19027 3117
rect 18288 3080 18736 3108
rect 18288 3068 18294 3080
rect 16899 3012 17724 3040
rect 16899 3009 16911 3012
rect 16853 3003 16911 3009
rect 17770 3000 17776 3052
rect 17828 3040 17834 3052
rect 18708 3049 18736 3080
rect 18969 3077 18981 3111
rect 19015 3108 19027 3111
rect 19880 3111 19938 3117
rect 19015 3080 19840 3108
rect 19015 3077 19027 3080
rect 18969 3071 19027 3077
rect 18693 3043 18751 3049
rect 17828 3012 17873 3040
rect 17972 3012 18644 3040
rect 17828 3000 17834 3012
rect 13863 2944 14688 2972
rect 14737 2975 14795 2981
rect 13863 2941 13875 2944
rect 13817 2935 13875 2941
rect 14737 2941 14749 2975
rect 14783 2972 14795 2975
rect 17129 2975 17187 2981
rect 14783 2944 17080 2972
rect 14783 2941 14795 2944
rect 14737 2935 14795 2941
rect 9582 2864 9588 2916
rect 9640 2904 9646 2916
rect 10594 2904 10600 2916
rect 9640 2876 10600 2904
rect 9640 2864 9646 2876
rect 10594 2864 10600 2876
rect 10652 2864 10658 2916
rect 10689 2907 10747 2913
rect 10689 2873 10701 2907
rect 10735 2873 10747 2907
rect 10689 2867 10747 2873
rect 12345 2907 12403 2913
rect 12345 2873 12357 2907
rect 12391 2904 12403 2907
rect 15657 2907 15715 2913
rect 15657 2904 15669 2907
rect 12391 2876 15669 2904
rect 12391 2873 12403 2876
rect 12345 2867 12403 2873
rect 15657 2873 15669 2876
rect 15703 2873 15715 2907
rect 16942 2904 16948 2916
rect 15657 2867 15715 2873
rect 15764 2876 16948 2904
rect 10704 2836 10732 2867
rect 9508 2808 10732 2836
rect 9401 2799 9459 2805
rect 11790 2796 11796 2848
rect 11848 2836 11854 2848
rect 13906 2836 13912 2848
rect 11848 2808 13912 2836
rect 11848 2796 11854 2808
rect 13906 2796 13912 2808
rect 13964 2796 13970 2848
rect 13998 2796 14004 2848
rect 14056 2836 14062 2848
rect 15764 2836 15792 2876
rect 16942 2864 16948 2876
rect 17000 2864 17006 2916
rect 17052 2904 17080 2944
rect 17129 2941 17141 2975
rect 17175 2972 17187 2975
rect 17972 2972 18000 3012
rect 17175 2944 18000 2972
rect 18049 2975 18107 2981
rect 17175 2941 17187 2944
rect 17129 2935 17187 2941
rect 18049 2941 18061 2975
rect 18095 2941 18107 2975
rect 18616 2972 18644 3012
rect 18693 3009 18705 3043
rect 18739 3009 18751 3043
rect 18693 3003 18751 3009
rect 19613 3043 19671 3049
rect 19613 3009 19625 3043
rect 19659 3040 19671 3043
rect 19702 3040 19708 3052
rect 19659 3012 19708 3040
rect 19659 3009 19671 3012
rect 19613 3003 19671 3009
rect 19702 3000 19708 3012
rect 19760 3000 19766 3052
rect 19812 3040 19840 3080
rect 19880 3077 19892 3111
rect 19926 3108 19938 3111
rect 21450 3108 21456 3120
rect 19926 3080 21456 3108
rect 19926 3077 19938 3080
rect 19880 3071 19938 3077
rect 21450 3068 21456 3080
rect 21508 3068 21514 3120
rect 23032 3108 23060 3148
rect 23198 3136 23204 3148
rect 23256 3136 23262 3188
rect 24581 3179 24639 3185
rect 24581 3145 24593 3179
rect 24627 3176 24639 3179
rect 27430 3176 27436 3188
rect 24627 3148 27436 3176
rect 24627 3145 24639 3148
rect 24581 3139 24639 3145
rect 27430 3136 27436 3148
rect 27488 3136 27494 3188
rect 29546 3176 29552 3188
rect 27540 3148 29552 3176
rect 23658 3108 23664 3120
rect 23032 3080 23664 3108
rect 23658 3068 23664 3080
rect 23716 3068 23722 3120
rect 26510 3068 26516 3120
rect 26568 3108 26574 3120
rect 27540 3108 27568 3148
rect 29546 3136 29552 3148
rect 29604 3136 29610 3188
rect 33042 3136 33048 3188
rect 33100 3176 33106 3188
rect 36909 3179 36967 3185
rect 33100 3148 35756 3176
rect 33100 3136 33106 3148
rect 26568 3080 27568 3108
rect 26568 3068 26574 3080
rect 30742 3068 30748 3120
rect 30800 3108 30806 3120
rect 30800 3080 31754 3108
rect 30800 3068 30806 3080
rect 21910 3040 21916 3052
rect 19812 3012 21916 3040
rect 21910 3000 21916 3012
rect 21968 3000 21974 3052
rect 22278 3040 22284 3052
rect 22239 3012 22284 3040
rect 22278 3000 22284 3012
rect 22336 3000 22342 3052
rect 22370 3000 22376 3052
rect 22428 3040 22434 3052
rect 23566 3040 23572 3052
rect 22428 3012 22692 3040
rect 23527 3012 23572 3040
rect 22428 3000 22434 3012
rect 22557 2975 22615 2981
rect 18616 2944 19656 2972
rect 18049 2935 18107 2941
rect 17954 2904 17960 2916
rect 17052 2876 17960 2904
rect 17954 2864 17960 2876
rect 18012 2864 18018 2916
rect 18064 2904 18092 2935
rect 19518 2904 19524 2916
rect 18064 2876 19524 2904
rect 19518 2864 19524 2876
rect 19576 2864 19582 2916
rect 14056 2808 15792 2836
rect 15841 2839 15899 2845
rect 14056 2796 14062 2808
rect 15841 2805 15853 2839
rect 15887 2836 15899 2839
rect 16574 2836 16580 2848
rect 15887 2808 16580 2836
rect 15887 2805 15899 2808
rect 15841 2799 15899 2805
rect 16574 2796 16580 2808
rect 16632 2796 16638 2848
rect 16850 2796 16856 2848
rect 16908 2836 16914 2848
rect 19150 2836 19156 2848
rect 16908 2808 19156 2836
rect 16908 2796 16914 2808
rect 19150 2796 19156 2808
rect 19208 2796 19214 2848
rect 19628 2836 19656 2944
rect 22557 2941 22569 2975
rect 22603 2941 22615 2975
rect 22664 2972 22692 3012
rect 23566 3000 23572 3012
rect 23624 3000 23630 3052
rect 25225 3043 25283 3049
rect 25225 3009 25237 3043
rect 25271 3040 25283 3043
rect 26145 3043 26203 3049
rect 25271 3012 26096 3040
rect 25271 3009 25283 3012
rect 25225 3003 25283 3009
rect 23753 2975 23811 2981
rect 23753 2972 23765 2975
rect 22664 2944 23765 2972
rect 22557 2935 22615 2941
rect 23753 2941 23765 2944
rect 23799 2972 23811 2975
rect 23934 2972 23940 2984
rect 23799 2944 23940 2972
rect 23799 2941 23811 2944
rect 23753 2935 23811 2941
rect 20622 2864 20628 2916
rect 20680 2904 20686 2916
rect 22186 2904 22192 2916
rect 20680 2876 22192 2904
rect 20680 2864 20686 2876
rect 22186 2864 22192 2876
rect 22244 2864 22250 2916
rect 22572 2904 22600 2935
rect 23934 2932 23940 2944
rect 23992 2932 23998 2984
rect 25409 2975 25467 2981
rect 25409 2972 25421 2975
rect 25240 2944 25421 2972
rect 25240 2916 25268 2944
rect 25409 2941 25421 2944
rect 25455 2941 25467 2975
rect 25409 2935 25467 2941
rect 23842 2904 23848 2916
rect 22572 2876 23848 2904
rect 23842 2864 23848 2876
rect 23900 2864 23906 2916
rect 25222 2864 25228 2916
rect 25280 2864 25286 2916
rect 26068 2904 26096 3012
rect 26145 3009 26157 3043
rect 26191 3040 26203 3043
rect 27338 3040 27344 3052
rect 26191 3012 27344 3040
rect 26191 3009 26203 3012
rect 26145 3003 26203 3009
rect 27338 3000 27344 3012
rect 27396 3000 27402 3052
rect 27522 3040 27528 3052
rect 27483 3012 27528 3040
rect 27522 3000 27528 3012
rect 27580 3000 27586 3052
rect 28445 3043 28503 3049
rect 28445 3009 28457 3043
rect 28491 3040 28503 3043
rect 28994 3040 29000 3052
rect 28491 3012 29000 3040
rect 28491 3009 28503 3012
rect 28445 3003 28503 3009
rect 28994 3000 29000 3012
rect 29052 3000 29058 3052
rect 30834 3040 30840 3052
rect 30795 3012 30840 3040
rect 30834 3000 30840 3012
rect 30892 3000 30898 3052
rect 31726 3040 31754 3080
rect 32214 3068 32220 3120
rect 32272 3108 32278 3120
rect 35618 3108 35624 3120
rect 32272 3080 33272 3108
rect 32272 3068 32278 3080
rect 33244 3049 33272 3080
rect 34440 3080 35624 3108
rect 32309 3043 32367 3049
rect 32309 3040 32321 3043
rect 31726 3012 32321 3040
rect 32309 3009 32321 3012
rect 32355 3009 32367 3043
rect 32309 3003 32367 3009
rect 33229 3043 33287 3049
rect 33229 3009 33241 3043
rect 33275 3040 33287 3043
rect 34440 3040 34468 3080
rect 35618 3068 35624 3080
rect 35676 3068 35682 3120
rect 33275 3012 34468 3040
rect 33275 3009 33287 3012
rect 33229 3003 33287 3009
rect 34514 3000 34520 3052
rect 34572 3040 34578 3052
rect 34885 3043 34943 3049
rect 34885 3040 34897 3043
rect 34572 3012 34897 3040
rect 34572 3000 34578 3012
rect 34885 3009 34897 3012
rect 34931 3009 34943 3043
rect 34885 3003 34943 3009
rect 35345 3043 35403 3049
rect 35345 3009 35357 3043
rect 35391 3040 35403 3043
rect 35728 3040 35756 3148
rect 36909 3145 36921 3179
rect 36955 3176 36967 3179
rect 37090 3176 37096 3188
rect 36955 3148 37096 3176
rect 36955 3145 36967 3148
rect 36909 3139 36967 3145
rect 37090 3136 37096 3148
rect 37148 3136 37154 3188
rect 37734 3136 37740 3188
rect 37792 3176 37798 3188
rect 37829 3179 37887 3185
rect 37829 3176 37841 3179
rect 37792 3148 37841 3176
rect 37792 3136 37798 3148
rect 37829 3145 37841 3148
rect 37875 3145 37887 3179
rect 37829 3139 37887 3145
rect 38197 3179 38255 3185
rect 38197 3145 38209 3179
rect 38243 3176 38255 3179
rect 38378 3176 38384 3188
rect 38243 3148 38384 3176
rect 38243 3145 38255 3148
rect 38197 3139 38255 3145
rect 38378 3136 38384 3148
rect 38436 3136 38442 3188
rect 38838 3136 38844 3188
rect 38896 3176 38902 3188
rect 38896 3148 40540 3176
rect 38896 3136 38902 3148
rect 36538 3108 36544 3120
rect 36499 3080 36544 3108
rect 36538 3068 36544 3080
rect 36596 3068 36602 3120
rect 36633 3111 36691 3117
rect 36633 3077 36645 3111
rect 36679 3108 36691 3111
rect 40218 3108 40224 3120
rect 36679 3080 40224 3108
rect 36679 3077 36691 3080
rect 36633 3071 36691 3077
rect 40218 3068 40224 3080
rect 40276 3068 40282 3120
rect 40402 3108 40408 3120
rect 40363 3080 40408 3108
rect 40402 3068 40408 3080
rect 40460 3068 40466 3120
rect 40512 3108 40540 3148
rect 40678 3136 40684 3188
rect 40736 3176 40742 3188
rect 44453 3179 44511 3185
rect 40736 3148 44404 3176
rect 40736 3136 40742 3148
rect 44376 3108 44404 3148
rect 44453 3145 44465 3179
rect 44499 3176 44511 3179
rect 44910 3176 44916 3188
rect 44499 3148 44916 3176
rect 44499 3145 44511 3148
rect 44453 3139 44511 3145
rect 44910 3136 44916 3148
rect 44968 3136 44974 3188
rect 45186 3176 45192 3188
rect 45147 3148 45192 3176
rect 45186 3136 45192 3148
rect 45244 3136 45250 3188
rect 46474 3176 46480 3188
rect 46435 3148 46480 3176
rect 46474 3136 46480 3148
rect 46532 3136 46538 3188
rect 47946 3176 47952 3188
rect 47907 3148 47952 3176
rect 47946 3136 47952 3148
rect 48004 3136 48010 3188
rect 48866 3176 48872 3188
rect 48827 3148 48872 3176
rect 48866 3136 48872 3148
rect 48924 3136 48930 3188
rect 49786 3176 49792 3188
rect 49747 3148 49792 3176
rect 49786 3136 49792 3148
rect 49844 3136 49850 3188
rect 50706 3176 50712 3188
rect 50667 3148 50712 3176
rect 50706 3136 50712 3148
rect 50764 3136 50770 3188
rect 52178 3176 52184 3188
rect 52139 3148 52184 3176
rect 52178 3136 52184 3148
rect 52236 3136 52242 3188
rect 55214 3136 55220 3188
rect 55272 3176 55278 3188
rect 55309 3179 55367 3185
rect 55309 3176 55321 3179
rect 55272 3148 55321 3176
rect 55272 3136 55278 3148
rect 55309 3145 55321 3148
rect 55355 3145 55367 3179
rect 55309 3139 55367 3145
rect 45097 3111 45155 3117
rect 45097 3108 45109 3111
rect 40512 3080 44312 3108
rect 44376 3080 45109 3108
rect 36262 3040 36268 3052
rect 35391 3012 35756 3040
rect 36223 3012 36268 3040
rect 35391 3009 35403 3012
rect 35345 3003 35403 3009
rect 36262 3000 36268 3012
rect 36320 3000 36326 3052
rect 36446 3049 36452 3052
rect 36413 3043 36452 3049
rect 36413 3009 36425 3043
rect 36413 3003 36452 3009
rect 36446 3000 36452 3003
rect 36504 3000 36510 3052
rect 36730 3043 36788 3049
rect 36730 3040 36742 3043
rect 36556 3012 36742 3040
rect 26418 2972 26424 2984
rect 26379 2944 26424 2972
rect 26418 2932 26424 2944
rect 26476 2932 26482 2984
rect 27801 2975 27859 2981
rect 27801 2941 27813 2975
rect 27847 2972 27859 2975
rect 27847 2944 28304 2972
rect 27847 2941 27859 2944
rect 27801 2935 27859 2941
rect 28166 2904 28172 2916
rect 26068 2876 28172 2904
rect 28166 2864 28172 2876
rect 28224 2864 28230 2916
rect 20254 2836 20260 2848
rect 19628 2808 20260 2836
rect 20254 2796 20260 2808
rect 20312 2796 20318 2848
rect 20898 2796 20904 2848
rect 20956 2836 20962 2848
rect 20993 2839 21051 2845
rect 20993 2836 21005 2839
rect 20956 2808 21005 2836
rect 20956 2796 20962 2808
rect 20993 2805 21005 2808
rect 21039 2805 21051 2839
rect 20993 2799 21051 2805
rect 22002 2796 22008 2848
rect 22060 2836 22066 2848
rect 23290 2836 23296 2848
rect 22060 2808 23296 2836
rect 22060 2796 22066 2808
rect 23290 2796 23296 2808
rect 23348 2796 23354 2848
rect 23382 2796 23388 2848
rect 23440 2836 23446 2848
rect 27154 2836 27160 2848
rect 23440 2808 27160 2836
rect 23440 2796 23446 2808
rect 27154 2796 27160 2808
rect 27212 2796 27218 2848
rect 28276 2836 28304 2944
rect 28350 2932 28356 2984
rect 28408 2972 28414 2984
rect 28721 2975 28779 2981
rect 28721 2972 28733 2975
rect 28408 2944 28733 2972
rect 28408 2932 28414 2944
rect 28721 2941 28733 2944
rect 28767 2941 28779 2975
rect 28721 2935 28779 2941
rect 29086 2932 29092 2984
rect 29144 2972 29150 2984
rect 29825 2975 29883 2981
rect 29825 2972 29837 2975
rect 29144 2944 29837 2972
rect 29144 2932 29150 2944
rect 29825 2941 29837 2944
rect 29871 2941 29883 2975
rect 29825 2935 29883 2941
rect 30742 2932 30748 2984
rect 30800 2972 30806 2984
rect 31021 2975 31079 2981
rect 31021 2972 31033 2975
rect 30800 2944 31033 2972
rect 30800 2932 30806 2944
rect 31021 2941 31033 2944
rect 31067 2941 31079 2975
rect 31021 2935 31079 2941
rect 31570 2932 31576 2984
rect 31628 2972 31634 2984
rect 32493 2975 32551 2981
rect 32493 2972 32505 2975
rect 31628 2944 32505 2972
rect 31628 2932 31634 2944
rect 32493 2941 32505 2944
rect 32539 2941 32551 2975
rect 33502 2972 33508 2984
rect 33463 2944 33508 2972
rect 32493 2935 32551 2941
rect 33502 2932 33508 2944
rect 33560 2932 33566 2984
rect 33870 2932 33876 2984
rect 33928 2972 33934 2984
rect 33928 2944 34183 2972
rect 33928 2932 33934 2944
rect 34155 2904 34183 2944
rect 34330 2932 34336 2984
rect 34388 2972 34394 2984
rect 35529 2975 35587 2981
rect 35529 2972 35541 2975
rect 34388 2944 35541 2972
rect 34388 2932 34394 2944
rect 35529 2941 35541 2944
rect 35575 2941 35587 2975
rect 35529 2935 35587 2941
rect 36078 2932 36084 2984
rect 36136 2972 36142 2984
rect 36556 2972 36584 3012
rect 36730 3009 36742 3012
rect 36776 3009 36788 3043
rect 38930 3040 38936 3052
rect 36730 3003 36788 3009
rect 38488 3012 38936 3040
rect 36136 2944 36584 2972
rect 36136 2932 36142 2944
rect 38102 2932 38108 2984
rect 38160 2972 38166 2984
rect 38488 2981 38516 3012
rect 38930 3000 38936 3012
rect 38988 3000 38994 3052
rect 39025 3043 39083 3049
rect 39025 3009 39037 3043
rect 39071 3040 39083 3043
rect 39298 3040 39304 3052
rect 39071 3012 39304 3040
rect 39071 3009 39083 3012
rect 39025 3003 39083 3009
rect 39298 3000 39304 3012
rect 39356 3000 39362 3052
rect 39574 3000 39580 3052
rect 39632 3040 39638 3052
rect 40037 3043 40095 3049
rect 40037 3040 40049 3043
rect 39632 3012 40049 3040
rect 39632 3000 39638 3012
rect 40037 3009 40049 3012
rect 40083 3009 40095 3043
rect 40037 3003 40095 3009
rect 40957 3043 41015 3049
rect 40957 3009 40969 3043
rect 41003 3009 41015 3043
rect 41138 3040 41144 3052
rect 41099 3012 41144 3040
rect 40957 3003 41015 3009
rect 38289 2975 38347 2981
rect 38289 2972 38301 2975
rect 38160 2944 38301 2972
rect 38160 2932 38166 2944
rect 38289 2941 38301 2944
rect 38335 2941 38347 2975
rect 38289 2935 38347 2941
rect 38473 2975 38531 2981
rect 38473 2941 38485 2975
rect 38519 2941 38531 2975
rect 38473 2935 38531 2941
rect 38562 2932 38568 2984
rect 38620 2972 38626 2984
rect 39209 2975 39267 2981
rect 39209 2972 39221 2975
rect 38620 2944 39221 2972
rect 38620 2932 38626 2944
rect 39209 2941 39221 2944
rect 39255 2941 39267 2975
rect 40972 2972 41000 3003
rect 41138 3000 41144 3012
rect 41196 3000 41202 3052
rect 41506 3000 41512 3052
rect 41564 3040 41570 3052
rect 41693 3043 41751 3049
rect 41693 3040 41705 3043
rect 41564 3012 41705 3040
rect 41564 3000 41570 3012
rect 41693 3009 41705 3012
rect 41739 3009 41751 3043
rect 41693 3003 41751 3009
rect 42061 3043 42119 3049
rect 42061 3009 42073 3043
rect 42107 3040 42119 3043
rect 42150 3040 42156 3052
rect 42107 3012 42156 3040
rect 42107 3009 42119 3012
rect 42061 3003 42119 3009
rect 42150 3000 42156 3012
rect 42208 3000 42214 3052
rect 42610 3040 42616 3052
rect 42571 3012 42616 3040
rect 42610 3000 42616 3012
rect 42668 3000 42674 3052
rect 42978 3000 42984 3052
rect 43036 3040 43042 3052
rect 43162 3040 43168 3052
rect 43036 3012 43168 3040
rect 43036 3000 43042 3012
rect 43162 3000 43168 3012
rect 43220 3040 43226 3052
rect 43257 3043 43315 3049
rect 43257 3040 43269 3043
rect 43220 3012 43269 3040
rect 43220 3000 43226 3012
rect 43257 3009 43269 3012
rect 43303 3009 43315 3043
rect 43622 3040 43628 3052
rect 43583 3012 43628 3040
rect 43257 3003 43315 3009
rect 43622 3000 43628 3012
rect 43680 3000 43686 3052
rect 44284 3049 44312 3080
rect 45097 3077 45109 3080
rect 45143 3077 45155 3111
rect 45097 3071 45155 3077
rect 45554 3068 45560 3120
rect 45612 3108 45618 3120
rect 49326 3108 49332 3120
rect 45612 3080 49332 3108
rect 45612 3068 45618 3080
rect 49326 3068 49332 3080
rect 49384 3068 49390 3120
rect 49510 3068 49516 3120
rect 49568 3108 49574 3120
rect 50617 3111 50675 3117
rect 50617 3108 50629 3111
rect 49568 3080 50629 3108
rect 49568 3068 49574 3080
rect 50617 3077 50629 3080
rect 50663 3077 50675 3111
rect 50617 3071 50675 3077
rect 50890 3068 50896 3120
rect 50948 3108 50954 3120
rect 52089 3111 52147 3117
rect 52089 3108 52101 3111
rect 50948 3080 52101 3108
rect 50948 3068 50954 3080
rect 52089 3077 52101 3080
rect 52135 3077 52147 3111
rect 52089 3071 52147 3077
rect 54481 3111 54539 3117
rect 54481 3077 54493 3111
rect 54527 3108 54539 3111
rect 54938 3108 54944 3120
rect 54527 3080 54944 3108
rect 54527 3077 54539 3080
rect 54481 3071 54539 3077
rect 54938 3068 54944 3080
rect 54996 3068 55002 3120
rect 58158 3108 58164 3120
rect 58119 3080 58164 3108
rect 58158 3068 58164 3080
rect 58216 3068 58222 3120
rect 44269 3043 44327 3049
rect 44269 3009 44281 3043
rect 44315 3009 44327 3043
rect 44269 3003 44327 3009
rect 44358 3000 44364 3052
rect 44416 3040 44422 3052
rect 45002 3040 45008 3052
rect 44416 3012 45008 3040
rect 44416 3000 44422 3012
rect 45002 3000 45008 3012
rect 45060 3000 45066 3052
rect 46198 3000 46204 3052
rect 46256 3040 46262 3052
rect 46385 3043 46443 3049
rect 46385 3040 46397 3043
rect 46256 3012 46397 3040
rect 46256 3000 46262 3012
rect 46385 3009 46397 3012
rect 46431 3009 46443 3043
rect 46385 3003 46443 3009
rect 47026 3000 47032 3052
rect 47084 3040 47090 3052
rect 47857 3043 47915 3049
rect 47857 3040 47869 3043
rect 47084 3012 47869 3040
rect 47084 3000 47090 3012
rect 47857 3009 47869 3012
rect 47903 3009 47915 3043
rect 47857 3003 47915 3009
rect 48406 3000 48412 3052
rect 48464 3040 48470 3052
rect 48777 3043 48835 3049
rect 48777 3040 48789 3043
rect 48464 3012 48789 3040
rect 48464 3000 48470 3012
rect 48777 3009 48789 3012
rect 48823 3009 48835 3043
rect 48777 3003 48835 3009
rect 48958 3000 48964 3052
rect 49016 3040 49022 3052
rect 49697 3043 49755 3049
rect 49697 3040 49709 3043
rect 49016 3012 49709 3040
rect 49016 3000 49022 3012
rect 49697 3009 49709 3012
rect 49743 3009 49755 3043
rect 49697 3003 49755 3009
rect 50154 3000 50160 3052
rect 50212 3040 50218 3052
rect 51353 3043 51411 3049
rect 51353 3040 51365 3043
rect 50212 3012 51365 3040
rect 50212 3000 50218 3012
rect 51353 3009 51365 3012
rect 51399 3009 51411 3043
rect 51353 3003 51411 3009
rect 51442 3000 51448 3052
rect 51500 3040 51506 3052
rect 53009 3043 53067 3049
rect 53009 3040 53021 3043
rect 51500 3012 53021 3040
rect 51500 3000 51506 3012
rect 53009 3009 53021 3012
rect 53055 3009 53067 3043
rect 53009 3003 53067 3009
rect 53926 3000 53932 3052
rect 53984 3040 53990 3052
rect 54113 3043 54171 3049
rect 54113 3040 54125 3043
rect 53984 3012 54125 3040
rect 53984 3000 53990 3012
rect 54113 3009 54125 3012
rect 54159 3009 54171 3043
rect 54113 3003 54171 3009
rect 54202 3000 54208 3052
rect 54260 3040 54266 3052
rect 55033 3043 55091 3049
rect 55033 3040 55045 3043
rect 54260 3012 55045 3040
rect 54260 3000 54266 3012
rect 55033 3009 55045 3012
rect 55079 3009 55091 3043
rect 55033 3003 55091 3009
rect 55306 3000 55312 3052
rect 55364 3040 55370 3052
rect 55861 3043 55919 3049
rect 55861 3040 55873 3043
rect 55364 3012 55873 3040
rect 55364 3000 55370 3012
rect 55861 3009 55873 3012
rect 55907 3009 55919 3043
rect 55861 3003 55919 3009
rect 57241 3043 57299 3049
rect 57241 3009 57253 3043
rect 57287 3040 57299 3043
rect 58250 3040 58256 3052
rect 57287 3012 58256 3040
rect 57287 3009 57299 3012
rect 57241 3003 57299 3009
rect 58250 3000 58256 3012
rect 58308 3000 58314 3052
rect 43346 2972 43352 2984
rect 39209 2935 39267 2941
rect 39776 2944 41000 2972
rect 43307 2944 43352 2972
rect 36814 2904 36820 2916
rect 34155 2876 36820 2904
rect 36814 2864 36820 2876
rect 36872 2864 36878 2916
rect 37458 2864 37464 2916
rect 37516 2904 37522 2916
rect 39776 2904 39804 2944
rect 43346 2932 43352 2944
rect 43404 2932 43410 2984
rect 43530 2972 43536 2984
rect 43491 2944 43536 2972
rect 43530 2932 43536 2944
rect 43588 2932 43594 2984
rect 45278 2932 45284 2984
rect 45336 2972 45342 2984
rect 45336 2944 46612 2972
rect 45336 2932 45342 2944
rect 37516 2876 38516 2904
rect 37516 2864 37522 2876
rect 29086 2836 29092 2848
rect 28276 2808 29092 2836
rect 29086 2796 29092 2808
rect 29144 2796 29150 2848
rect 32490 2796 32496 2848
rect 32548 2836 32554 2848
rect 34514 2836 34520 2848
rect 32548 2808 34520 2836
rect 32548 2796 32554 2808
rect 34514 2796 34520 2808
rect 34572 2796 34578 2848
rect 38488 2836 38516 2876
rect 38626 2876 39804 2904
rect 38626 2836 38654 2876
rect 40954 2864 40960 2916
rect 41012 2904 41018 2916
rect 41012 2876 41184 2904
rect 41012 2864 41018 2876
rect 38488 2808 38654 2836
rect 41156 2836 41184 2876
rect 43438 2864 43444 2916
rect 43496 2904 43502 2916
rect 45370 2904 45376 2916
rect 43496 2876 45376 2904
rect 43496 2864 43502 2876
rect 45370 2864 45376 2876
rect 45428 2864 45434 2916
rect 46584 2904 46612 2944
rect 47670 2932 47676 2984
rect 47728 2972 47734 2984
rect 51537 2975 51595 2981
rect 51537 2972 51549 2975
rect 47728 2944 51549 2972
rect 47728 2932 47734 2944
rect 51537 2941 51549 2944
rect 51583 2941 51595 2975
rect 51537 2935 51595 2941
rect 53282 2932 53288 2984
rect 53340 2972 53346 2984
rect 56045 2975 56103 2981
rect 56045 2972 56057 2975
rect 53340 2944 56057 2972
rect 53340 2932 53346 2944
rect 56045 2941 56057 2944
rect 56091 2941 56103 2975
rect 56045 2935 56103 2941
rect 57057 2975 57115 2981
rect 57057 2941 57069 2975
rect 57103 2972 57115 2975
rect 58345 2975 58403 2981
rect 58345 2972 58357 2975
rect 57103 2944 58357 2972
rect 57103 2941 57115 2944
rect 57057 2935 57115 2941
rect 58345 2941 58357 2944
rect 58391 2941 58403 2975
rect 58345 2935 58403 2941
rect 49602 2904 49608 2916
rect 46584 2876 49608 2904
rect 49602 2864 49608 2876
rect 49660 2864 49666 2916
rect 49694 2864 49700 2916
rect 49752 2904 49758 2916
rect 50798 2904 50804 2916
rect 49752 2876 50804 2904
rect 49752 2864 49758 2876
rect 50798 2864 50804 2876
rect 50856 2864 50862 2916
rect 53193 2907 53251 2913
rect 53193 2904 53205 2907
rect 51046 2876 53205 2904
rect 41598 2836 41604 2848
rect 41156 2808 41604 2836
rect 41598 2796 41604 2808
rect 41656 2796 41662 2848
rect 42334 2796 42340 2848
rect 42392 2836 42398 2848
rect 44174 2836 44180 2848
rect 42392 2808 44180 2836
rect 42392 2796 42398 2808
rect 44174 2796 44180 2808
rect 44232 2796 44238 2848
rect 47854 2796 47860 2848
rect 47912 2836 47918 2848
rect 50430 2836 50436 2848
rect 47912 2808 50436 2836
rect 47912 2796 47918 2808
rect 50430 2796 50436 2808
rect 50488 2796 50494 2848
rect 50522 2796 50528 2848
rect 50580 2836 50586 2848
rect 51046 2836 51074 2876
rect 53193 2873 53205 2876
rect 53239 2873 53251 2907
rect 53193 2867 53251 2873
rect 53466 2864 53472 2916
rect 53524 2904 53530 2916
rect 57425 2907 57483 2913
rect 57425 2904 57437 2907
rect 53524 2876 57437 2904
rect 53524 2864 53530 2876
rect 57425 2873 57437 2876
rect 57471 2873 57483 2907
rect 57425 2867 57483 2873
rect 50580 2808 51074 2836
rect 50580 2796 50586 2808
rect 1104 2746 58880 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 58880 2746
rect 1104 2672 58880 2694
rect 3329 2635 3387 2641
rect 3329 2601 3341 2635
rect 3375 2632 3387 2635
rect 7190 2632 7196 2644
rect 3375 2604 7196 2632
rect 3375 2601 3387 2604
rect 3329 2595 3387 2601
rect 7190 2592 7196 2604
rect 7248 2592 7254 2644
rect 7374 2592 7380 2644
rect 7432 2632 7438 2644
rect 9030 2632 9036 2644
rect 7432 2604 9036 2632
rect 7432 2592 7438 2604
rect 9030 2592 9036 2604
rect 9088 2592 9094 2644
rect 11238 2632 11244 2644
rect 9692 2604 11244 2632
rect 5997 2567 6055 2573
rect 5997 2533 6009 2567
rect 6043 2564 6055 2567
rect 7650 2564 7656 2576
rect 6043 2536 7656 2564
rect 6043 2533 6055 2536
rect 5997 2527 6055 2533
rect 7650 2524 7656 2536
rect 7708 2524 7714 2576
rect 9692 2573 9720 2604
rect 11238 2592 11244 2604
rect 11296 2592 11302 2644
rect 11885 2635 11943 2641
rect 11885 2601 11897 2635
rect 11931 2632 11943 2635
rect 13998 2632 14004 2644
rect 11931 2604 14004 2632
rect 11931 2601 11943 2604
rect 11885 2595 11943 2601
rect 13998 2592 14004 2604
rect 14056 2592 14062 2644
rect 14461 2635 14519 2641
rect 14461 2601 14473 2635
rect 14507 2632 14519 2635
rect 17402 2632 17408 2644
rect 14507 2604 17408 2632
rect 14507 2601 14519 2604
rect 14461 2595 14519 2601
rect 17402 2592 17408 2604
rect 17460 2592 17466 2644
rect 19426 2632 19432 2644
rect 18524 2604 19432 2632
rect 9677 2567 9735 2573
rect 9677 2533 9689 2567
rect 9723 2533 9735 2567
rect 9677 2527 9735 2533
rect 10413 2567 10471 2573
rect 10413 2533 10425 2567
rect 10459 2564 10471 2567
rect 11054 2564 11060 2576
rect 10459 2536 11060 2564
rect 10459 2533 10471 2536
rect 10413 2527 10471 2533
rect 11054 2524 11060 2536
rect 11112 2524 11118 2576
rect 11149 2567 11207 2573
rect 11149 2533 11161 2567
rect 11195 2564 11207 2567
rect 12618 2564 12624 2576
rect 11195 2536 12624 2564
rect 11195 2533 11207 2536
rect 11149 2527 11207 2533
rect 12618 2524 12624 2536
rect 12676 2524 12682 2576
rect 18524 2564 18552 2604
rect 19426 2592 19432 2604
rect 19484 2592 19490 2644
rect 19518 2592 19524 2644
rect 19576 2632 19582 2644
rect 21358 2632 21364 2644
rect 19576 2604 21364 2632
rect 19576 2592 19582 2604
rect 21358 2592 21364 2604
rect 21416 2592 21422 2644
rect 26786 2592 26792 2644
rect 26844 2632 26850 2644
rect 26844 2604 31248 2632
rect 26844 2592 26850 2604
rect 20622 2564 20628 2576
rect 14936 2536 18552 2564
rect 18708 2536 20628 2564
rect 7834 2496 7840 2508
rect 5000 2468 7840 2496
rect 1578 2428 1584 2440
rect 1539 2400 1584 2428
rect 1578 2388 1584 2400
rect 1636 2388 1642 2440
rect 3237 2431 3295 2437
rect 3237 2397 3249 2431
rect 3283 2428 3295 2431
rect 4522 2428 4528 2440
rect 3283 2400 4528 2428
rect 3283 2397 3295 2400
rect 3237 2391 3295 2397
rect 4522 2388 4528 2400
rect 4580 2388 4586 2440
rect 1854 2360 1860 2372
rect 1815 2332 1860 2360
rect 1854 2320 1860 2332
rect 1912 2320 1918 2372
rect 4341 2363 4399 2369
rect 4341 2329 4353 2363
rect 4387 2360 4399 2363
rect 5000 2360 5028 2468
rect 7834 2456 7840 2468
rect 7892 2456 7898 2508
rect 9306 2496 9312 2508
rect 9232 2468 9312 2496
rect 5261 2431 5319 2437
rect 5261 2397 5273 2431
rect 5307 2428 5319 2431
rect 6917 2431 6975 2437
rect 5307 2400 6684 2428
rect 5307 2397 5319 2400
rect 5261 2391 5319 2397
rect 4387 2332 5028 2360
rect 5077 2363 5135 2369
rect 4387 2329 4399 2332
rect 4341 2323 4399 2329
rect 5077 2329 5089 2363
rect 5123 2360 5135 2363
rect 5718 2360 5724 2372
rect 5123 2332 5724 2360
rect 5123 2329 5135 2332
rect 5077 2323 5135 2329
rect 5718 2320 5724 2332
rect 5776 2320 5782 2372
rect 5813 2363 5871 2369
rect 5813 2329 5825 2363
rect 5859 2329 5871 2363
rect 6656 2360 6684 2400
rect 6917 2397 6929 2431
rect 6963 2428 6975 2431
rect 9232 2428 9260 2468
rect 9306 2456 9312 2468
rect 9364 2456 9370 2508
rect 13630 2496 13636 2508
rect 10244 2468 13636 2496
rect 10244 2437 10272 2468
rect 13630 2456 13636 2468
rect 13688 2456 13694 2508
rect 10229 2431 10287 2437
rect 6963 2400 9260 2428
rect 9324 2400 10180 2428
rect 6963 2397 6975 2400
rect 6917 2391 6975 2397
rect 7374 2360 7380 2372
rect 6656 2332 7380 2360
rect 5813 2323 5871 2329
rect 4430 2292 4436 2304
rect 4391 2264 4436 2292
rect 4430 2252 4436 2264
rect 4488 2252 4494 2304
rect 5828 2292 5856 2323
rect 7374 2320 7380 2332
rect 7432 2320 7438 2372
rect 7650 2360 7656 2372
rect 7611 2332 7656 2360
rect 7650 2320 7656 2332
rect 7708 2320 7714 2372
rect 8389 2363 8447 2369
rect 8389 2329 8401 2363
rect 8435 2360 8447 2363
rect 9324 2360 9352 2400
rect 9490 2360 9496 2372
rect 8435 2332 9352 2360
rect 9451 2332 9496 2360
rect 8435 2329 8447 2332
rect 8389 2323 8447 2329
rect 9490 2320 9496 2332
rect 9548 2320 9554 2372
rect 10152 2360 10180 2400
rect 10229 2397 10241 2431
rect 10275 2397 10287 2431
rect 10229 2391 10287 2397
rect 10965 2431 11023 2437
rect 10965 2397 10977 2431
rect 11011 2428 11023 2431
rect 11790 2428 11796 2440
rect 11011 2400 11796 2428
rect 11011 2397 11023 2400
rect 10965 2391 11023 2397
rect 11790 2388 11796 2400
rect 11848 2388 11854 2440
rect 12342 2428 12348 2440
rect 12303 2400 12348 2428
rect 12342 2388 12348 2400
rect 12400 2388 12406 2440
rect 12986 2388 12992 2440
rect 13044 2428 13050 2440
rect 14936 2437 14964 2536
rect 15197 2499 15255 2505
rect 15197 2465 15209 2499
rect 15243 2496 15255 2499
rect 16850 2496 16856 2508
rect 15243 2468 16856 2496
rect 15243 2465 15255 2468
rect 15197 2459 15255 2465
rect 16850 2456 16856 2468
rect 16908 2456 16914 2508
rect 17037 2499 17095 2505
rect 17037 2465 17049 2499
rect 17083 2496 17095 2499
rect 17770 2496 17776 2508
rect 17083 2468 17776 2496
rect 17083 2465 17095 2468
rect 17037 2459 17095 2465
rect 17770 2456 17776 2468
rect 17828 2456 17834 2508
rect 18708 2505 18736 2536
rect 20622 2524 20628 2536
rect 20680 2524 20686 2576
rect 28810 2564 28816 2576
rect 26160 2536 28816 2564
rect 18693 2499 18751 2505
rect 18693 2465 18705 2499
rect 18739 2465 18751 2499
rect 20165 2499 20223 2505
rect 18693 2459 18751 2465
rect 19168 2468 20116 2496
rect 13265 2431 13323 2437
rect 13265 2428 13277 2431
rect 13044 2400 13277 2428
rect 13044 2388 13050 2400
rect 13265 2397 13277 2400
rect 13311 2397 13323 2431
rect 13265 2391 13323 2397
rect 14921 2431 14979 2437
rect 14921 2397 14933 2431
rect 14967 2397 14979 2431
rect 14921 2391 14979 2397
rect 15841 2431 15899 2437
rect 15841 2397 15853 2431
rect 15887 2428 15899 2431
rect 17310 2428 17316 2440
rect 15887 2400 17316 2428
rect 15887 2397 15899 2400
rect 15841 2391 15899 2397
rect 17310 2388 17316 2400
rect 17368 2388 17374 2440
rect 17494 2428 17500 2440
rect 17455 2400 17500 2428
rect 17494 2388 17500 2400
rect 17552 2388 17558 2440
rect 18414 2428 18420 2440
rect 18375 2400 18420 2428
rect 18414 2388 18420 2400
rect 18472 2388 18478 2440
rect 11422 2360 11428 2372
rect 10152 2332 11428 2360
rect 11422 2320 11428 2332
rect 11480 2320 11486 2372
rect 12621 2363 12679 2369
rect 12621 2329 12633 2363
rect 12667 2329 12679 2363
rect 12621 2323 12679 2329
rect 13541 2363 13599 2369
rect 13541 2329 13553 2363
rect 13587 2360 13599 2363
rect 15746 2360 15752 2372
rect 13587 2332 15752 2360
rect 13587 2329 13599 2332
rect 13541 2323 13599 2329
rect 6914 2292 6920 2304
rect 5828 2264 6920 2292
rect 6914 2252 6920 2264
rect 6972 2252 6978 2304
rect 7009 2295 7067 2301
rect 7009 2261 7021 2295
rect 7055 2292 7067 2295
rect 7466 2292 7472 2304
rect 7055 2264 7472 2292
rect 7055 2261 7067 2264
rect 7009 2255 7067 2261
rect 7466 2252 7472 2264
rect 7524 2252 7530 2304
rect 7742 2292 7748 2304
rect 7703 2264 7748 2292
rect 7742 2252 7748 2264
rect 7800 2252 7806 2304
rect 8478 2292 8484 2304
rect 8439 2264 8484 2292
rect 8478 2252 8484 2264
rect 8536 2252 8542 2304
rect 9214 2252 9220 2304
rect 9272 2292 9278 2304
rect 10870 2292 10876 2304
rect 9272 2264 10876 2292
rect 9272 2252 9278 2264
rect 10870 2252 10876 2264
rect 10928 2252 10934 2304
rect 12636 2292 12664 2323
rect 15746 2320 15752 2332
rect 15804 2320 15810 2372
rect 16117 2363 16175 2369
rect 16117 2329 16129 2363
rect 16163 2360 16175 2363
rect 17773 2363 17831 2369
rect 16163 2332 16574 2360
rect 16163 2329 16175 2332
rect 16117 2323 16175 2329
rect 15010 2292 15016 2304
rect 12636 2264 15016 2292
rect 15010 2252 15016 2264
rect 15068 2252 15074 2304
rect 16546 2292 16574 2332
rect 17773 2329 17785 2363
rect 17819 2360 17831 2363
rect 19168 2360 19196 2468
rect 19886 2428 19892 2440
rect 19847 2400 19892 2428
rect 19886 2388 19892 2400
rect 19944 2388 19950 2440
rect 20088 2428 20116 2468
rect 20165 2465 20177 2499
rect 20211 2496 20223 2499
rect 22002 2496 22008 2508
rect 20211 2468 22008 2496
rect 20211 2465 20223 2468
rect 20165 2459 20223 2465
rect 22002 2456 22008 2468
rect 22060 2456 22066 2508
rect 22925 2499 22983 2505
rect 22925 2465 22937 2499
rect 22971 2496 22983 2499
rect 24394 2496 24400 2508
rect 22971 2468 24400 2496
rect 22971 2465 22983 2468
rect 22925 2459 22983 2465
rect 24394 2456 24400 2468
rect 24452 2456 24458 2508
rect 20717 2431 20775 2437
rect 20088 2400 20668 2428
rect 20070 2360 20076 2372
rect 17819 2332 19196 2360
rect 19306 2332 20076 2360
rect 17819 2329 17831 2332
rect 17773 2323 17831 2329
rect 19306 2292 19334 2332
rect 20070 2320 20076 2332
rect 20128 2320 20134 2372
rect 19426 2292 19432 2304
rect 16546 2264 19334 2292
rect 19387 2264 19432 2292
rect 19426 2252 19432 2264
rect 19484 2252 19490 2304
rect 19518 2252 19524 2304
rect 19576 2292 19582 2304
rect 20438 2292 20444 2304
rect 19576 2264 20444 2292
rect 19576 2252 19582 2264
rect 20438 2252 20444 2264
rect 20496 2252 20502 2304
rect 20640 2292 20668 2400
rect 20717 2397 20729 2431
rect 20763 2428 20775 2431
rect 20990 2428 20996 2440
rect 20763 2400 20996 2428
rect 20763 2397 20775 2400
rect 20717 2391 20775 2397
rect 20990 2388 20996 2400
rect 21048 2388 21054 2440
rect 22646 2428 22652 2440
rect 22607 2400 22652 2428
rect 22646 2388 22652 2400
rect 22704 2388 22710 2440
rect 23569 2431 23627 2437
rect 23569 2397 23581 2431
rect 23615 2397 23627 2431
rect 23569 2391 23627 2397
rect 21269 2363 21327 2369
rect 21269 2329 21281 2363
rect 21315 2360 21327 2363
rect 23474 2360 23480 2372
rect 21315 2332 23480 2360
rect 21315 2329 21327 2332
rect 21269 2323 21327 2329
rect 23474 2320 23480 2332
rect 23532 2320 23538 2372
rect 23584 2360 23612 2391
rect 23658 2388 23664 2440
rect 23716 2428 23722 2440
rect 26160 2437 26188 2536
rect 28810 2524 28816 2536
rect 28868 2524 28874 2576
rect 28077 2499 28135 2505
rect 28077 2465 28089 2499
rect 28123 2496 28135 2499
rect 29362 2496 29368 2508
rect 28123 2468 29368 2496
rect 28123 2465 28135 2468
rect 28077 2459 28135 2465
rect 29362 2456 29368 2468
rect 29420 2456 29426 2508
rect 25225 2431 25283 2437
rect 25225 2428 25237 2431
rect 23716 2400 25237 2428
rect 23716 2388 23722 2400
rect 25225 2397 25237 2400
rect 25271 2397 25283 2431
rect 25225 2391 25283 2397
rect 26145 2431 26203 2437
rect 26145 2397 26157 2431
rect 26191 2397 26203 2431
rect 26145 2391 26203 2397
rect 27801 2431 27859 2437
rect 27801 2397 27813 2431
rect 27847 2428 27859 2431
rect 27890 2428 27896 2440
rect 27847 2400 27896 2428
rect 27847 2397 27859 2400
rect 27801 2391 27859 2397
rect 27890 2388 27896 2400
rect 27948 2388 27954 2440
rect 28721 2431 28779 2437
rect 28721 2397 28733 2431
rect 28767 2428 28779 2431
rect 28902 2428 28908 2440
rect 28767 2400 28908 2428
rect 28767 2397 28779 2400
rect 28721 2391 28779 2397
rect 28902 2388 28908 2400
rect 28960 2388 28966 2440
rect 29178 2388 29184 2440
rect 29236 2428 29242 2440
rect 30193 2431 30251 2437
rect 30193 2428 30205 2431
rect 29236 2400 30205 2428
rect 29236 2388 29242 2400
rect 30193 2397 30205 2400
rect 30239 2397 30251 2431
rect 30193 2391 30251 2397
rect 30926 2388 30932 2440
rect 30984 2428 30990 2440
rect 31113 2431 31171 2437
rect 31113 2428 31125 2431
rect 30984 2400 31125 2428
rect 30984 2388 30990 2400
rect 31113 2397 31125 2400
rect 31159 2397 31171 2431
rect 31220 2428 31248 2604
rect 34330 2592 34336 2644
rect 34388 2632 34394 2644
rect 34388 2604 38608 2632
rect 34388 2592 34394 2604
rect 34238 2524 34244 2576
rect 34296 2564 34302 2576
rect 34296 2536 36124 2564
rect 34296 2524 34302 2536
rect 31294 2456 31300 2508
rect 31352 2496 31358 2508
rect 32493 2499 32551 2505
rect 32493 2496 32505 2499
rect 31352 2468 32505 2496
rect 31352 2456 31358 2468
rect 32493 2465 32505 2468
rect 32539 2465 32551 2499
rect 32493 2459 32551 2465
rect 34514 2456 34520 2508
rect 34572 2496 34578 2508
rect 35989 2499 36047 2505
rect 35989 2496 36001 2499
rect 34572 2468 36001 2496
rect 34572 2456 34578 2468
rect 35989 2465 36001 2468
rect 36035 2465 36047 2499
rect 35989 2459 36047 2465
rect 32309 2431 32367 2437
rect 32309 2428 32321 2431
rect 31220 2400 32321 2428
rect 31113 2391 31171 2397
rect 32309 2397 32321 2400
rect 32355 2397 32367 2431
rect 32309 2391 32367 2397
rect 32398 2388 32404 2440
rect 32456 2428 32462 2440
rect 33229 2431 33287 2437
rect 33229 2428 33241 2431
rect 32456 2400 33241 2428
rect 32456 2388 32462 2400
rect 33229 2397 33241 2400
rect 33275 2397 33287 2431
rect 34882 2428 34888 2440
rect 34843 2400 34888 2428
rect 33229 2391 33287 2397
rect 34882 2388 34888 2400
rect 34940 2388 34946 2440
rect 35805 2431 35863 2437
rect 35805 2428 35817 2431
rect 34992 2400 35817 2428
rect 23750 2360 23756 2372
rect 23584 2332 23756 2360
rect 23750 2320 23756 2332
rect 23808 2320 23814 2372
rect 23845 2363 23903 2369
rect 23845 2329 23857 2363
rect 23891 2360 23903 2363
rect 24946 2360 24952 2372
rect 23891 2332 24952 2360
rect 23891 2329 23903 2332
rect 23845 2323 23903 2329
rect 24946 2320 24952 2332
rect 25004 2320 25010 2372
rect 25498 2360 25504 2372
rect 25459 2332 25504 2360
rect 25498 2320 25504 2332
rect 25556 2320 25562 2372
rect 26421 2363 26479 2369
rect 26421 2329 26433 2363
rect 26467 2360 26479 2363
rect 28810 2360 28816 2372
rect 26467 2332 28816 2360
rect 26467 2329 26479 2332
rect 26421 2323 26479 2329
rect 28810 2320 28816 2332
rect 28868 2320 28874 2372
rect 28997 2363 29055 2369
rect 28997 2329 29009 2363
rect 29043 2360 29055 2363
rect 29914 2360 29920 2372
rect 29043 2332 29920 2360
rect 29043 2329 29055 2332
rect 28997 2323 29055 2329
rect 29914 2320 29920 2332
rect 29972 2320 29978 2372
rect 30466 2360 30472 2372
rect 30427 2332 30472 2360
rect 30466 2320 30472 2332
rect 30524 2320 30530 2372
rect 31018 2320 31024 2372
rect 31076 2360 31082 2372
rect 31389 2363 31447 2369
rect 31389 2360 31401 2363
rect 31076 2332 31401 2360
rect 31076 2320 31082 2332
rect 31389 2329 31401 2332
rect 31435 2329 31447 2363
rect 31389 2323 31447 2329
rect 31846 2320 31852 2372
rect 31904 2360 31910 2372
rect 33505 2363 33563 2369
rect 33505 2360 33517 2363
rect 31904 2332 33517 2360
rect 31904 2320 31910 2332
rect 33505 2329 33517 2332
rect 33551 2329 33563 2363
rect 33505 2323 33563 2329
rect 33870 2320 33876 2372
rect 33928 2360 33934 2372
rect 34992 2360 35020 2400
rect 35805 2397 35817 2400
rect 35851 2397 35863 2431
rect 36096 2428 36124 2536
rect 36906 2456 36912 2508
rect 36964 2496 36970 2508
rect 38580 2505 38608 2604
rect 40862 2592 40868 2644
rect 40920 2632 40926 2644
rect 40920 2604 41414 2632
rect 40920 2592 40926 2604
rect 41386 2564 41414 2604
rect 42794 2592 42800 2644
rect 42852 2632 42858 2644
rect 45002 2632 45008 2644
rect 42852 2604 45008 2632
rect 42852 2592 42858 2604
rect 45002 2592 45008 2604
rect 45060 2592 45066 2644
rect 45370 2632 45376 2644
rect 45331 2604 45376 2632
rect 45370 2592 45376 2604
rect 45428 2592 45434 2644
rect 46106 2592 46112 2644
rect 46164 2632 46170 2644
rect 46201 2635 46259 2641
rect 46201 2632 46213 2635
rect 46164 2604 46213 2632
rect 46164 2592 46170 2604
rect 46201 2601 46213 2604
rect 46247 2601 46259 2635
rect 47118 2632 47124 2644
rect 47079 2604 47124 2632
rect 46201 2595 46259 2601
rect 47118 2592 47124 2604
rect 47176 2592 47182 2644
rect 47762 2592 47768 2644
rect 47820 2632 47826 2644
rect 47949 2635 48007 2641
rect 47949 2632 47961 2635
rect 47820 2604 47961 2632
rect 47820 2592 47826 2604
rect 47949 2601 47961 2604
rect 47995 2601 48007 2635
rect 47949 2595 48007 2601
rect 48682 2592 48688 2644
rect 48740 2632 48746 2644
rect 48869 2635 48927 2641
rect 48869 2632 48881 2635
rect 48740 2604 48881 2632
rect 48740 2592 48746 2604
rect 48869 2601 48881 2604
rect 48915 2601 48927 2635
rect 48869 2595 48927 2601
rect 49050 2592 49056 2644
rect 49108 2632 49114 2644
rect 58250 2632 58256 2644
rect 49108 2604 55720 2632
rect 58211 2604 58256 2632
rect 49108 2592 49114 2604
rect 50617 2567 50675 2573
rect 50617 2564 50629 2567
rect 41386 2536 50629 2564
rect 50617 2533 50629 2536
rect 50663 2533 50675 2567
rect 50617 2527 50675 2533
rect 50706 2524 50712 2576
rect 50764 2564 50770 2576
rect 52089 2567 52147 2573
rect 52089 2564 52101 2567
rect 50764 2536 52101 2564
rect 50764 2524 50770 2536
rect 52089 2533 52101 2536
rect 52135 2533 52147 2567
rect 52089 2527 52147 2533
rect 37645 2499 37703 2505
rect 37645 2496 37657 2499
rect 36964 2468 37657 2496
rect 36964 2456 36970 2468
rect 37645 2465 37657 2468
rect 37691 2465 37703 2499
rect 37645 2459 37703 2465
rect 38565 2499 38623 2505
rect 38565 2465 38577 2499
rect 38611 2465 38623 2499
rect 41325 2499 41383 2505
rect 41325 2496 41337 2499
rect 38565 2459 38623 2465
rect 38672 2468 41337 2496
rect 37461 2431 37519 2437
rect 37461 2428 37473 2431
rect 36096 2400 37473 2428
rect 35805 2391 35863 2397
rect 37461 2397 37473 2400
rect 37507 2397 37519 2431
rect 37461 2391 37519 2397
rect 37918 2388 37924 2440
rect 37976 2428 37982 2440
rect 38381 2431 38439 2437
rect 38381 2428 38393 2431
rect 37976 2400 38393 2428
rect 37976 2388 37982 2400
rect 38381 2397 38393 2400
rect 38427 2397 38439 2431
rect 38381 2391 38439 2397
rect 33928 2332 35020 2360
rect 35161 2363 35219 2369
rect 33928 2320 33934 2332
rect 35161 2329 35173 2363
rect 35207 2329 35219 2363
rect 35161 2323 35219 2329
rect 21634 2292 21640 2304
rect 20640 2264 21640 2292
rect 21634 2252 21640 2264
rect 21692 2252 21698 2304
rect 22005 2295 22063 2301
rect 22005 2261 22017 2295
rect 22051 2292 22063 2295
rect 23382 2292 23388 2304
rect 22051 2264 23388 2292
rect 22051 2261 22063 2264
rect 22005 2255 22063 2261
rect 23382 2252 23388 2264
rect 23440 2252 23446 2304
rect 24581 2295 24639 2301
rect 24581 2261 24593 2295
rect 24627 2292 24639 2295
rect 26142 2292 26148 2304
rect 24627 2264 26148 2292
rect 24627 2261 24639 2264
rect 24581 2255 24639 2261
rect 26142 2252 26148 2264
rect 26200 2252 26206 2304
rect 26878 2252 26884 2304
rect 26936 2292 26942 2304
rect 27157 2295 27215 2301
rect 27157 2292 27169 2295
rect 26936 2264 27169 2292
rect 26936 2252 26942 2264
rect 27157 2261 27169 2264
rect 27203 2261 27215 2295
rect 27157 2255 27215 2261
rect 32122 2252 32128 2304
rect 32180 2292 32186 2304
rect 35176 2292 35204 2323
rect 36630 2320 36636 2372
rect 36688 2360 36694 2372
rect 38672 2360 38700 2468
rect 41325 2465 41337 2468
rect 41371 2465 41383 2499
rect 41325 2459 41383 2465
rect 42978 2456 42984 2508
rect 43036 2456 43042 2508
rect 45002 2456 45008 2508
rect 45060 2496 45066 2508
rect 45060 2468 49188 2496
rect 45060 2456 45066 2468
rect 40218 2388 40224 2440
rect 40276 2428 40282 2440
rect 41049 2431 41107 2437
rect 41049 2428 41061 2431
rect 40276 2400 41061 2428
rect 40276 2388 40282 2400
rect 41049 2397 41061 2400
rect 41095 2397 41107 2431
rect 42610 2428 42616 2440
rect 42571 2400 42616 2428
rect 41049 2391 41107 2397
rect 42610 2388 42616 2400
rect 42668 2388 42674 2440
rect 42794 2437 42800 2440
rect 42761 2431 42800 2437
rect 42761 2397 42773 2431
rect 42761 2391 42800 2397
rect 42794 2388 42800 2391
rect 42852 2388 42858 2440
rect 42889 2431 42947 2437
rect 42889 2397 42901 2431
rect 42935 2428 42947 2431
rect 42996 2428 43024 2456
rect 42935 2400 43024 2428
rect 43119 2431 43177 2437
rect 42935 2397 42947 2400
rect 42889 2391 42947 2397
rect 43119 2397 43131 2431
rect 43165 2428 43177 2431
rect 43530 2428 43536 2440
rect 43165 2400 43536 2428
rect 43165 2397 43177 2400
rect 43119 2391 43177 2397
rect 43530 2388 43536 2400
rect 43588 2388 43594 2440
rect 44450 2428 44456 2440
rect 43732 2400 44456 2428
rect 36688 2332 38700 2360
rect 36688 2320 36694 2332
rect 39298 2320 39304 2372
rect 39356 2360 39362 2372
rect 40129 2363 40187 2369
rect 40129 2360 40141 2363
rect 39356 2332 40141 2360
rect 39356 2320 39362 2332
rect 40129 2329 40141 2332
rect 40175 2329 40187 2363
rect 40129 2323 40187 2329
rect 42981 2363 43039 2369
rect 42981 2329 42993 2363
rect 43027 2360 43039 2363
rect 43732 2360 43760 2400
rect 44450 2388 44456 2400
rect 44508 2388 44514 2440
rect 45186 2428 45192 2440
rect 45147 2400 45192 2428
rect 45186 2388 45192 2400
rect 45244 2388 45250 2440
rect 46474 2388 46480 2440
rect 46532 2428 46538 2440
rect 47857 2431 47915 2437
rect 47857 2428 47869 2431
rect 46532 2400 47869 2428
rect 46532 2388 46538 2400
rect 47857 2397 47869 2400
rect 47903 2397 47915 2431
rect 49160 2428 49188 2468
rect 49234 2456 49240 2508
rect 49292 2496 49298 2508
rect 49292 2468 50568 2496
rect 49292 2456 49298 2468
rect 49694 2428 49700 2440
rect 49160 2400 49700 2428
rect 47857 2391 47915 2397
rect 49694 2388 49700 2400
rect 49752 2388 49758 2440
rect 50430 2428 50436 2440
rect 50391 2400 50436 2428
rect 50430 2388 50436 2400
rect 50488 2388 50494 2440
rect 50540 2428 50568 2468
rect 50982 2456 50988 2508
rect 51040 2496 51046 2508
rect 55692 2505 55720 2604
rect 58250 2592 58256 2604
rect 58308 2592 58314 2644
rect 54021 2499 54079 2505
rect 54021 2496 54033 2499
rect 51040 2468 54033 2496
rect 51040 2456 51046 2468
rect 54021 2465 54033 2468
rect 54067 2465 54079 2499
rect 54021 2459 54079 2465
rect 55677 2499 55735 2505
rect 55677 2465 55689 2499
rect 55723 2465 55735 2499
rect 55677 2459 55735 2465
rect 51169 2431 51227 2437
rect 51169 2428 51181 2431
rect 50540 2400 51181 2428
rect 51169 2397 51181 2400
rect 51215 2397 51227 2431
rect 51169 2391 51227 2397
rect 53650 2388 53656 2440
rect 53708 2428 53714 2440
rect 53837 2431 53895 2437
rect 53837 2428 53849 2431
rect 53708 2400 53849 2428
rect 53708 2388 53714 2400
rect 53837 2397 53849 2400
rect 53883 2397 53895 2431
rect 53837 2391 53895 2397
rect 55030 2388 55036 2440
rect 55088 2428 55094 2440
rect 55493 2431 55551 2437
rect 55493 2428 55505 2431
rect 55088 2400 55505 2428
rect 55088 2388 55094 2400
rect 55493 2397 55505 2400
rect 55539 2397 55551 2431
rect 55493 2391 55551 2397
rect 57057 2431 57115 2437
rect 57057 2397 57069 2431
rect 57103 2428 57115 2431
rect 57238 2428 57244 2440
rect 57103 2400 57244 2428
rect 57103 2397 57115 2400
rect 57057 2391 57115 2397
rect 57238 2388 57244 2400
rect 57296 2388 57302 2440
rect 58158 2428 58164 2440
rect 58119 2400 58164 2428
rect 58158 2388 58164 2400
rect 58216 2388 58222 2440
rect 43898 2360 43904 2372
rect 43027 2332 43760 2360
rect 43859 2332 43904 2360
rect 43027 2329 43039 2332
rect 42981 2323 43039 2329
rect 43898 2320 43904 2332
rect 43956 2320 43962 2372
rect 45922 2320 45928 2372
rect 45980 2360 45986 2372
rect 46109 2363 46167 2369
rect 46109 2360 46121 2363
rect 45980 2332 46121 2360
rect 45980 2320 45986 2332
rect 46109 2329 46121 2332
rect 46155 2329 46167 2363
rect 46109 2323 46167 2329
rect 47029 2363 47087 2369
rect 47029 2329 47041 2363
rect 47075 2329 47087 2363
rect 47029 2323 47087 2329
rect 32180 2264 35204 2292
rect 32180 2252 32186 2264
rect 35526 2252 35532 2304
rect 35584 2292 35590 2304
rect 40221 2295 40279 2301
rect 40221 2292 40233 2295
rect 35584 2264 40233 2292
rect 35584 2252 35590 2264
rect 40221 2261 40233 2264
rect 40267 2261 40279 2295
rect 40221 2255 40279 2261
rect 42242 2252 42248 2304
rect 42300 2292 42306 2304
rect 43257 2295 43315 2301
rect 43257 2292 43269 2295
rect 42300 2264 43269 2292
rect 42300 2252 42306 2264
rect 43257 2261 43269 2264
rect 43303 2261 43315 2295
rect 43257 2255 43315 2261
rect 43346 2252 43352 2304
rect 43404 2292 43410 2304
rect 43993 2295 44051 2301
rect 43993 2292 44005 2295
rect 43404 2264 44005 2292
rect 43404 2252 43410 2264
rect 43993 2261 44005 2264
rect 44039 2261 44051 2295
rect 43993 2255 44051 2261
rect 44174 2252 44180 2304
rect 44232 2292 44238 2304
rect 47044 2292 47072 2323
rect 47302 2320 47308 2372
rect 47360 2360 47366 2372
rect 48777 2363 48835 2369
rect 48777 2360 48789 2363
rect 47360 2332 48789 2360
rect 47360 2320 47366 2332
rect 48777 2329 48789 2332
rect 48823 2329 48835 2363
rect 51905 2363 51963 2369
rect 51905 2360 51917 2363
rect 48777 2323 48835 2329
rect 51092 2332 51917 2360
rect 44232 2264 47072 2292
rect 44232 2252 44238 2264
rect 50062 2252 50068 2304
rect 50120 2292 50126 2304
rect 51092 2292 51120 2332
rect 51905 2329 51917 2332
rect 51951 2329 51963 2363
rect 51905 2323 51963 2329
rect 52546 2320 52552 2372
rect 52604 2360 52610 2372
rect 53009 2363 53067 2369
rect 53009 2360 53021 2363
rect 52604 2332 53021 2360
rect 52604 2320 52610 2332
rect 53009 2329 53021 2332
rect 53055 2329 53067 2363
rect 57330 2360 57336 2372
rect 57291 2332 57336 2360
rect 53009 2323 53067 2329
rect 57330 2320 57336 2332
rect 57388 2320 57394 2372
rect 51258 2292 51264 2304
rect 50120 2264 51120 2292
rect 51219 2264 51264 2292
rect 50120 2252 50126 2264
rect 51258 2252 51264 2264
rect 51316 2252 51322 2304
rect 53098 2292 53104 2304
rect 53059 2264 53104 2292
rect 53098 2252 53104 2264
rect 53156 2252 53162 2304
rect 1104 2202 58880 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 58880 2202
rect 1104 2128 58880 2150
rect 1578 2048 1584 2100
rect 1636 2088 1642 2100
rect 1636 2060 17264 2088
rect 1636 2048 1642 2060
rect 4430 1980 4436 2032
rect 4488 2020 4494 2032
rect 8662 2020 8668 2032
rect 4488 1992 8668 2020
rect 4488 1980 4494 1992
rect 8662 1980 8668 1992
rect 8720 1980 8726 2032
rect 9490 1980 9496 2032
rect 9548 2020 9554 2032
rect 12802 2020 12808 2032
rect 9548 1992 12808 2020
rect 9548 1980 9554 1992
rect 12802 1980 12808 1992
rect 12860 1980 12866 2032
rect 8478 1912 8484 1964
rect 8536 1952 8542 1964
rect 11330 1952 11336 1964
rect 8536 1924 11336 1952
rect 8536 1912 8542 1924
rect 11330 1912 11336 1924
rect 11388 1912 11394 1964
rect 17236 1952 17264 2060
rect 19426 2048 19432 2100
rect 19484 2088 19490 2100
rect 27982 2088 27988 2100
rect 19484 2060 27988 2088
rect 19484 2048 19490 2060
rect 27982 2048 27988 2060
rect 28040 2048 28046 2100
rect 41046 2048 41052 2100
rect 41104 2088 41110 2100
rect 43346 2088 43352 2100
rect 41104 2060 43352 2088
rect 41104 2048 41110 2060
rect 43346 2048 43352 2060
rect 43404 2048 43410 2100
rect 43622 2048 43628 2100
rect 43680 2088 43686 2100
rect 50706 2088 50712 2100
rect 43680 2060 50712 2088
rect 43680 2048 43686 2060
rect 50706 2048 50712 2060
rect 50764 2048 50770 2100
rect 18414 1980 18420 2032
rect 18472 2020 18478 2032
rect 22830 2020 22836 2032
rect 18472 1992 22836 2020
rect 18472 1980 18478 1992
rect 22830 1980 22836 1992
rect 22888 1980 22894 2032
rect 23750 1980 23756 2032
rect 23808 2020 23814 2032
rect 23808 1992 35020 2020
rect 23808 1980 23814 1992
rect 26694 1952 26700 1964
rect 17236 1924 26700 1952
rect 26694 1912 26700 1924
rect 26752 1912 26758 1964
rect 26970 1912 26976 1964
rect 27028 1952 27034 1964
rect 34882 1952 34888 1964
rect 27028 1924 34888 1952
rect 27028 1912 27034 1924
rect 34882 1912 34888 1924
rect 34940 1912 34946 1964
rect 7650 1844 7656 1896
rect 7708 1884 7714 1896
rect 11146 1884 11152 1896
rect 7708 1856 11152 1884
rect 7708 1844 7714 1856
rect 11146 1844 11152 1856
rect 11204 1844 11210 1896
rect 7742 1776 7748 1828
rect 7800 1816 7806 1828
rect 12710 1816 12716 1828
rect 7800 1788 12716 1816
rect 7800 1776 7806 1788
rect 12710 1776 12716 1788
rect 12768 1776 12774 1828
rect 13170 1776 13176 1828
rect 13228 1816 13234 1828
rect 23658 1816 23664 1828
rect 13228 1788 23664 1816
rect 13228 1776 13234 1788
rect 23658 1776 23664 1788
rect 23716 1776 23722 1828
rect 34992 1816 35020 1992
rect 36998 1980 37004 2032
rect 37056 2020 37062 2032
rect 42242 2020 42248 2032
rect 37056 1992 42248 2020
rect 37056 1980 37062 1992
rect 42242 1980 42248 1992
rect 42300 1980 42306 2032
rect 39758 1912 39764 1964
rect 39816 1952 39822 1964
rect 51258 1952 51264 1964
rect 39816 1924 51264 1952
rect 39816 1912 39822 1924
rect 51258 1912 51264 1924
rect 51316 1912 51322 1964
rect 36906 1844 36912 1896
rect 36964 1884 36970 1896
rect 53098 1884 53104 1896
rect 36964 1856 53104 1884
rect 36964 1844 36970 1856
rect 53098 1844 53104 1856
rect 53156 1844 53162 1896
rect 34992 1788 38654 1816
rect 7466 1708 7472 1760
rect 7524 1748 7530 1760
rect 13262 1748 13268 1760
rect 7524 1720 13268 1748
rect 7524 1708 7530 1720
rect 13262 1708 13268 1720
rect 13320 1708 13326 1760
rect 17310 1708 17316 1760
rect 17368 1748 17374 1760
rect 20162 1748 20168 1760
rect 17368 1720 20168 1748
rect 17368 1708 17374 1720
rect 20162 1708 20168 1720
rect 20220 1708 20226 1760
rect 26050 1708 26056 1760
rect 26108 1748 26114 1760
rect 38626 1748 38654 1788
rect 43070 1748 43076 1760
rect 26108 1720 28994 1748
rect 38626 1720 43076 1748
rect 26108 1708 26114 1720
rect 28966 1680 28994 1720
rect 43070 1708 43076 1720
rect 43128 1708 43134 1760
rect 36906 1680 36912 1692
rect 28966 1652 36912 1680
rect 36906 1640 36912 1652
rect 36964 1640 36970 1692
rect 37918 1640 37924 1692
rect 37976 1680 37982 1692
rect 43898 1680 43904 1692
rect 37976 1652 43904 1680
rect 37976 1640 37982 1652
rect 43898 1640 43904 1652
rect 43956 1640 43962 1692
rect 26418 1504 26424 1556
rect 26476 1544 26482 1556
rect 28534 1544 28540 1556
rect 26476 1516 28540 1544
rect 26476 1504 26482 1516
rect 28534 1504 28540 1516
rect 28592 1504 28598 1556
rect 35710 1504 35716 1556
rect 35768 1544 35774 1556
rect 36722 1544 36728 1556
rect 35768 1516 36728 1544
rect 35768 1504 35774 1516
rect 36722 1504 36728 1516
rect 36780 1504 36786 1556
rect 6914 1436 6920 1488
rect 6972 1476 6978 1488
rect 10042 1476 10048 1488
rect 6972 1448 10048 1476
rect 6972 1436 6978 1448
rect 10042 1436 10048 1448
rect 10100 1436 10106 1488
rect 5718 1368 5724 1420
rect 5776 1408 5782 1420
rect 9490 1408 9496 1420
rect 5776 1380 9496 1408
rect 5776 1368 5782 1380
rect 9490 1368 9496 1380
rect 9548 1368 9554 1420
rect 26142 1368 26148 1420
rect 26200 1408 26206 1420
rect 28258 1408 28264 1420
rect 26200 1380 28264 1408
rect 26200 1368 26206 1380
rect 28258 1368 28264 1380
rect 28316 1368 28322 1420
rect 35986 1368 35992 1420
rect 36044 1408 36050 1420
rect 37458 1408 37464 1420
rect 36044 1380 37464 1408
rect 36044 1368 36050 1380
rect 37458 1368 37464 1380
rect 37516 1368 37522 1420
rect 36814 1300 36820 1352
rect 36872 1340 36878 1352
rect 37826 1340 37832 1352
rect 36872 1312 37832 1340
rect 36872 1300 36878 1312
rect 37826 1300 37832 1312
rect 37884 1300 37890 1352
rect 46934 1300 46940 1352
rect 46992 1340 46998 1352
rect 55950 1340 55956 1352
rect 46992 1312 55956 1340
rect 46992 1300 46998 1312
rect 55950 1300 55956 1312
rect 56008 1300 56014 1352
rect 35434 1164 35440 1216
rect 35492 1204 35498 1216
rect 38562 1204 38568 1216
rect 35492 1176 38568 1204
rect 35492 1164 35498 1176
rect 38562 1164 38568 1176
rect 38620 1164 38626 1216
rect 39022 1028 39028 1080
rect 39080 1068 39086 1080
rect 45186 1068 45192 1080
rect 39080 1040 45192 1068
rect 39080 1028 39086 1040
rect 45186 1028 45192 1040
rect 45244 1028 45250 1080
<< via1 >>
rect 30104 61752 30156 61804
rect 49424 61752 49476 61804
rect 33416 61684 33468 61736
rect 42708 61684 42760 61736
rect 11060 61616 11112 61668
rect 19432 61616 19484 61668
rect 28448 61616 28500 61668
rect 46848 61616 46900 61668
rect 21180 61548 21232 61600
rect 40224 61548 40276 61600
rect 41880 61548 41932 61600
rect 51448 61548 51500 61600
rect 4214 61446 4266 61498
rect 4278 61446 4330 61498
rect 4342 61446 4394 61498
rect 4406 61446 4458 61498
rect 4470 61446 4522 61498
rect 34934 61446 34986 61498
rect 34998 61446 35050 61498
rect 35062 61446 35114 61498
rect 35126 61446 35178 61498
rect 35190 61446 35242 61498
rect 7656 61344 7708 61396
rect 40224 61387 40276 61396
rect 15844 61276 15896 61328
rect 1676 61183 1728 61192
rect 1676 61149 1685 61183
rect 1685 61149 1719 61183
rect 1719 61149 1728 61183
rect 1676 61140 1728 61149
rect 2780 61183 2832 61192
rect 2780 61149 2789 61183
rect 2789 61149 2823 61183
rect 2823 61149 2832 61183
rect 2780 61140 2832 61149
rect 4620 61140 4672 61192
rect 5080 61183 5132 61192
rect 5080 61149 5089 61183
rect 5089 61149 5123 61183
rect 5123 61149 5132 61183
rect 5080 61140 5132 61149
rect 5724 61183 5776 61192
rect 5724 61149 5733 61183
rect 5733 61149 5767 61183
rect 5767 61149 5776 61183
rect 5724 61140 5776 61149
rect 6644 61183 6696 61192
rect 6644 61149 6653 61183
rect 6653 61149 6687 61183
rect 6687 61149 6696 61183
rect 6644 61140 6696 61149
rect 7564 61183 7616 61192
rect 7564 61149 7573 61183
rect 7573 61149 7607 61183
rect 7607 61149 7616 61183
rect 7564 61140 7616 61149
rect 9680 61140 9732 61192
rect 10232 61183 10284 61192
rect 10232 61149 10241 61183
rect 10241 61149 10275 61183
rect 10275 61149 10284 61183
rect 10232 61140 10284 61149
rect 5632 61072 5684 61124
rect 6920 61115 6972 61124
rect 6920 61081 6929 61115
rect 6929 61081 6963 61115
rect 6963 61081 6972 61115
rect 6920 61072 6972 61081
rect 8944 61072 8996 61124
rect 18236 61276 18288 61328
rect 22100 61276 22152 61328
rect 22836 61208 22888 61260
rect 40224 61353 40233 61387
rect 40233 61353 40267 61387
rect 40267 61353 40276 61387
rect 40224 61344 40276 61353
rect 42616 61344 42668 61396
rect 46848 61387 46900 61396
rect 46848 61353 46857 61387
rect 46857 61353 46891 61387
rect 46891 61353 46900 61387
rect 46848 61344 46900 61353
rect 49424 61387 49476 61396
rect 49424 61353 49433 61387
rect 49433 61353 49467 61387
rect 49467 61353 49476 61387
rect 49424 61344 49476 61353
rect 51448 61387 51500 61396
rect 51448 61353 51457 61387
rect 51457 61353 51491 61387
rect 51491 61353 51500 61387
rect 51448 61344 51500 61353
rect 11152 61140 11204 61192
rect 11980 61183 12032 61192
rect 11980 61149 11989 61183
rect 11989 61149 12023 61183
rect 12023 61149 12032 61183
rect 11980 61140 12032 61149
rect 12716 61183 12768 61192
rect 12716 61149 12725 61183
rect 12725 61149 12759 61183
rect 12759 61149 12768 61183
rect 12716 61140 12768 61149
rect 12992 61183 13044 61192
rect 12992 61149 13001 61183
rect 13001 61149 13035 61183
rect 13035 61149 13044 61183
rect 12992 61140 13044 61149
rect 14924 61183 14976 61192
rect 14924 61149 14933 61183
rect 14933 61149 14967 61183
rect 14967 61149 14976 61183
rect 14924 61140 14976 61149
rect 16120 61183 16172 61192
rect 16120 61149 16129 61183
rect 16129 61149 16163 61183
rect 16163 61149 16172 61183
rect 16120 61140 16172 61149
rect 17224 61183 17276 61192
rect 17224 61149 17233 61183
rect 17233 61149 17267 61183
rect 17267 61149 17276 61183
rect 17224 61140 17276 61149
rect 17960 61183 18012 61192
rect 17960 61149 17969 61183
rect 17969 61149 18003 61183
rect 18003 61149 18012 61183
rect 17960 61140 18012 61149
rect 18696 61183 18748 61192
rect 18696 61149 18705 61183
rect 18705 61149 18739 61183
rect 18739 61149 18748 61183
rect 18696 61140 18748 61149
rect 19800 61183 19852 61192
rect 19800 61149 19809 61183
rect 19809 61149 19843 61183
rect 19843 61149 19852 61183
rect 19800 61140 19852 61149
rect 20720 61140 20772 61192
rect 21272 61183 21324 61192
rect 21272 61149 21281 61183
rect 21281 61149 21315 61183
rect 21315 61149 21324 61183
rect 21272 61140 21324 61149
rect 22376 61183 22428 61192
rect 22376 61149 22385 61183
rect 22385 61149 22419 61183
rect 22419 61149 22428 61183
rect 22376 61140 22428 61149
rect 35900 61208 35952 61260
rect 23848 61183 23900 61192
rect 14648 61072 14700 61124
rect 15200 61115 15252 61124
rect 15200 61081 15209 61115
rect 15209 61081 15243 61115
rect 15243 61081 15252 61115
rect 15200 61072 15252 61081
rect 17408 61072 17460 61124
rect 18880 61115 18932 61124
rect 18880 61081 18889 61115
rect 18889 61081 18923 61115
rect 18923 61081 18932 61115
rect 18880 61072 18932 61081
rect 20444 61072 20496 61124
rect 21088 61072 21140 61124
rect 23848 61149 23857 61183
rect 23857 61149 23891 61183
rect 23891 61149 23900 61183
rect 23848 61140 23900 61149
rect 25136 61140 25188 61192
rect 26240 61183 26292 61192
rect 26240 61149 26249 61183
rect 26249 61149 26283 61183
rect 26283 61149 26292 61183
rect 26240 61140 26292 61149
rect 26608 61140 26660 61192
rect 28080 61140 28132 61192
rect 29828 61183 29880 61192
rect 29828 61149 29837 61183
rect 29837 61149 29871 61183
rect 29871 61149 29880 61183
rect 29828 61140 29880 61149
rect 31208 61183 31260 61192
rect 31208 61149 31217 61183
rect 31217 61149 31251 61183
rect 31251 61149 31260 61183
rect 31208 61140 31260 61149
rect 31760 61140 31812 61192
rect 32864 61140 32916 61192
rect 33508 61140 33560 61192
rect 34704 61140 34756 61192
rect 41512 61208 41564 61260
rect 53380 61251 53432 61260
rect 53380 61217 53389 61251
rect 53389 61217 53423 61251
rect 53423 61217 53432 61251
rect 53380 61208 53432 61217
rect 37280 61140 37332 61192
rect 37648 61140 37700 61192
rect 38660 61140 38712 61192
rect 39488 61140 39540 61192
rect 40592 61140 40644 61192
rect 42064 61140 42116 61192
rect 42800 61140 42852 61192
rect 43628 61140 43680 61192
rect 44548 61140 44600 61192
rect 45560 61140 45612 61192
rect 46112 61140 46164 61192
rect 47216 61140 47268 61192
rect 48320 61140 48372 61192
rect 48688 61140 48740 61192
rect 49700 61140 49752 61192
rect 51080 61140 51132 61192
rect 51632 61140 51684 61192
rect 53196 61183 53248 61192
rect 53196 61149 53205 61183
rect 53205 61149 53239 61183
rect 53239 61149 53248 61183
rect 53196 61140 53248 61149
rect 54116 61183 54168 61192
rect 54116 61149 54125 61183
rect 54125 61149 54159 61183
rect 54159 61149 54168 61183
rect 54116 61140 54168 61149
rect 55496 61183 55548 61192
rect 55496 61149 55505 61183
rect 55505 61149 55539 61183
rect 55539 61149 55548 61183
rect 55496 61140 55548 61149
rect 56048 61140 56100 61192
rect 57520 61140 57572 61192
rect 22744 61115 22796 61124
rect 22744 61081 22753 61115
rect 22753 61081 22787 61115
rect 22787 61081 22796 61115
rect 22744 61072 22796 61081
rect 24768 61072 24820 61124
rect 28172 61072 28224 61124
rect 33140 61072 33192 61124
rect 34520 61072 34572 61124
rect 35900 61115 35952 61124
rect 35900 61081 35909 61115
rect 35909 61081 35943 61115
rect 35943 61081 35952 61115
rect 35900 61072 35952 61081
rect 38016 61072 38068 61124
rect 39948 61072 40000 61124
rect 42892 61115 42944 61124
rect 42892 61081 42901 61115
rect 42901 61081 42935 61115
rect 42935 61081 42944 61115
rect 42892 61072 42944 61081
rect 55772 61115 55824 61124
rect 4712 61004 4764 61056
rect 5172 61047 5224 61056
rect 5172 61013 5181 61047
rect 5181 61013 5215 61047
rect 5215 61013 5224 61047
rect 5172 61004 5224 61013
rect 5908 61047 5960 61056
rect 5908 61013 5917 61047
rect 5917 61013 5951 61047
rect 5951 61013 5960 61047
rect 5908 61004 5960 61013
rect 11060 61047 11112 61056
rect 11060 61013 11069 61047
rect 11069 61013 11103 61047
rect 11103 61013 11112 61047
rect 11060 61004 11112 61013
rect 12164 61047 12216 61056
rect 12164 61013 12173 61047
rect 12173 61013 12207 61047
rect 12207 61013 12216 61047
rect 12164 61004 12216 61013
rect 17316 61047 17368 61056
rect 17316 61013 17325 61047
rect 17325 61013 17359 61047
rect 17359 61013 17368 61047
rect 17316 61004 17368 61013
rect 20904 61004 20956 61056
rect 25412 61047 25464 61056
rect 25412 61013 25421 61047
rect 25421 61013 25455 61047
rect 25455 61013 25464 61047
rect 25412 61004 25464 61013
rect 27344 61047 27396 61056
rect 27344 61013 27353 61047
rect 27353 61013 27387 61047
rect 27387 61013 27396 61047
rect 27344 61004 27396 61013
rect 28356 61047 28408 61056
rect 28356 61013 28365 61047
rect 28365 61013 28399 61047
rect 28399 61013 28408 61047
rect 28356 61004 28408 61013
rect 29920 61047 29972 61056
rect 29920 61013 29929 61047
rect 29929 61013 29963 61047
rect 29963 61013 29972 61047
rect 29920 61004 29972 61013
rect 31300 61047 31352 61056
rect 31300 61013 31309 61047
rect 31309 61013 31343 61047
rect 31343 61013 31352 61047
rect 31300 61004 31352 61013
rect 32588 61004 32640 61056
rect 33416 61047 33468 61056
rect 33416 61013 33425 61047
rect 33425 61013 33459 61047
rect 33459 61013 33468 61047
rect 33416 61004 33468 61013
rect 35072 61047 35124 61056
rect 35072 61013 35081 61047
rect 35081 61013 35115 61047
rect 35115 61013 35124 61047
rect 35072 61004 35124 61013
rect 36084 61004 36136 61056
rect 39120 61047 39172 61056
rect 39120 61013 39129 61047
rect 39129 61013 39163 61047
rect 39163 61013 39172 61047
rect 39120 61004 39172 61013
rect 40316 61004 40368 61056
rect 41696 61047 41748 61056
rect 41696 61013 41705 61047
rect 41705 61013 41739 61047
rect 41739 61013 41748 61047
rect 41696 61004 41748 61013
rect 44456 61047 44508 61056
rect 44456 61013 44465 61047
rect 44465 61013 44499 61047
rect 44499 61013 44508 61047
rect 44456 61004 44508 61013
rect 45376 61047 45428 61056
rect 45376 61013 45385 61047
rect 45385 61013 45419 61047
rect 45419 61013 45428 61047
rect 45376 61004 45428 61013
rect 46112 61047 46164 61056
rect 46112 61013 46121 61047
rect 46121 61013 46155 61047
rect 46155 61013 46164 61047
rect 46112 61004 46164 61013
rect 46848 61004 46900 61056
rect 50068 61004 50120 61056
rect 53196 61004 53248 61056
rect 54300 61047 54352 61056
rect 54300 61013 54309 61047
rect 54309 61013 54343 61047
rect 54343 61013 54352 61047
rect 54300 61004 54352 61013
rect 55772 61081 55781 61115
rect 55781 61081 55815 61115
rect 55815 61081 55824 61115
rect 55772 61072 55824 61081
rect 56692 61004 56744 61056
rect 19574 60902 19626 60954
rect 19638 60902 19690 60954
rect 19702 60902 19754 60954
rect 19766 60902 19818 60954
rect 19830 60902 19882 60954
rect 50294 60902 50346 60954
rect 50358 60902 50410 60954
rect 50422 60902 50474 60954
rect 50486 60902 50538 60954
rect 50550 60902 50602 60954
rect 5172 60800 5224 60852
rect 23480 60800 23532 60852
rect 23756 60800 23808 60852
rect 44456 60800 44508 60852
rect 3240 60775 3292 60784
rect 3240 60741 3249 60775
rect 3249 60741 3283 60775
rect 3283 60741 3292 60775
rect 3240 60732 3292 60741
rect 3976 60775 4028 60784
rect 3976 60741 3985 60775
rect 3985 60741 4019 60775
rect 4019 60741 4028 60775
rect 3976 60732 4028 60741
rect 8300 60732 8352 60784
rect 13544 60775 13596 60784
rect 13544 60741 13553 60775
rect 13553 60741 13587 60775
rect 13587 60741 13596 60775
rect 13544 60732 13596 60741
rect 14280 60775 14332 60784
rect 14280 60741 14289 60775
rect 14289 60741 14323 60775
rect 14323 60741 14332 60775
rect 14280 60732 14332 60741
rect 15752 60775 15804 60784
rect 15752 60741 15761 60775
rect 15761 60741 15795 60775
rect 15795 60741 15804 60775
rect 15752 60732 15804 60741
rect 15844 60732 15896 60784
rect 1584 60707 1636 60716
rect 1584 60673 1593 60707
rect 1593 60673 1627 60707
rect 1627 60673 1636 60707
rect 1584 60664 1636 60673
rect 9036 60707 9088 60716
rect 9036 60673 9045 60707
rect 9045 60673 9079 60707
rect 9079 60673 9088 60707
rect 9036 60664 9088 60673
rect 19340 60732 19392 60784
rect 23296 60732 23348 60784
rect 24400 60732 24452 60784
rect 27528 60775 27580 60784
rect 27528 60741 27537 60775
rect 27537 60741 27571 60775
rect 27571 60741 27580 60775
rect 27528 60732 27580 60741
rect 28816 60732 28868 60784
rect 30380 60732 30432 60784
rect 36360 60775 36412 60784
rect 36360 60741 36369 60775
rect 36369 60741 36403 60775
rect 36403 60741 36412 60775
rect 36360 60732 36412 60741
rect 41420 60732 41472 60784
rect 46664 60775 46716 60784
rect 46664 60741 46673 60775
rect 46673 60741 46707 60775
rect 46707 60741 46716 60775
rect 46664 60732 46716 60741
rect 50160 60732 50212 60784
rect 52460 60732 52512 60784
rect 22100 60707 22152 60716
rect 22100 60673 22109 60707
rect 22109 60673 22143 60707
rect 22143 60673 22152 60707
rect 22100 60664 22152 60673
rect 22560 60707 22612 60716
rect 22560 60673 22563 60707
rect 22563 60673 22612 60707
rect 5540 60596 5592 60648
rect 4620 60528 4672 60580
rect 18420 60528 18472 60580
rect 20628 60528 20680 60580
rect 3332 60503 3384 60512
rect 3332 60469 3341 60503
rect 3341 60469 3375 60503
rect 3375 60469 3384 60503
rect 3332 60460 3384 60469
rect 9220 60503 9272 60512
rect 9220 60469 9229 60503
rect 9229 60469 9263 60503
rect 9263 60469 9272 60503
rect 9220 60460 9272 60469
rect 13636 60503 13688 60512
rect 13636 60469 13645 60503
rect 13645 60469 13679 60503
rect 13679 60469 13688 60503
rect 13636 60460 13688 60469
rect 14372 60503 14424 60512
rect 14372 60469 14381 60503
rect 14381 60469 14415 60503
rect 14415 60469 14424 60503
rect 14372 60460 14424 60469
rect 17868 60460 17920 60512
rect 20536 60460 20588 60512
rect 22560 60664 22612 60673
rect 23204 60707 23256 60716
rect 23204 60673 23213 60707
rect 23213 60673 23247 60707
rect 23247 60673 23256 60707
rect 23204 60664 23256 60673
rect 54668 60707 54720 60716
rect 54668 60673 54677 60707
rect 54677 60673 54711 60707
rect 54711 60673 54720 60707
rect 54668 60664 54720 60673
rect 55404 60707 55456 60716
rect 55404 60673 55413 60707
rect 55413 60673 55447 60707
rect 55447 60673 55456 60707
rect 55404 60664 55456 60673
rect 56140 60707 56192 60716
rect 56140 60673 56149 60707
rect 56149 60673 56183 60707
rect 56183 60673 56192 60707
rect 56140 60664 56192 60673
rect 56876 60707 56928 60716
rect 56876 60673 56885 60707
rect 56885 60673 56919 60707
rect 56919 60673 56928 60707
rect 56876 60664 56928 60673
rect 58072 60707 58124 60716
rect 58072 60673 58081 60707
rect 58081 60673 58115 60707
rect 58115 60673 58124 60707
rect 58072 60664 58124 60673
rect 40776 60596 40828 60648
rect 22468 60460 22520 60512
rect 22928 60460 22980 60512
rect 23388 60503 23440 60512
rect 23388 60469 23397 60503
rect 23397 60469 23431 60503
rect 23431 60469 23440 60503
rect 23388 60460 23440 60469
rect 25228 60460 25280 60512
rect 29000 60460 29052 60512
rect 29828 60460 29880 60512
rect 30564 60503 30616 60512
rect 30564 60469 30573 60503
rect 30573 60469 30607 60503
rect 30607 60469 30616 60503
rect 30564 60460 30616 60469
rect 33048 60460 33100 60512
rect 35072 60460 35124 60512
rect 35716 60460 35768 60512
rect 40868 60460 40920 60512
rect 44180 60460 44232 60512
rect 50436 60503 50488 60512
rect 50436 60469 50445 60503
rect 50445 60469 50479 60503
rect 50479 60469 50488 60503
rect 50436 60460 50488 60469
rect 53104 60503 53156 60512
rect 53104 60469 53113 60503
rect 53113 60469 53147 60503
rect 53147 60469 53156 60503
rect 53104 60460 53156 60469
rect 54852 60503 54904 60512
rect 54852 60469 54861 60503
rect 54861 60469 54895 60503
rect 54895 60469 54904 60503
rect 54852 60460 54904 60469
rect 55588 60503 55640 60512
rect 55588 60469 55597 60503
rect 55597 60469 55631 60503
rect 55631 60469 55640 60503
rect 55588 60460 55640 60469
rect 57060 60503 57112 60512
rect 57060 60469 57069 60503
rect 57069 60469 57103 60503
rect 57103 60469 57112 60503
rect 57060 60460 57112 60469
rect 58256 60503 58308 60512
rect 58256 60469 58265 60503
rect 58265 60469 58299 60503
rect 58299 60469 58308 60503
rect 58256 60460 58308 60469
rect 4214 60358 4266 60410
rect 4278 60358 4330 60410
rect 4342 60358 4394 60410
rect 4406 60358 4458 60410
rect 4470 60358 4522 60410
rect 34934 60358 34986 60410
rect 34998 60358 35050 60410
rect 35062 60358 35114 60410
rect 35126 60358 35178 60410
rect 35190 60358 35242 60410
rect 3332 60256 3384 60308
rect 20260 60256 20312 60308
rect 20720 60256 20772 60308
rect 55588 60256 55640 60308
rect 13636 60188 13688 60240
rect 17868 60163 17920 60172
rect 2596 60095 2648 60104
rect 2596 60061 2605 60095
rect 2605 60061 2639 60095
rect 2639 60061 2648 60095
rect 2596 60052 2648 60061
rect 5632 60052 5684 60104
rect 7656 60095 7708 60104
rect 7656 60061 7665 60095
rect 7665 60061 7699 60095
rect 7699 60061 7708 60095
rect 7656 60052 7708 60061
rect 1676 60027 1728 60036
rect 1676 59993 1685 60027
rect 1685 59993 1719 60027
rect 1719 59993 1728 60027
rect 1676 59984 1728 59993
rect 2044 60027 2096 60036
rect 2044 59993 2053 60027
rect 2053 59993 2087 60027
rect 2087 59993 2096 60027
rect 2044 59984 2096 59993
rect 2504 59916 2556 59968
rect 17592 59984 17644 60036
rect 8024 59916 8076 59968
rect 17500 59959 17552 59968
rect 17500 59925 17509 59959
rect 17509 59925 17543 59959
rect 17543 59925 17552 59959
rect 17500 59916 17552 59925
rect 17868 60129 17877 60163
rect 17877 60129 17911 60163
rect 17911 60129 17920 60163
rect 17868 60120 17920 60129
rect 21364 60188 21416 60240
rect 22652 60188 22704 60240
rect 23388 60188 23440 60240
rect 26884 60120 26936 60172
rect 30196 60188 30248 60240
rect 41144 60231 41196 60240
rect 18420 60095 18472 60104
rect 18420 60061 18429 60095
rect 18429 60061 18463 60095
rect 18463 60061 18472 60095
rect 18420 60052 18472 60061
rect 18604 60095 18656 60104
rect 18604 60061 18613 60095
rect 18613 60061 18647 60095
rect 18647 60061 18656 60095
rect 18604 60052 18656 60061
rect 19984 60052 20036 60104
rect 20444 60095 20496 60104
rect 20444 60061 20453 60095
rect 20453 60061 20487 60095
rect 20487 60061 20496 60095
rect 20444 60052 20496 60061
rect 20536 60052 20588 60104
rect 20720 60095 20772 60104
rect 20720 60061 20729 60095
rect 20729 60061 20763 60095
rect 20763 60061 20772 60095
rect 20720 60052 20772 60061
rect 21824 60052 21876 60104
rect 22008 60095 22060 60104
rect 22008 60061 22017 60095
rect 22017 60061 22051 60095
rect 22051 60061 22060 60095
rect 22008 60052 22060 60061
rect 22100 60095 22152 60104
rect 22100 60061 22109 60095
rect 22109 60061 22143 60095
rect 22143 60061 22152 60095
rect 22376 60095 22428 60104
rect 22100 60052 22152 60061
rect 22376 60061 22385 60095
rect 22385 60061 22419 60095
rect 22419 60061 22428 60095
rect 22376 60052 22428 60061
rect 22468 60052 22520 60104
rect 22836 60095 22888 60104
rect 19248 59984 19300 60036
rect 21272 59984 21324 60036
rect 22836 60061 22845 60095
rect 22845 60061 22879 60095
rect 22879 60061 22888 60095
rect 22836 60052 22888 60061
rect 23480 60095 23532 60104
rect 23480 60061 23489 60095
rect 23489 60061 23523 60095
rect 23523 60061 23532 60095
rect 23480 60052 23532 60061
rect 23756 60095 23808 60104
rect 23756 60061 23765 60095
rect 23765 60061 23799 60095
rect 23799 60061 23808 60095
rect 23756 60052 23808 60061
rect 23940 60052 23992 60104
rect 28080 60095 28132 60104
rect 28080 60061 28089 60095
rect 28089 60061 28123 60095
rect 28123 60061 28132 60095
rect 28080 60052 28132 60061
rect 28172 60095 28224 60104
rect 28172 60061 28182 60095
rect 28182 60061 28216 60095
rect 28216 60061 28224 60095
rect 28448 60095 28500 60104
rect 28172 60052 28224 60061
rect 28448 60061 28457 60095
rect 28457 60061 28491 60095
rect 28491 60061 28500 60095
rect 28448 60052 28500 60061
rect 29000 60120 29052 60172
rect 30380 60095 30432 60104
rect 30380 60061 30389 60095
rect 30389 60061 30423 60095
rect 30423 60061 30432 60095
rect 30380 60052 30432 60061
rect 41144 60197 41153 60231
rect 41153 60197 41187 60231
rect 41187 60197 41196 60231
rect 41144 60188 41196 60197
rect 32496 60095 32548 60104
rect 32496 60061 32505 60095
rect 32505 60061 32539 60095
rect 32539 60061 32548 60095
rect 32496 60052 32548 60061
rect 32680 60095 32732 60104
rect 32680 60061 32689 60095
rect 32689 60061 32723 60095
rect 32723 60061 32732 60095
rect 32680 60052 32732 60061
rect 33048 60095 33100 60104
rect 33048 60061 33057 60095
rect 33057 60061 33091 60095
rect 33091 60061 33100 60095
rect 33048 60052 33100 60061
rect 34520 60052 34572 60104
rect 21640 59959 21692 59968
rect 21640 59925 21649 59959
rect 21649 59925 21683 59959
rect 21683 59925 21692 59959
rect 21640 59916 21692 59925
rect 23572 59984 23624 60036
rect 30012 59984 30064 60036
rect 30656 60027 30708 60036
rect 30656 59993 30665 60027
rect 30665 59993 30699 60027
rect 30699 59993 30708 60027
rect 30656 59984 30708 59993
rect 41512 60120 41564 60172
rect 40592 60095 40644 60104
rect 40592 60061 40601 60095
rect 40601 60061 40635 60095
rect 40635 60061 40644 60095
rect 40592 60052 40644 60061
rect 40868 60095 40920 60104
rect 40868 60061 40877 60095
rect 40877 60061 40911 60095
rect 40911 60061 40920 60095
rect 40868 60052 40920 60061
rect 40960 60095 41012 60104
rect 40960 60061 40974 60095
rect 40974 60061 41008 60095
rect 41008 60061 41012 60095
rect 42156 60095 42208 60104
rect 40960 60052 41012 60061
rect 42156 60061 42165 60095
rect 42165 60061 42199 60095
rect 42199 60061 42208 60095
rect 42156 60052 42208 60061
rect 42340 60095 42392 60104
rect 42340 60061 42349 60095
rect 42349 60061 42383 60095
rect 42383 60061 42392 60095
rect 42340 60052 42392 60061
rect 40776 60027 40828 60036
rect 40776 59993 40785 60027
rect 40785 59993 40819 60027
rect 40819 59993 40828 60027
rect 40776 59984 40828 59993
rect 50436 60188 50488 60240
rect 53932 60120 53984 60172
rect 56508 60095 56560 60104
rect 56508 60061 56517 60095
rect 56517 60061 56551 60095
rect 56551 60061 56560 60095
rect 56508 60052 56560 60061
rect 57244 60095 57296 60104
rect 57244 60061 57253 60095
rect 57253 60061 57287 60095
rect 57287 60061 57296 60095
rect 57244 60052 57296 60061
rect 57980 60052 58032 60104
rect 43536 59984 43588 60036
rect 58256 59984 58308 60036
rect 24400 59916 24452 59968
rect 28540 59916 28592 59968
rect 28724 59959 28776 59968
rect 28724 59925 28733 59959
rect 28733 59925 28767 59959
rect 28767 59925 28776 59959
rect 28724 59916 28776 59925
rect 31024 59959 31076 59968
rect 31024 59925 31033 59959
rect 31033 59925 31067 59959
rect 31067 59925 31076 59959
rect 31024 59916 31076 59925
rect 32312 59959 32364 59968
rect 32312 59925 32321 59959
rect 32321 59925 32355 59959
rect 32355 59925 32364 59959
rect 32312 59916 32364 59925
rect 41972 59959 42024 59968
rect 41972 59925 41981 59959
rect 41981 59925 42015 59959
rect 42015 59925 42024 59959
rect 41972 59916 42024 59925
rect 54116 59916 54168 59968
rect 19574 59814 19626 59866
rect 19638 59814 19690 59866
rect 19702 59814 19754 59866
rect 19766 59814 19818 59866
rect 19830 59814 19882 59866
rect 50294 59814 50346 59866
rect 50358 59814 50410 59866
rect 50422 59814 50474 59866
rect 50486 59814 50538 59866
rect 50550 59814 50602 59866
rect 14372 59712 14424 59764
rect 32496 59712 32548 59764
rect 32680 59712 32732 59764
rect 33048 59712 33100 59764
rect 42340 59712 42392 59764
rect 1768 59644 1820 59696
rect 18236 59644 18288 59696
rect 1676 59619 1728 59628
rect 1676 59585 1685 59619
rect 1685 59585 1719 59619
rect 1719 59585 1728 59619
rect 1676 59576 1728 59585
rect 17960 59576 18012 59628
rect 17592 59508 17644 59560
rect 19248 59508 19300 59560
rect 1952 59415 2004 59424
rect 1952 59381 1961 59415
rect 1961 59381 1995 59415
rect 1995 59381 2004 59415
rect 1952 59372 2004 59381
rect 2320 59372 2372 59424
rect 19984 59576 20036 59628
rect 21456 59644 21508 59696
rect 23388 59687 23440 59696
rect 21088 59619 21140 59628
rect 21088 59585 21097 59619
rect 21097 59585 21131 59619
rect 21131 59585 21140 59619
rect 21088 59576 21140 59585
rect 22100 59619 22152 59628
rect 22100 59585 22109 59619
rect 22109 59585 22143 59619
rect 22143 59585 22152 59619
rect 22100 59576 22152 59585
rect 22744 59576 22796 59628
rect 20168 59372 20220 59424
rect 22376 59440 22428 59492
rect 23388 59653 23397 59687
rect 23397 59653 23431 59687
rect 23431 59653 23440 59687
rect 23388 59644 23440 59653
rect 30104 59687 30156 59696
rect 30104 59653 30113 59687
rect 30113 59653 30147 59687
rect 30147 59653 30156 59687
rect 30104 59644 30156 59653
rect 23296 59576 23348 59628
rect 23664 59619 23716 59628
rect 23664 59585 23667 59619
rect 23667 59585 23716 59619
rect 23664 59576 23716 59585
rect 28448 59576 28500 59628
rect 29736 59619 29788 59628
rect 29736 59585 29745 59619
rect 29745 59585 29779 59619
rect 29779 59585 29788 59619
rect 29736 59576 29788 59585
rect 29828 59619 29880 59628
rect 29828 59585 29838 59619
rect 29838 59585 29872 59619
rect 29872 59585 29880 59619
rect 29828 59576 29880 59585
rect 30012 59619 30064 59628
rect 30012 59585 30021 59619
rect 30021 59585 30055 59619
rect 30055 59585 30064 59619
rect 30012 59576 30064 59585
rect 30196 59619 30248 59628
rect 30196 59585 30210 59619
rect 30210 59585 30244 59619
rect 30244 59585 30248 59619
rect 30196 59576 30248 59585
rect 28540 59551 28592 59560
rect 23480 59440 23532 59492
rect 28540 59517 28549 59551
rect 28549 59517 28583 59551
rect 28583 59517 28592 59551
rect 28540 59508 28592 59517
rect 28632 59508 28684 59560
rect 30104 59508 30156 59560
rect 56416 59644 56468 59696
rect 30564 59576 30616 59628
rect 42156 59576 42208 59628
rect 42340 59576 42392 59628
rect 53104 59576 53156 59628
rect 58072 59619 58124 59628
rect 58072 59585 58081 59619
rect 58081 59585 58115 59619
rect 58115 59585 58124 59619
rect 58072 59576 58124 59585
rect 30656 59508 30708 59560
rect 42708 59551 42760 59560
rect 42708 59517 42717 59551
rect 42717 59517 42751 59551
rect 42751 59517 42760 59551
rect 42708 59508 42760 59517
rect 42800 59508 42852 59560
rect 43536 59551 43588 59560
rect 43536 59517 43545 59551
rect 43545 59517 43579 59551
rect 43579 59517 43588 59551
rect 43536 59508 43588 59517
rect 21180 59372 21232 59424
rect 21456 59372 21508 59424
rect 23664 59372 23716 59424
rect 24492 59372 24544 59424
rect 29736 59372 29788 59424
rect 30288 59372 30340 59424
rect 30564 59440 30616 59492
rect 32956 59440 33008 59492
rect 40592 59440 40644 59492
rect 30472 59372 30524 59424
rect 31576 59372 31628 59424
rect 57152 59372 57204 59424
rect 58992 59372 59044 59424
rect 4214 59270 4266 59322
rect 4278 59270 4330 59322
rect 4342 59270 4394 59322
rect 4406 59270 4458 59322
rect 4470 59270 4522 59322
rect 34934 59270 34986 59322
rect 34998 59270 35050 59322
rect 35062 59270 35114 59322
rect 35126 59270 35178 59322
rect 35190 59270 35242 59322
rect 1952 59032 2004 59084
rect 848 58964 900 59016
rect 19524 59100 19576 59152
rect 41788 59075 41840 59084
rect 41788 59041 41797 59075
rect 41797 59041 41831 59075
rect 41831 59041 41840 59075
rect 41788 59032 41840 59041
rect 58072 59075 58124 59084
rect 58072 59041 58081 59075
rect 58081 59041 58115 59075
rect 58115 59041 58124 59075
rect 58072 59032 58124 59041
rect 19708 59007 19760 59016
rect 19708 58973 19717 59007
rect 19717 58973 19751 59007
rect 19751 58973 19760 59007
rect 19708 58964 19760 58973
rect 21456 58964 21508 59016
rect 41236 58964 41288 59016
rect 41880 59007 41932 59016
rect 41880 58973 41889 59007
rect 41889 58973 41923 59007
rect 41923 58973 41932 59007
rect 41880 58964 41932 58973
rect 57152 59007 57204 59016
rect 57152 58973 57161 59007
rect 57161 58973 57195 59007
rect 57195 58973 57204 59007
rect 57152 58964 57204 58973
rect 57888 59007 57940 59016
rect 57888 58973 57897 59007
rect 57897 58973 57931 59007
rect 57931 58973 57940 59007
rect 57888 58964 57940 58973
rect 17960 58828 18012 58880
rect 19984 58828 20036 58880
rect 42340 58828 42392 58880
rect 19574 58726 19626 58778
rect 19638 58726 19690 58778
rect 19702 58726 19754 58778
rect 19766 58726 19818 58778
rect 19830 58726 19882 58778
rect 50294 58726 50346 58778
rect 50358 58726 50410 58778
rect 50422 58726 50474 58778
rect 50486 58726 50538 58778
rect 50550 58726 50602 58778
rect 2044 58624 2096 58676
rect 1584 58531 1636 58540
rect 1584 58497 1593 58531
rect 1593 58497 1627 58531
rect 1627 58497 1636 58531
rect 1584 58488 1636 58497
rect 37924 58531 37976 58540
rect 37924 58497 37933 58531
rect 37933 58497 37967 58531
rect 37967 58497 37976 58531
rect 37924 58488 37976 58497
rect 38016 58531 38068 58540
rect 38016 58497 38025 58531
rect 38025 58497 38059 58531
rect 38059 58497 38068 58531
rect 38016 58488 38068 58497
rect 4804 58420 4856 58472
rect 36912 58420 36964 58472
rect 37188 58352 37240 58404
rect 58164 58599 58216 58608
rect 41512 58531 41564 58540
rect 41512 58497 41521 58531
rect 41521 58497 41555 58531
rect 41555 58497 41564 58531
rect 41512 58488 41564 58497
rect 42616 58488 42668 58540
rect 58164 58565 58173 58599
rect 58173 58565 58207 58599
rect 58207 58565 58216 58599
rect 58164 58556 58216 58565
rect 56692 58488 56744 58540
rect 37556 58327 37608 58336
rect 37556 58293 37565 58327
rect 37565 58293 37599 58327
rect 37599 58293 37608 58327
rect 37556 58284 37608 58293
rect 37924 58284 37976 58336
rect 40960 58420 41012 58472
rect 41788 58463 41840 58472
rect 41788 58429 41797 58463
rect 41797 58429 41831 58463
rect 41831 58429 41840 58463
rect 41788 58420 41840 58429
rect 41328 58284 41380 58336
rect 52460 58284 52512 58336
rect 4214 58182 4266 58234
rect 4278 58182 4330 58234
rect 4342 58182 4394 58234
rect 4406 58182 4458 58234
rect 4470 58182 4522 58234
rect 34934 58182 34986 58234
rect 34998 58182 35050 58234
rect 35062 58182 35114 58234
rect 35126 58182 35178 58234
rect 35190 58182 35242 58234
rect 35348 58080 35400 58132
rect 41512 58080 41564 58132
rect 1584 57919 1636 57928
rect 1584 57885 1593 57919
rect 1593 57885 1627 57919
rect 1627 57885 1636 57919
rect 1584 57876 1636 57885
rect 35624 57919 35676 57928
rect 35624 57885 35633 57919
rect 35633 57885 35667 57919
rect 35667 57885 35676 57919
rect 35624 57876 35676 57885
rect 10140 57808 10192 57860
rect 34704 57808 34756 57860
rect 35716 57740 35768 57792
rect 35992 57919 36044 57928
rect 35992 57885 36001 57919
rect 36001 57885 36035 57919
rect 36035 57885 36044 57919
rect 36268 57919 36320 57928
rect 35992 57876 36044 57885
rect 36268 57885 36277 57919
rect 36277 57885 36311 57919
rect 36311 57885 36320 57919
rect 36268 57876 36320 57885
rect 52460 57876 52512 57928
rect 57980 57851 58032 57860
rect 57980 57817 57989 57851
rect 57989 57817 58023 57851
rect 58023 57817 58032 57851
rect 57980 57808 58032 57817
rect 58072 57783 58124 57792
rect 58072 57749 58081 57783
rect 58081 57749 58115 57783
rect 58115 57749 58124 57783
rect 58072 57740 58124 57749
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 34612 57468 34664 57520
rect 35992 57468 36044 57520
rect 1584 57443 1636 57452
rect 1584 57409 1593 57443
rect 1593 57409 1627 57443
rect 1627 57409 1636 57443
rect 1584 57400 1636 57409
rect 34520 57400 34572 57452
rect 35624 57332 35676 57384
rect 37924 57332 37976 57384
rect 4712 57264 4764 57316
rect 15936 57264 15988 57316
rect 1768 57239 1820 57248
rect 1768 57205 1777 57239
rect 1777 57205 1811 57239
rect 1811 57205 1820 57239
rect 1768 57196 1820 57205
rect 5540 57196 5592 57248
rect 31484 57196 31536 57248
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 29368 56992 29420 57044
rect 30656 56992 30708 57044
rect 17040 56856 17092 56908
rect 22100 56856 22152 56908
rect 26884 56856 26936 56908
rect 32956 56856 33008 56908
rect 33048 56831 33100 56840
rect 33048 56797 33057 56831
rect 33057 56797 33091 56831
rect 33091 56797 33100 56831
rect 33048 56788 33100 56797
rect 1676 56763 1728 56772
rect 1676 56729 1685 56763
rect 1685 56729 1719 56763
rect 1719 56729 1728 56763
rect 1676 56720 1728 56729
rect 2044 56763 2096 56772
rect 2044 56729 2053 56763
rect 2053 56729 2087 56763
rect 2087 56729 2096 56763
rect 2044 56720 2096 56729
rect 36268 56788 36320 56840
rect 41328 56788 41380 56840
rect 43996 56788 44048 56840
rect 57888 56831 57940 56840
rect 57888 56797 57897 56831
rect 57897 56797 57931 56831
rect 57931 56797 57940 56831
rect 57888 56788 57940 56797
rect 49608 56720 49660 56772
rect 51724 56720 51776 56772
rect 32496 56695 32548 56704
rect 32496 56661 32505 56695
rect 32505 56661 32539 56695
rect 32539 56661 32548 56695
rect 32496 56652 32548 56661
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 1768 56448 1820 56500
rect 2044 56380 2096 56432
rect 23572 56380 23624 56432
rect 24216 56380 24268 56432
rect 24400 56355 24452 56364
rect 24400 56321 24409 56355
rect 24409 56321 24443 56355
rect 24443 56321 24452 56355
rect 24400 56312 24452 56321
rect 24768 56355 24820 56364
rect 24768 56321 24777 56355
rect 24777 56321 24811 56355
rect 24811 56321 24820 56355
rect 24768 56312 24820 56321
rect 25320 56312 25372 56364
rect 24032 56244 24084 56296
rect 29368 56312 29420 56364
rect 41236 56380 41288 56432
rect 58164 56423 58216 56432
rect 58164 56389 58173 56423
rect 58173 56389 58207 56423
rect 58207 56389 58216 56423
rect 58164 56380 58216 56389
rect 29736 56244 29788 56296
rect 46848 56312 46900 56364
rect 40960 56244 41012 56296
rect 23848 56151 23900 56160
rect 23848 56117 23857 56151
rect 23857 56117 23891 56151
rect 23891 56117 23900 56151
rect 23848 56108 23900 56117
rect 29000 56108 29052 56160
rect 41328 56108 41380 56160
rect 49608 56108 49660 56160
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 58348 55947 58400 55956
rect 58348 55913 58357 55947
rect 58357 55913 58391 55947
rect 58391 55913 58400 55947
rect 58348 55904 58400 55913
rect 1768 55836 1820 55888
rect 40868 55836 40920 55888
rect 31024 55768 31076 55820
rect 25320 55743 25372 55752
rect 25320 55709 25329 55743
rect 25329 55709 25363 55743
rect 25363 55709 25372 55743
rect 25320 55700 25372 55709
rect 1676 55675 1728 55684
rect 1676 55641 1685 55675
rect 1685 55641 1719 55675
rect 1719 55641 1728 55675
rect 1676 55632 1728 55641
rect 24308 55632 24360 55684
rect 25688 55743 25740 55752
rect 25688 55709 25697 55743
rect 25697 55709 25731 55743
rect 25731 55709 25740 55743
rect 25688 55700 25740 55709
rect 29736 55700 29788 55752
rect 35348 55632 35400 55684
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 1768 55403 1820 55412
rect 1768 55369 1777 55403
rect 1777 55369 1811 55403
rect 1811 55369 1820 55403
rect 1768 55360 1820 55369
rect 40500 55292 40552 55344
rect 41236 55360 41288 55412
rect 44180 55292 44232 55344
rect 1584 55267 1636 55276
rect 1584 55233 1593 55267
rect 1593 55233 1627 55267
rect 1627 55233 1636 55267
rect 1584 55224 1636 55233
rect 40868 55267 40920 55276
rect 40868 55233 40877 55267
rect 40877 55233 40911 55267
rect 40911 55233 40920 55267
rect 40868 55224 40920 55233
rect 40960 55224 41012 55276
rect 41236 55267 41288 55276
rect 41236 55233 41250 55267
rect 41250 55233 41284 55267
rect 41284 55233 41288 55267
rect 41236 55224 41288 55233
rect 42064 55224 42116 55276
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 24860 54748 24912 54800
rect 25320 54748 25372 54800
rect 28724 54680 28776 54732
rect 1676 54587 1728 54596
rect 1676 54553 1685 54587
rect 1685 54553 1719 54587
rect 1719 54553 1728 54587
rect 1676 54544 1728 54553
rect 22836 54587 22888 54596
rect 22836 54553 22845 54587
rect 22845 54553 22879 54587
rect 22879 54553 22888 54587
rect 22836 54544 22888 54553
rect 25688 54612 25740 54664
rect 58348 54655 58400 54664
rect 58348 54621 58357 54655
rect 58357 54621 58391 54655
rect 58391 54621 58400 54655
rect 58348 54612 58400 54621
rect 28080 54476 28132 54528
rect 39396 54476 39448 54528
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 1584 54179 1636 54188
rect 1584 54145 1593 54179
rect 1593 54145 1627 54179
rect 1627 54145 1636 54179
rect 1584 54136 1636 54145
rect 1768 53975 1820 53984
rect 1768 53941 1777 53975
rect 1777 53941 1811 53975
rect 1811 53941 1820 53975
rect 1768 53932 1820 53941
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 40868 53703 40920 53712
rect 40868 53669 40877 53703
rect 40877 53669 40911 53703
rect 40911 53669 40920 53703
rect 40868 53660 40920 53669
rect 1768 53524 1820 53576
rect 41236 53524 41288 53576
rect 24952 53456 25004 53508
rect 40500 53499 40552 53508
rect 40500 53465 40509 53499
rect 40509 53465 40543 53499
rect 40543 53465 40552 53499
rect 40500 53456 40552 53465
rect 46112 53456 46164 53508
rect 23480 53388 23532 53440
rect 24584 53388 24636 53440
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 24952 53184 25004 53236
rect 45376 53116 45428 53168
rect 1676 53091 1728 53100
rect 1676 53057 1685 53091
rect 1685 53057 1719 53091
rect 1719 53057 1728 53091
rect 1676 53048 1728 53057
rect 23940 53091 23992 53100
rect 23940 53057 23949 53091
rect 23949 53057 23983 53091
rect 23983 53057 23992 53091
rect 23940 53048 23992 53057
rect 24584 53091 24636 53100
rect 24584 53057 24593 53091
rect 24593 53057 24627 53091
rect 24627 53057 24636 53091
rect 24584 53048 24636 53057
rect 23940 52844 23992 52896
rect 58348 52887 58400 52896
rect 58348 52853 58357 52887
rect 58357 52853 58391 52887
rect 58391 52853 58400 52887
rect 58348 52844 58400 52853
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 24952 52683 25004 52692
rect 24952 52649 24961 52683
rect 24961 52649 24995 52683
rect 24995 52649 25004 52683
rect 24952 52640 25004 52649
rect 10784 52504 10836 52556
rect 1584 52479 1636 52488
rect 1584 52445 1593 52479
rect 1593 52445 1627 52479
rect 1627 52445 1636 52479
rect 1584 52436 1636 52445
rect 20720 52368 20772 52420
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 1676 52003 1728 52012
rect 1676 51969 1685 52003
rect 1685 51969 1719 52003
rect 1719 51969 1728 52003
rect 1676 51960 1728 51969
rect 8024 52003 8076 52012
rect 8024 51969 8033 52003
rect 8033 51969 8067 52003
rect 8067 51969 8076 52003
rect 8024 51960 8076 51969
rect 4068 51892 4120 51944
rect 20720 51960 20772 52012
rect 7840 51799 7892 51808
rect 7840 51765 7849 51799
rect 7849 51765 7883 51799
rect 7883 51765 7892 51799
rect 7840 51756 7892 51765
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 24124 51552 24176 51604
rect 17868 51484 17920 51536
rect 41144 51416 41196 51468
rect 1676 51323 1728 51332
rect 1676 51289 1685 51323
rect 1685 51289 1719 51323
rect 1719 51289 1728 51323
rect 1676 51280 1728 51289
rect 3976 51280 4028 51332
rect 20260 51280 20312 51332
rect 21180 51348 21232 51400
rect 58348 51391 58400 51400
rect 58348 51357 58357 51391
rect 58357 51357 58391 51391
rect 58391 51357 58400 51391
rect 58348 51348 58400 51357
rect 20444 51212 20496 51264
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 4620 51008 4672 51060
rect 3976 50983 4028 50992
rect 3976 50949 3985 50983
rect 3985 50949 4019 50983
rect 4019 50949 4028 50983
rect 3976 50940 4028 50949
rect 2596 50804 2648 50856
rect 4068 50915 4120 50924
rect 4068 50881 4082 50915
rect 4082 50881 4116 50915
rect 4116 50881 4120 50915
rect 4068 50872 4120 50881
rect 6276 50668 6328 50720
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 29920 50396 29972 50448
rect 41788 50396 41840 50448
rect 10140 50328 10192 50380
rect 29828 50328 29880 50380
rect 39488 50328 39540 50380
rect 55772 50328 55824 50380
rect 57428 50260 57480 50312
rect 1676 50235 1728 50244
rect 1676 50201 1685 50235
rect 1685 50201 1719 50235
rect 1719 50201 1728 50235
rect 1676 50192 1728 50201
rect 2044 50192 2096 50244
rect 57888 50124 57940 50176
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 1584 49827 1636 49836
rect 1584 49793 1593 49827
rect 1593 49793 1627 49827
rect 1627 49793 1636 49827
rect 1584 49784 1636 49793
rect 13084 49716 13136 49768
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 1584 49215 1636 49224
rect 1584 49181 1593 49215
rect 1593 49181 1627 49215
rect 1627 49181 1636 49215
rect 1584 49172 1636 49181
rect 57980 49147 58032 49156
rect 57980 49113 57989 49147
rect 57989 49113 58023 49147
rect 58023 49113 58032 49147
rect 57980 49104 58032 49113
rect 59084 49104 59136 49156
rect 18604 49036 18656 49088
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 1676 48739 1728 48748
rect 1676 48705 1685 48739
rect 1685 48705 1719 48739
rect 1719 48705 1728 48739
rect 1676 48696 1728 48705
rect 1952 48560 2004 48612
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 17868 48220 17920 48272
rect 2044 48127 2096 48136
rect 2044 48093 2053 48127
rect 2053 48093 2087 48127
rect 2087 48093 2096 48127
rect 2044 48084 2096 48093
rect 2872 48152 2924 48204
rect 4068 48152 4120 48204
rect 2412 48127 2464 48136
rect 2412 48093 2426 48127
rect 2426 48093 2460 48127
rect 2460 48093 2464 48127
rect 2412 48084 2464 48093
rect 57796 48084 57848 48136
rect 58164 48059 58216 48068
rect 1860 47948 1912 48000
rect 58164 48025 58173 48059
rect 58173 48025 58207 48059
rect 58207 48025 58216 48059
rect 58164 48016 58216 48025
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 53380 47744 53432 47796
rect 58072 47744 58124 47796
rect 1676 47651 1728 47660
rect 1676 47617 1685 47651
rect 1685 47617 1719 47651
rect 1719 47617 1728 47651
rect 1676 47608 1728 47617
rect 25412 47608 25464 47660
rect 40132 47608 40184 47660
rect 58072 47651 58124 47660
rect 58072 47617 58081 47651
rect 58081 47617 58115 47651
rect 58115 47617 58124 47651
rect 58072 47608 58124 47617
rect 10784 47540 10836 47592
rect 26240 47540 26292 47592
rect 35808 47540 35860 47592
rect 53196 47540 53248 47592
rect 6184 47472 6236 47524
rect 58808 47404 58860 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 1584 47039 1636 47048
rect 1584 47005 1593 47039
rect 1593 47005 1627 47039
rect 1627 47005 1636 47039
rect 1584 46996 1636 47005
rect 10324 46928 10376 46980
rect 32588 46928 32640 46980
rect 37924 46928 37976 46980
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 1584 46563 1636 46572
rect 1584 46529 1593 46563
rect 1593 46529 1627 46563
rect 1627 46529 1636 46563
rect 1584 46520 1636 46529
rect 36360 46316 36412 46368
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 58164 46019 58216 46028
rect 58164 45985 58173 46019
rect 58173 45985 58207 46019
rect 58207 45985 58216 46019
rect 58164 45976 58216 45985
rect 57704 45908 57756 45960
rect 1676 45883 1728 45892
rect 1676 45849 1685 45883
rect 1685 45849 1719 45883
rect 1719 45849 1728 45883
rect 1676 45840 1728 45849
rect 15200 45772 15252 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 15200 45500 15252 45552
rect 20720 45500 20772 45552
rect 35348 45500 35400 45552
rect 17408 45475 17460 45484
rect 17408 45441 17414 45475
rect 17414 45441 17448 45475
rect 17448 45441 17460 45475
rect 17408 45432 17460 45441
rect 23480 45432 23532 45484
rect 24216 45432 24268 45484
rect 36360 45475 36412 45484
rect 36360 45441 36369 45475
rect 36369 45441 36403 45475
rect 36403 45441 36412 45475
rect 36360 45432 36412 45441
rect 36636 45475 36688 45484
rect 36636 45441 36645 45475
rect 36645 45441 36679 45475
rect 36679 45441 36688 45475
rect 36636 45432 36688 45441
rect 37464 45432 37516 45484
rect 38016 45475 38068 45484
rect 38016 45441 38025 45475
rect 38025 45441 38059 45475
rect 38059 45441 38068 45475
rect 38016 45432 38068 45441
rect 35992 45364 36044 45416
rect 37188 45364 37240 45416
rect 57060 45432 57112 45484
rect 58072 45475 58124 45484
rect 58072 45441 58081 45475
rect 58081 45441 58115 45475
rect 58115 45441 58124 45475
rect 58072 45432 58124 45441
rect 36912 45339 36964 45348
rect 17684 45271 17736 45280
rect 17684 45237 17693 45271
rect 17693 45237 17727 45271
rect 17727 45237 17736 45271
rect 17684 45228 17736 45237
rect 36912 45305 36921 45339
rect 36921 45305 36955 45339
rect 36955 45305 36964 45339
rect 36912 45296 36964 45305
rect 58624 45228 58676 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 1584 44863 1636 44872
rect 1584 44829 1593 44863
rect 1593 44829 1627 44863
rect 1627 44829 1636 44863
rect 1584 44820 1636 44829
rect 56784 44820 56836 44872
rect 36820 44752 36872 44804
rect 57244 44795 57296 44804
rect 57244 44761 57253 44795
rect 57253 44761 57287 44795
rect 57287 44761 57296 44795
rect 57244 44752 57296 44761
rect 57888 44752 57940 44804
rect 58716 44752 58768 44804
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 34060 44480 34112 44532
rect 9220 44412 9272 44464
rect 1676 44387 1728 44396
rect 1676 44353 1685 44387
rect 1685 44353 1719 44387
rect 1719 44353 1728 44387
rect 1676 44344 1728 44353
rect 34060 44387 34112 44396
rect 34060 44353 34069 44387
rect 34069 44353 34103 44387
rect 34103 44353 34112 44387
rect 34060 44344 34112 44353
rect 34152 44344 34204 44396
rect 21456 44276 21508 44328
rect 45744 44344 45796 44396
rect 9588 44208 9640 44260
rect 34612 44251 34664 44260
rect 34612 44217 34621 44251
rect 34621 44217 34655 44251
rect 34655 44217 34664 44251
rect 34612 44208 34664 44217
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 34244 43911 34296 43920
rect 34244 43877 34253 43911
rect 34253 43877 34287 43911
rect 34287 43877 34296 43911
rect 34244 43868 34296 43877
rect 9588 43800 9640 43852
rect 1676 43707 1728 43716
rect 1676 43673 1685 43707
rect 1685 43673 1719 43707
rect 1719 43673 1728 43707
rect 1676 43664 1728 43673
rect 33048 43664 33100 43716
rect 57612 43732 57664 43784
rect 32312 43596 32364 43648
rect 33692 43596 33744 43648
rect 35900 43664 35952 43716
rect 58164 43707 58216 43716
rect 58164 43673 58173 43707
rect 58173 43673 58207 43707
rect 58207 43673 58216 43707
rect 58164 43664 58216 43673
rect 35348 43596 35400 43648
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 33232 43392 33284 43444
rect 33692 43392 33744 43444
rect 54852 43324 54904 43376
rect 1584 43299 1636 43308
rect 1584 43265 1593 43299
rect 1593 43265 1627 43299
rect 1627 43265 1636 43299
rect 1584 43256 1636 43265
rect 32312 43299 32364 43308
rect 32312 43265 32321 43299
rect 32321 43265 32355 43299
rect 32355 43265 32364 43299
rect 32312 43256 32364 43265
rect 32772 43299 32824 43308
rect 32772 43265 32775 43299
rect 32775 43265 32824 43299
rect 32772 43256 32824 43265
rect 1768 43095 1820 43104
rect 1768 43061 1777 43095
rect 1777 43061 1811 43095
rect 1811 43061 1820 43095
rect 1768 43052 1820 43061
rect 32956 43052 33008 43104
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 32772 42712 32824 42764
rect 33048 42687 33100 42696
rect 33048 42653 33057 42687
rect 33057 42653 33091 42687
rect 33091 42653 33100 42687
rect 33048 42644 33100 42653
rect 33140 42687 33192 42696
rect 33140 42653 33149 42687
rect 33149 42653 33183 42687
rect 33183 42653 33192 42687
rect 33140 42644 33192 42653
rect 33692 42687 33744 42696
rect 32772 42508 32824 42560
rect 33692 42653 33701 42687
rect 33701 42653 33735 42687
rect 33735 42653 33744 42687
rect 33692 42644 33744 42653
rect 33876 42687 33928 42696
rect 33876 42653 33885 42687
rect 33885 42653 33919 42687
rect 33919 42653 33928 42687
rect 33876 42644 33928 42653
rect 34244 42644 34296 42696
rect 34796 42644 34848 42696
rect 37280 42687 37332 42696
rect 37280 42653 37289 42687
rect 37289 42653 37323 42687
rect 37323 42653 37332 42687
rect 37280 42644 37332 42653
rect 37464 42619 37516 42628
rect 37464 42585 37473 42619
rect 37473 42585 37507 42619
rect 37507 42585 37516 42619
rect 37464 42576 37516 42585
rect 54300 42576 54352 42628
rect 57060 42619 57112 42628
rect 57060 42585 57069 42619
rect 57069 42585 57103 42619
rect 57103 42585 57112 42619
rect 57060 42576 57112 42585
rect 57980 42619 58032 42628
rect 57980 42585 57989 42619
rect 57989 42585 58023 42619
rect 58023 42585 58032 42619
rect 57980 42576 58032 42585
rect 58348 42619 58400 42628
rect 58348 42585 58357 42619
rect 58357 42585 58391 42619
rect 58391 42585 58400 42619
rect 58348 42576 58400 42585
rect 57336 42551 57388 42560
rect 57336 42517 57345 42551
rect 57345 42517 57379 42551
rect 57379 42517 57388 42551
rect 57336 42508 57388 42517
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 1768 42304 1820 42356
rect 33876 42304 33928 42356
rect 1584 42211 1636 42220
rect 1584 42177 1593 42211
rect 1593 42177 1627 42211
rect 1627 42177 1636 42211
rect 1584 42168 1636 42177
rect 2136 41964 2188 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 54668 41556 54720 41608
rect 1676 41531 1728 41540
rect 1676 41497 1685 41531
rect 1685 41497 1719 41531
rect 1719 41497 1728 41531
rect 1676 41488 1728 41497
rect 57244 41531 57296 41540
rect 57244 41497 57253 41531
rect 57253 41497 57287 41531
rect 57287 41497 57296 41531
rect 57244 41488 57296 41497
rect 57888 41488 57940 41540
rect 58440 41488 58492 41540
rect 26884 41420 26936 41472
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 1676 41123 1728 41132
rect 1676 41089 1685 41123
rect 1685 41089 1719 41123
rect 1719 41089 1728 41123
rect 1676 41080 1728 41089
rect 21180 40876 21232 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 57520 40468 57572 40520
rect 1676 40443 1728 40452
rect 1676 40409 1685 40443
rect 1685 40409 1719 40443
rect 1719 40409 1728 40443
rect 1676 40400 1728 40409
rect 18604 40400 18656 40452
rect 22468 40400 22520 40452
rect 36636 40400 36688 40452
rect 45100 40400 45152 40452
rect 57060 40443 57112 40452
rect 57060 40409 57069 40443
rect 57069 40409 57103 40443
rect 57103 40409 57112 40443
rect 57060 40400 57112 40409
rect 23296 40332 23348 40384
rect 47584 40332 47636 40384
rect 57888 40332 57940 40384
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 20904 40128 20956 40180
rect 23480 40128 23532 40180
rect 25320 40128 25372 40180
rect 21180 40103 21232 40112
rect 21180 40069 21189 40103
rect 21189 40069 21223 40103
rect 21223 40069 21232 40103
rect 21180 40060 21232 40069
rect 20996 39992 21048 40044
rect 2780 39924 2832 39976
rect 23756 39992 23808 40044
rect 21732 39788 21784 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 2228 39516 2280 39568
rect 2412 39516 2464 39568
rect 22284 39516 22336 39568
rect 2320 39423 2372 39432
rect 2320 39389 2329 39423
rect 2329 39389 2363 39423
rect 2363 39389 2372 39423
rect 2320 39380 2372 39389
rect 2780 39423 2832 39432
rect 2780 39389 2783 39423
rect 2783 39389 2832 39423
rect 2780 39380 2832 39389
rect 1676 39355 1728 39364
rect 1676 39321 1685 39355
rect 1685 39321 1719 39355
rect 1719 39321 1728 39355
rect 1676 39312 1728 39321
rect 2412 39244 2464 39296
rect 13084 39312 13136 39364
rect 23572 39312 23624 39364
rect 57060 39355 57112 39364
rect 57060 39321 57069 39355
rect 57069 39321 57103 39355
rect 57103 39321 57112 39355
rect 57060 39312 57112 39321
rect 57980 39355 58032 39364
rect 57980 39321 57989 39355
rect 57989 39321 58023 39355
rect 58023 39321 58032 39355
rect 57980 39312 58032 39321
rect 2596 39244 2648 39296
rect 33784 39244 33836 39296
rect 58072 39287 58124 39296
rect 58072 39253 58081 39287
rect 58081 39253 58115 39287
rect 58115 39253 58124 39287
rect 58072 39244 58124 39253
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 1676 38947 1728 38956
rect 1676 38913 1685 38947
rect 1685 38913 1719 38947
rect 1719 38913 1728 38947
rect 1676 38904 1728 38913
rect 22928 38947 22980 38956
rect 22928 38913 22937 38947
rect 22937 38913 22971 38947
rect 22971 38913 22980 38947
rect 22928 38904 22980 38913
rect 23296 39015 23348 39024
rect 23296 38981 23302 39015
rect 23302 38981 23336 39015
rect 23336 38981 23348 39015
rect 23296 38972 23348 38981
rect 23204 38947 23256 38956
rect 23204 38913 23213 38947
rect 23213 38913 23247 38947
rect 23247 38913 23256 38947
rect 23204 38904 23256 38913
rect 50712 39040 50764 39092
rect 58072 39040 58124 39092
rect 37004 38836 37056 38888
rect 1860 38811 1912 38820
rect 1860 38777 1869 38811
rect 1869 38777 1903 38811
rect 1903 38777 1912 38811
rect 1860 38768 1912 38777
rect 23112 38768 23164 38820
rect 24768 38700 24820 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 1860 38360 1912 38412
rect 16304 38496 16356 38548
rect 19156 38428 19208 38480
rect 23020 38496 23072 38548
rect 19432 38360 19484 38412
rect 19984 38360 20036 38412
rect 20628 38360 20680 38412
rect 39580 38360 39632 38412
rect 2780 38335 2832 38344
rect 2780 38301 2789 38335
rect 2789 38301 2823 38335
rect 2823 38301 2832 38335
rect 20168 38335 20220 38344
rect 2780 38292 2832 38301
rect 20168 38301 20177 38335
rect 20177 38301 20211 38335
rect 20211 38301 20220 38335
rect 20168 38292 20220 38301
rect 1676 38267 1728 38276
rect 1676 38233 1685 38267
rect 1685 38233 1719 38267
rect 1719 38233 1728 38267
rect 1676 38224 1728 38233
rect 20168 38156 20220 38208
rect 20536 38292 20588 38344
rect 21732 38335 21784 38344
rect 21732 38301 21741 38335
rect 21741 38301 21775 38335
rect 21775 38301 21784 38335
rect 21732 38292 21784 38301
rect 22928 38292 22980 38344
rect 46848 38292 46900 38344
rect 21088 38224 21140 38276
rect 58164 38267 58216 38276
rect 58164 38233 58173 38267
rect 58173 38233 58207 38267
rect 58207 38233 58216 38267
rect 58164 38224 58216 38233
rect 21824 38156 21876 38208
rect 22008 38156 22060 38208
rect 23020 38156 23072 38208
rect 26148 38156 26200 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 5908 37952 5960 38004
rect 2872 37884 2924 37936
rect 6184 37884 6236 37936
rect 1952 37816 2004 37868
rect 2228 37748 2280 37800
rect 3056 37816 3108 37868
rect 19340 37859 19392 37868
rect 19340 37825 19349 37859
rect 19349 37825 19383 37859
rect 19383 37825 19392 37859
rect 19340 37816 19392 37825
rect 2320 37680 2372 37732
rect 2596 37655 2648 37664
rect 2596 37621 2605 37655
rect 2605 37621 2639 37655
rect 2639 37621 2648 37655
rect 2596 37612 2648 37621
rect 19708 37859 19760 37868
rect 19708 37825 19717 37859
rect 19717 37825 19751 37859
rect 19751 37825 19760 37859
rect 19708 37816 19760 37825
rect 20260 37816 20312 37868
rect 20812 37859 20864 37868
rect 20812 37825 20821 37859
rect 20821 37825 20855 37859
rect 20855 37825 20864 37859
rect 20812 37816 20864 37825
rect 20904 37816 20956 37868
rect 21088 37859 21140 37868
rect 21088 37825 21097 37859
rect 21097 37825 21131 37859
rect 21131 37825 21140 37859
rect 21088 37816 21140 37825
rect 23020 37952 23072 38004
rect 22928 37927 22980 37936
rect 22928 37893 22937 37927
rect 22937 37893 22971 37927
rect 22971 37893 22980 37927
rect 22928 37884 22980 37893
rect 23020 37859 23072 37868
rect 23020 37825 23029 37859
rect 23029 37825 23063 37859
rect 23063 37825 23072 37859
rect 23020 37816 23072 37825
rect 25228 37927 25280 37936
rect 22560 37748 22612 37800
rect 20444 37680 20496 37732
rect 21272 37680 21324 37732
rect 25228 37893 25237 37927
rect 25237 37893 25271 37927
rect 25271 37893 25280 37927
rect 25228 37884 25280 37893
rect 25320 37859 25372 37868
rect 23940 37748 23992 37800
rect 24124 37791 24176 37800
rect 24124 37757 24133 37791
rect 24133 37757 24167 37791
rect 24167 37757 24176 37791
rect 24124 37748 24176 37757
rect 25320 37825 25329 37859
rect 25329 37825 25363 37859
rect 25363 37825 25372 37859
rect 25320 37816 25372 37825
rect 26148 37952 26200 38004
rect 37464 37884 37516 37936
rect 29736 37816 29788 37868
rect 58072 37859 58124 37868
rect 58072 37825 58081 37859
rect 58081 37825 58115 37859
rect 58115 37825 58124 37859
rect 58072 37816 58124 37825
rect 44180 37748 44232 37800
rect 20352 37612 20404 37664
rect 20628 37655 20680 37664
rect 20628 37621 20637 37655
rect 20637 37621 20671 37655
rect 20671 37621 20680 37655
rect 20628 37612 20680 37621
rect 24400 37655 24452 37664
rect 24400 37621 24409 37655
rect 24409 37621 24443 37655
rect 24443 37621 24452 37655
rect 24400 37612 24452 37621
rect 58532 37612 58584 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 2596 37408 2648 37460
rect 16304 37408 16356 37460
rect 16488 37408 16540 37460
rect 20720 37408 20772 37460
rect 20812 37408 20864 37460
rect 54208 37408 54260 37460
rect 20260 37340 20312 37392
rect 23112 37340 23164 37392
rect 2688 37272 2740 37324
rect 3056 37272 3108 37324
rect 1676 37247 1728 37256
rect 1676 37213 1685 37247
rect 1685 37213 1719 37247
rect 1719 37213 1728 37247
rect 1676 37204 1728 37213
rect 5540 37111 5592 37120
rect 5540 37077 5549 37111
rect 5549 37077 5583 37111
rect 5583 37077 5592 37111
rect 5540 37068 5592 37077
rect 6000 37247 6052 37256
rect 6000 37213 6009 37247
rect 6009 37213 6043 37247
rect 6043 37213 6052 37247
rect 6276 37247 6328 37256
rect 6000 37204 6052 37213
rect 6276 37213 6285 37247
rect 6285 37213 6319 37247
rect 6319 37213 6328 37247
rect 6276 37204 6328 37213
rect 9036 37272 9088 37324
rect 21088 37315 21140 37324
rect 21088 37281 21097 37315
rect 21097 37281 21131 37315
rect 21131 37281 21140 37315
rect 21088 37272 21140 37281
rect 6736 37247 6788 37256
rect 6736 37213 6745 37247
rect 6745 37213 6779 37247
rect 6779 37213 6788 37247
rect 6736 37204 6788 37213
rect 19340 37204 19392 37256
rect 20536 37204 20588 37256
rect 21916 37204 21968 37256
rect 53840 37247 53892 37256
rect 53840 37213 53849 37247
rect 53849 37213 53883 37247
rect 53883 37213 53892 37247
rect 53840 37204 53892 37213
rect 54116 37247 54168 37256
rect 54116 37213 54125 37247
rect 54125 37213 54159 37247
rect 54159 37213 54168 37247
rect 54116 37204 54168 37213
rect 54300 37247 54352 37256
rect 54300 37213 54303 37247
rect 54303 37213 54352 37247
rect 54300 37204 54352 37213
rect 54484 37204 54536 37256
rect 18788 37136 18840 37188
rect 20996 37136 21048 37188
rect 54024 37179 54076 37188
rect 54024 37145 54033 37179
rect 54033 37145 54067 37179
rect 54067 37145 54076 37179
rect 54024 37136 54076 37145
rect 58164 37179 58216 37188
rect 58164 37145 58173 37179
rect 58173 37145 58207 37179
rect 58207 37145 58216 37179
rect 58164 37136 58216 37145
rect 9036 37068 9088 37120
rect 19248 37068 19300 37120
rect 49976 37068 50028 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 6000 36864 6052 36916
rect 42892 36864 42944 36916
rect 18880 36796 18932 36848
rect 20076 36796 20128 36848
rect 20260 36796 20312 36848
rect 20536 36796 20588 36848
rect 28448 36796 28500 36848
rect 36268 36796 36320 36848
rect 53932 36839 53984 36848
rect 53932 36805 53941 36839
rect 53941 36805 53975 36839
rect 53975 36805 53984 36839
rect 53932 36796 53984 36805
rect 1584 36771 1636 36780
rect 1584 36737 1593 36771
rect 1593 36737 1627 36771
rect 1627 36737 1636 36771
rect 1584 36728 1636 36737
rect 18420 36771 18472 36780
rect 18420 36737 18429 36771
rect 18429 36737 18463 36771
rect 18463 36737 18472 36771
rect 18420 36728 18472 36737
rect 18788 36771 18840 36780
rect 18788 36737 18797 36771
rect 18797 36737 18831 36771
rect 18831 36737 18840 36771
rect 18788 36728 18840 36737
rect 19432 36771 19484 36780
rect 19432 36737 19441 36771
rect 19441 36737 19475 36771
rect 19475 36737 19484 36771
rect 19432 36728 19484 36737
rect 20996 36728 21048 36780
rect 20168 36660 20220 36712
rect 23848 36703 23900 36712
rect 19340 36592 19392 36644
rect 23848 36669 23857 36703
rect 23857 36669 23891 36703
rect 23891 36669 23900 36703
rect 23848 36660 23900 36669
rect 24032 36771 24084 36780
rect 24032 36737 24041 36771
rect 24041 36737 24075 36771
rect 24075 36737 24084 36771
rect 24032 36728 24084 36737
rect 25504 36728 25556 36780
rect 53656 36771 53708 36780
rect 53656 36737 53665 36771
rect 53665 36737 53699 36771
rect 53699 36737 53708 36771
rect 53656 36728 53708 36737
rect 37280 36660 37332 36712
rect 49976 36592 50028 36644
rect 54024 36592 54076 36644
rect 54208 36635 54260 36644
rect 54208 36601 54217 36635
rect 54217 36601 54251 36635
rect 54251 36601 54260 36635
rect 54208 36592 54260 36601
rect 2596 36524 2648 36576
rect 20076 36524 20128 36576
rect 23480 36524 23532 36576
rect 24584 36524 24636 36576
rect 53840 36524 53892 36576
rect 55036 36524 55088 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 23480 36320 23532 36372
rect 23848 36363 23900 36372
rect 23848 36329 23857 36363
rect 23857 36329 23891 36363
rect 23891 36329 23900 36363
rect 23848 36320 23900 36329
rect 6736 36252 6788 36304
rect 20628 36252 20680 36304
rect 20996 36252 21048 36304
rect 23204 36252 23256 36304
rect 20720 36227 20772 36236
rect 20720 36193 20729 36227
rect 20729 36193 20763 36227
rect 20763 36193 20772 36227
rect 20720 36184 20772 36193
rect 2504 36159 2556 36168
rect 2504 36125 2513 36159
rect 2513 36125 2547 36159
rect 2547 36125 2556 36159
rect 2504 36116 2556 36125
rect 2872 36159 2924 36168
rect 2872 36125 2886 36159
rect 2886 36125 2920 36159
rect 2920 36125 2924 36159
rect 2872 36116 2924 36125
rect 3056 36116 3108 36168
rect 20168 36159 20220 36168
rect 20168 36125 20177 36159
rect 20177 36125 20211 36159
rect 20211 36125 20220 36159
rect 20168 36116 20220 36125
rect 20444 36159 20496 36168
rect 20444 36125 20453 36159
rect 20453 36125 20487 36159
rect 20487 36125 20496 36159
rect 20444 36116 20496 36125
rect 22192 36159 22244 36168
rect 22192 36125 22201 36159
rect 22201 36125 22235 36159
rect 22235 36125 22244 36159
rect 22192 36116 22244 36125
rect 22468 36159 22520 36168
rect 22468 36125 22477 36159
rect 22477 36125 22511 36159
rect 22511 36125 22520 36159
rect 22468 36116 22520 36125
rect 23296 36159 23348 36168
rect 23296 36125 23305 36159
rect 23305 36125 23339 36159
rect 23339 36125 23348 36159
rect 23296 36116 23348 36125
rect 23388 36116 23440 36168
rect 33232 36184 33284 36236
rect 24584 36159 24636 36168
rect 24584 36125 24593 36159
rect 24593 36125 24627 36159
rect 24627 36125 24636 36159
rect 24584 36116 24636 36125
rect 24768 36159 24820 36168
rect 24768 36125 24777 36159
rect 24777 36125 24811 36159
rect 24811 36125 24820 36159
rect 24768 36116 24820 36125
rect 1676 36091 1728 36100
rect 1676 36057 1685 36091
rect 1685 36057 1719 36091
rect 1719 36057 1728 36091
rect 1676 36048 1728 36057
rect 2412 36048 2464 36100
rect 2780 36091 2832 36100
rect 2780 36057 2789 36091
rect 2789 36057 2823 36091
rect 2823 36057 2832 36091
rect 2780 36048 2832 36057
rect 15752 35980 15804 36032
rect 16488 35980 16540 36032
rect 22744 36023 22796 36032
rect 22744 35989 22753 36023
rect 22753 35989 22787 36023
rect 22787 35989 22796 36023
rect 22744 35980 22796 35989
rect 23572 36091 23624 36100
rect 23572 36057 23581 36091
rect 23581 36057 23615 36091
rect 23615 36057 23624 36091
rect 23572 36048 23624 36057
rect 25412 36048 25464 36100
rect 57980 36091 58032 36100
rect 57980 36057 57989 36091
rect 57989 36057 58023 36091
rect 58023 36057 58032 36091
rect 57980 36048 58032 36057
rect 58900 36048 58952 36100
rect 24952 35980 25004 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 1768 35819 1820 35828
rect 1768 35785 1777 35819
rect 1777 35785 1811 35819
rect 1811 35785 1820 35819
rect 1768 35776 1820 35785
rect 19340 35776 19392 35828
rect 19248 35751 19300 35760
rect 19248 35717 19257 35751
rect 19257 35717 19291 35751
rect 19291 35717 19300 35751
rect 19248 35708 19300 35717
rect 20168 35776 20220 35828
rect 33048 35776 33100 35828
rect 37280 35776 37332 35828
rect 1676 35683 1728 35692
rect 1676 35649 1685 35683
rect 1685 35649 1719 35683
rect 1719 35649 1728 35683
rect 1676 35640 1728 35649
rect 16580 35640 16632 35692
rect 24676 35708 24728 35760
rect 29736 35708 29788 35760
rect 19340 35504 19392 35556
rect 21088 35640 21140 35692
rect 24124 35640 24176 35692
rect 40592 35683 40644 35692
rect 40592 35649 40601 35683
rect 40601 35649 40635 35683
rect 40635 35649 40644 35683
rect 40592 35640 40644 35649
rect 23388 35615 23440 35624
rect 23388 35581 23397 35615
rect 23397 35581 23431 35615
rect 23431 35581 23440 35615
rect 23388 35572 23440 35581
rect 40408 35572 40460 35624
rect 22192 35504 22244 35556
rect 40592 35504 40644 35556
rect 41696 35572 41748 35624
rect 48964 35504 49016 35556
rect 20076 35479 20128 35488
rect 20076 35445 20085 35479
rect 20085 35445 20119 35479
rect 20119 35445 20128 35479
rect 20076 35436 20128 35445
rect 33048 35436 33100 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 2688 35232 2740 35284
rect 13820 35232 13872 35284
rect 22744 35275 22796 35284
rect 22744 35241 22753 35275
rect 22753 35241 22787 35275
rect 22787 35241 22796 35275
rect 22744 35232 22796 35241
rect 2780 35164 2832 35216
rect 23296 35164 23348 35216
rect 31760 35164 31812 35216
rect 40684 35232 40736 35284
rect 47676 35232 47728 35284
rect 22284 35028 22336 35080
rect 24860 35028 24912 35080
rect 31760 35028 31812 35080
rect 53196 35164 53248 35216
rect 40500 35096 40552 35148
rect 40316 35071 40368 35080
rect 40316 35037 40325 35071
rect 40325 35037 40359 35071
rect 40359 35037 40368 35071
rect 40316 35028 40368 35037
rect 40408 35071 40460 35080
rect 40408 35037 40417 35071
rect 40417 35037 40451 35071
rect 40451 35037 40460 35071
rect 40408 35028 40460 35037
rect 51632 35028 51684 35080
rect 1676 35003 1728 35012
rect 1676 34969 1685 35003
rect 1685 34969 1719 35003
rect 1719 34969 1728 35003
rect 1676 34960 1728 34969
rect 23204 34960 23256 35012
rect 58164 35003 58216 35012
rect 58164 34969 58173 35003
rect 58173 34969 58207 35003
rect 58207 34969 58216 35003
rect 58164 34960 58216 34969
rect 23020 34935 23072 34944
rect 23020 34901 23029 34935
rect 23029 34901 23063 34935
rect 23063 34901 23072 34935
rect 23020 34892 23072 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 19340 34688 19392 34740
rect 39120 34688 39172 34740
rect 58992 34688 59044 34740
rect 19984 34620 20036 34672
rect 22376 34620 22428 34672
rect 19432 34552 19484 34604
rect 22836 34552 22888 34604
rect 57888 34552 57940 34604
rect 20996 34416 21048 34468
rect 23204 34416 23256 34468
rect 23572 34416 23624 34468
rect 40408 34416 40460 34468
rect 43260 34416 43312 34468
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 21732 34144 21784 34196
rect 17316 34076 17368 34128
rect 21548 34076 21600 34128
rect 21364 33983 21416 33992
rect 21364 33949 21373 33983
rect 21373 33949 21407 33983
rect 21407 33949 21416 33983
rect 21364 33940 21416 33949
rect 21548 33983 21600 33992
rect 21548 33949 21555 33983
rect 21555 33949 21600 33983
rect 21548 33940 21600 33949
rect 22192 34076 22244 34128
rect 23020 33983 23072 33992
rect 1676 33915 1728 33924
rect 1676 33881 1685 33915
rect 1685 33881 1719 33915
rect 1719 33881 1728 33915
rect 1676 33872 1728 33881
rect 21272 33872 21324 33924
rect 1768 33847 1820 33856
rect 1768 33813 1777 33847
rect 1777 33813 1811 33847
rect 1811 33813 1820 33847
rect 1768 33804 1820 33813
rect 17132 33804 17184 33856
rect 23020 33949 23029 33983
rect 23029 33949 23063 33983
rect 23063 33949 23072 33983
rect 23020 33940 23072 33949
rect 24492 33940 24544 33992
rect 25320 33940 25372 33992
rect 24032 33872 24084 33924
rect 24860 33915 24912 33924
rect 24860 33881 24869 33915
rect 24869 33881 24903 33915
rect 24903 33881 24912 33915
rect 24860 33872 24912 33881
rect 46296 34008 46348 34060
rect 22744 33804 22796 33856
rect 26976 33872 27028 33924
rect 25228 33847 25280 33856
rect 25228 33813 25237 33847
rect 25237 33813 25271 33847
rect 25271 33813 25280 33847
rect 25228 33804 25280 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 1768 33600 1820 33652
rect 17132 33600 17184 33652
rect 22284 33600 22336 33652
rect 34152 33600 34204 33652
rect 2320 33532 2372 33584
rect 12164 33532 12216 33584
rect 1676 33507 1728 33516
rect 1676 33473 1685 33507
rect 1685 33473 1719 33507
rect 1719 33473 1728 33507
rect 1676 33464 1728 33473
rect 16948 33260 17000 33312
rect 20904 33260 20956 33312
rect 21088 33507 21140 33516
rect 21088 33473 21097 33507
rect 21097 33473 21131 33507
rect 21131 33473 21140 33507
rect 21456 33532 21508 33584
rect 21088 33464 21140 33473
rect 22192 33507 22244 33516
rect 22192 33473 22199 33507
rect 22199 33473 22244 33507
rect 22192 33464 22244 33473
rect 36084 33575 36136 33584
rect 22376 33507 22428 33516
rect 22376 33473 22385 33507
rect 22385 33473 22419 33507
rect 22419 33473 22428 33507
rect 22376 33464 22428 33473
rect 22560 33464 22612 33516
rect 22836 33464 22888 33516
rect 36084 33541 36093 33575
rect 36093 33541 36127 33575
rect 36127 33541 36136 33575
rect 36084 33532 36136 33541
rect 32220 33464 32272 33516
rect 35808 33507 35860 33516
rect 35808 33473 35818 33507
rect 35818 33473 35852 33507
rect 35852 33473 35860 33507
rect 35808 33464 35860 33473
rect 35992 33507 36044 33516
rect 35992 33473 36001 33507
rect 36001 33473 36035 33507
rect 36035 33473 36044 33507
rect 40408 33600 40460 33652
rect 35992 33464 36044 33473
rect 40408 33396 40460 33448
rect 23296 33328 23348 33380
rect 35992 33328 36044 33380
rect 22652 33303 22704 33312
rect 22652 33269 22661 33303
rect 22661 33269 22695 33303
rect 22695 33269 22704 33303
rect 22652 33260 22704 33269
rect 37648 33260 37700 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 20904 33056 20956 33108
rect 21732 33056 21784 33108
rect 22652 32988 22704 33040
rect 25228 32988 25280 33040
rect 58164 32963 58216 32972
rect 58164 32929 58173 32963
rect 58173 32929 58207 32963
rect 58207 32929 58216 32963
rect 58164 32920 58216 32929
rect 21824 32895 21876 32904
rect 21824 32861 21833 32895
rect 21833 32861 21867 32895
rect 21867 32861 21876 32895
rect 21824 32852 21876 32861
rect 23204 32852 23256 32904
rect 24768 32895 24820 32904
rect 24768 32861 24777 32895
rect 24777 32861 24811 32895
rect 24811 32861 24820 32895
rect 24768 32852 24820 32861
rect 37556 32852 37608 32904
rect 56140 32852 56192 32904
rect 1676 32827 1728 32836
rect 1676 32793 1685 32827
rect 1685 32793 1719 32827
rect 1719 32793 1728 32827
rect 1676 32784 1728 32793
rect 22192 32784 22244 32836
rect 57060 32827 57112 32836
rect 16580 32716 16632 32768
rect 22100 32716 22152 32768
rect 57060 32793 57069 32827
rect 57069 32793 57103 32827
rect 57103 32793 57112 32827
rect 57060 32784 57112 32793
rect 55864 32716 55916 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 16488 32444 16540 32496
rect 22284 32444 22336 32496
rect 1676 32419 1728 32428
rect 1676 32385 1685 32419
rect 1685 32385 1719 32419
rect 1719 32385 1728 32419
rect 1676 32376 1728 32385
rect 22008 32376 22060 32428
rect 29184 32376 29236 32428
rect 22744 32172 22796 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 20260 31900 20312 31952
rect 22928 31900 22980 31952
rect 22744 31807 22796 31816
rect 22744 31773 22753 31807
rect 22753 31773 22787 31807
rect 22787 31773 22796 31807
rect 22744 31764 22796 31773
rect 23296 31900 23348 31952
rect 58256 31900 58308 31952
rect 21732 31696 21784 31748
rect 49148 31764 49200 31816
rect 58164 31807 58216 31816
rect 58164 31773 58173 31807
rect 58173 31773 58207 31807
rect 58207 31773 58216 31807
rect 58164 31764 58216 31773
rect 23296 31671 23348 31680
rect 23296 31637 23305 31671
rect 23305 31637 23339 31671
rect 23339 31637 23348 31671
rect 23296 31628 23348 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 19248 31424 19300 31476
rect 24584 31424 24636 31476
rect 1676 31331 1728 31340
rect 1676 31297 1685 31331
rect 1685 31297 1719 31331
rect 1719 31297 1728 31331
rect 1676 31288 1728 31297
rect 24124 31331 24176 31340
rect 24124 31297 24133 31331
rect 24133 31297 24167 31331
rect 24167 31297 24176 31331
rect 24124 31288 24176 31297
rect 24216 31331 24268 31340
rect 24216 31297 24226 31331
rect 24226 31297 24260 31331
rect 24260 31297 24268 31331
rect 24216 31288 24268 31297
rect 21272 31220 21324 31272
rect 22744 31220 22796 31272
rect 10324 31152 10376 31204
rect 21824 31152 21876 31204
rect 24584 31331 24636 31340
rect 24584 31297 24617 31331
rect 24617 31297 24636 31331
rect 58072 31331 58124 31340
rect 24584 31288 24636 31297
rect 58072 31297 58081 31331
rect 58081 31297 58115 31331
rect 58115 31297 58124 31331
rect 58072 31288 58124 31297
rect 24768 31195 24820 31204
rect 24768 31161 24777 31195
rect 24777 31161 24811 31195
rect 24811 31161 24820 31195
rect 24768 31152 24820 31161
rect 44180 31084 44232 31136
rect 49792 31084 49844 31136
rect 59176 31084 59228 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 23296 30880 23348 30932
rect 24216 30880 24268 30932
rect 29092 30880 29144 30932
rect 19340 30744 19392 30796
rect 34704 30744 34756 30796
rect 23112 30719 23164 30728
rect 1676 30651 1728 30660
rect 1676 30617 1685 30651
rect 1685 30617 1719 30651
rect 1719 30617 1728 30651
rect 1676 30608 1728 30617
rect 17684 30608 17736 30660
rect 23112 30685 23121 30719
rect 23121 30685 23155 30719
rect 23155 30685 23164 30719
rect 23112 30676 23164 30685
rect 23204 30676 23256 30728
rect 23572 30719 23624 30728
rect 20352 30608 20404 30660
rect 22284 30608 22336 30660
rect 23572 30685 23581 30719
rect 23581 30685 23615 30719
rect 23615 30685 23624 30719
rect 23572 30676 23624 30685
rect 32220 30608 32272 30660
rect 17960 30540 18012 30592
rect 24860 30540 24912 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 17960 30336 18012 30388
rect 19340 30379 19392 30388
rect 15108 30268 15160 30320
rect 19340 30345 19349 30379
rect 19349 30345 19383 30379
rect 19383 30345 19392 30379
rect 19340 30336 19392 30345
rect 1584 30243 1636 30252
rect 1584 30209 1593 30243
rect 1593 30209 1627 30243
rect 1627 30209 1636 30243
rect 1584 30200 1636 30209
rect 18880 30243 18932 30252
rect 18880 30209 18887 30243
rect 18887 30209 18932 30243
rect 1768 30175 1820 30184
rect 1768 30141 1777 30175
rect 1777 30141 1811 30175
rect 1811 30141 1820 30175
rect 1768 30132 1820 30141
rect 18880 30200 18932 30209
rect 18972 30243 19024 30252
rect 18972 30209 18981 30243
rect 18981 30209 19015 30243
rect 19015 30209 19024 30243
rect 18972 30200 19024 30209
rect 19248 30200 19300 30252
rect 22284 30243 22336 30252
rect 22284 30209 22293 30243
rect 22293 30209 22327 30243
rect 22327 30209 22336 30243
rect 22284 30200 22336 30209
rect 22560 30243 22612 30252
rect 22560 30209 22569 30243
rect 22569 30209 22603 30243
rect 22603 30209 22612 30243
rect 22560 30200 22612 30209
rect 21640 30132 21692 30184
rect 22468 30132 22520 30184
rect 24124 30064 24176 30116
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 22560 29792 22612 29844
rect 23112 29835 23164 29844
rect 23112 29801 23121 29835
rect 23121 29801 23155 29835
rect 23155 29801 23164 29835
rect 23112 29792 23164 29801
rect 13820 29656 13872 29708
rect 1952 29588 2004 29640
rect 2596 29588 2648 29640
rect 9956 29588 10008 29640
rect 21548 29631 21600 29640
rect 21548 29597 21557 29631
rect 21557 29597 21591 29631
rect 21591 29597 21600 29631
rect 21548 29588 21600 29597
rect 21916 29631 21968 29640
rect 21916 29597 21925 29631
rect 21925 29597 21959 29631
rect 21959 29597 21968 29631
rect 21916 29588 21968 29597
rect 1860 29563 1912 29572
rect 1860 29529 1869 29563
rect 1869 29529 1903 29563
rect 1903 29529 1912 29563
rect 1860 29520 1912 29529
rect 18972 29520 19024 29572
rect 21824 29563 21876 29572
rect 21824 29529 21833 29563
rect 21833 29529 21867 29563
rect 21867 29529 21876 29563
rect 33140 29656 33192 29708
rect 35532 29656 35584 29708
rect 51724 29656 51776 29708
rect 58164 29699 58216 29708
rect 58164 29665 58173 29699
rect 58173 29665 58207 29699
rect 58207 29665 58216 29699
rect 58164 29656 58216 29665
rect 23020 29588 23072 29640
rect 57152 29588 57204 29640
rect 21824 29520 21876 29529
rect 22744 29563 22796 29572
rect 22744 29529 22753 29563
rect 22753 29529 22787 29563
rect 22787 29529 22796 29563
rect 22744 29520 22796 29529
rect 23388 29520 23440 29572
rect 57060 29563 57112 29572
rect 57060 29529 57069 29563
rect 57069 29529 57103 29563
rect 57103 29529 57112 29563
rect 57060 29520 57112 29529
rect 24952 29452 25004 29504
rect 44824 29452 44876 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 1584 29248 1636 29300
rect 21548 29248 21600 29300
rect 49056 29248 49108 29300
rect 15108 29112 15160 29164
rect 21732 29112 21784 29164
rect 23020 29112 23072 29164
rect 9680 29044 9732 29096
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 5540 28568 5592 28620
rect 29276 28568 29328 28620
rect 1860 28475 1912 28484
rect 1860 28441 1869 28475
rect 1869 28441 1903 28475
rect 1903 28441 1912 28475
rect 1860 28432 1912 28441
rect 2964 28500 3016 28552
rect 8944 28500 8996 28552
rect 9680 28432 9732 28484
rect 12808 28500 12860 28552
rect 22652 28500 22704 28552
rect 23296 28500 23348 28552
rect 29092 28500 29144 28552
rect 46480 28500 46532 28552
rect 55588 28500 55640 28552
rect 34060 28432 34112 28484
rect 58164 28475 58216 28484
rect 58164 28441 58173 28475
rect 58173 28441 58207 28475
rect 58207 28441 58216 28475
rect 58164 28432 58216 28441
rect 20444 28364 20496 28416
rect 47308 28364 47360 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 22836 28092 22888 28144
rect 2228 28024 2280 28076
rect 23112 28067 23164 28076
rect 23112 28033 23121 28067
rect 23121 28033 23155 28067
rect 23155 28033 23164 28067
rect 23112 28024 23164 28033
rect 23572 28092 23624 28144
rect 1768 27999 1820 28008
rect 1768 27965 1777 27999
rect 1777 27965 1811 27999
rect 1811 27965 1820 27999
rect 1768 27956 1820 27965
rect 23296 27956 23348 28008
rect 37280 28024 37332 28076
rect 23020 27820 23072 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 23664 27616 23716 27668
rect 2136 27480 2188 27532
rect 1584 27455 1636 27464
rect 1584 27421 1593 27455
rect 1593 27421 1627 27455
rect 1627 27421 1636 27455
rect 1584 27412 1636 27421
rect 23020 27412 23072 27464
rect 23296 27455 23348 27464
rect 23296 27421 23303 27455
rect 23303 27421 23348 27455
rect 23296 27412 23348 27421
rect 1860 27387 1912 27396
rect 1860 27353 1869 27387
rect 1869 27353 1903 27387
rect 1903 27353 1912 27387
rect 1860 27344 1912 27353
rect 23388 27387 23440 27396
rect 23388 27353 23397 27387
rect 23397 27353 23431 27387
rect 23431 27353 23440 27387
rect 23388 27344 23440 27353
rect 31116 27548 31168 27600
rect 33784 27548 33836 27600
rect 57980 27455 58032 27464
rect 57980 27421 57989 27455
rect 57989 27421 58023 27455
rect 58023 27421 58032 27455
rect 57980 27412 58032 27421
rect 22836 27276 22888 27328
rect 58072 27319 58124 27328
rect 58072 27285 58081 27319
rect 58081 27285 58115 27319
rect 58115 27285 58124 27319
rect 58072 27276 58124 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 1584 27072 1636 27124
rect 28356 27072 28408 27124
rect 41696 27072 41748 27124
rect 18880 27004 18932 27056
rect 50988 27004 51040 27056
rect 1584 26979 1636 26988
rect 1584 26945 1593 26979
rect 1593 26945 1627 26979
rect 1627 26945 1636 26979
rect 1584 26936 1636 26945
rect 2504 26979 2556 26988
rect 2504 26945 2513 26979
rect 2513 26945 2547 26979
rect 2547 26945 2556 26979
rect 2504 26936 2556 26945
rect 2596 26979 2648 26988
rect 2596 26945 2606 26979
rect 2606 26945 2640 26979
rect 2640 26945 2648 26979
rect 2596 26936 2648 26945
rect 7840 26936 7892 26988
rect 22836 26979 22888 26988
rect 22836 26945 22845 26979
rect 22845 26945 22879 26979
rect 22879 26945 22888 26979
rect 22836 26936 22888 26945
rect 23204 26936 23256 26988
rect 33140 26936 33192 26988
rect 47492 26936 47544 26988
rect 1768 26911 1820 26920
rect 1768 26877 1777 26911
rect 1777 26877 1811 26911
rect 1811 26877 1820 26911
rect 1768 26868 1820 26877
rect 20720 26868 20772 26920
rect 26884 26868 26936 26920
rect 27804 26868 27856 26920
rect 36636 26868 36688 26920
rect 55864 26868 55916 26920
rect 27252 26800 27304 26852
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 58164 26435 58216 26444
rect 58164 26401 58173 26435
rect 58173 26401 58207 26435
rect 58207 26401 58216 26435
rect 58164 26392 58216 26401
rect 57888 26367 57940 26376
rect 57888 26333 57897 26367
rect 57897 26333 57931 26367
rect 57931 26333 57940 26367
rect 57888 26324 57940 26333
rect 28448 26256 28500 26308
rect 29644 26256 29696 26308
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 1768 25823 1820 25832
rect 1768 25789 1777 25823
rect 1777 25789 1811 25823
rect 1811 25789 1820 25823
rect 1768 25780 1820 25789
rect 9680 25848 9732 25900
rect 10692 25891 10744 25900
rect 10692 25857 10701 25891
rect 10701 25857 10735 25891
rect 10735 25857 10744 25891
rect 10692 25848 10744 25857
rect 17224 25848 17276 25900
rect 58072 25891 58124 25900
rect 58072 25857 58081 25891
rect 58081 25857 58115 25891
rect 58115 25857 58124 25891
rect 58072 25848 58124 25857
rect 18420 25780 18472 25832
rect 34520 25780 34572 25832
rect 23112 25712 23164 25764
rect 40316 25712 40368 25764
rect 23296 25644 23348 25696
rect 48872 25644 48924 25696
rect 57980 25644 58032 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 17224 25440 17276 25492
rect 22560 25440 22612 25492
rect 27436 25440 27488 25492
rect 2504 25279 2556 25288
rect 2504 25245 2513 25279
rect 2513 25245 2547 25279
rect 2547 25245 2556 25279
rect 2504 25236 2556 25245
rect 2596 25279 2648 25288
rect 2596 25245 2606 25279
rect 2606 25245 2640 25279
rect 2640 25245 2648 25279
rect 2596 25236 2648 25245
rect 44456 25236 44508 25288
rect 1860 25211 1912 25220
rect 1860 25177 1869 25211
rect 1869 25177 1903 25211
rect 1903 25177 1912 25211
rect 1860 25168 1912 25177
rect 2872 25168 2924 25220
rect 58164 25211 58216 25220
rect 58164 25177 58173 25211
rect 58173 25177 58207 25211
rect 58207 25177 58216 25211
rect 58164 25168 58216 25177
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 3056 24760 3108 24812
rect 58072 24803 58124 24812
rect 58072 24769 58081 24803
rect 58081 24769 58115 24803
rect 58115 24769 58124 24803
rect 58072 24760 58124 24769
rect 1768 24735 1820 24744
rect 1768 24701 1777 24735
rect 1777 24701 1811 24735
rect 1811 24701 1820 24735
rect 1768 24692 1820 24701
rect 58256 24599 58308 24608
rect 58256 24565 58265 24599
rect 58265 24565 58299 24599
rect 58299 24565 58308 24599
rect 58256 24556 58308 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 3056 24395 3108 24404
rect 3056 24361 3065 24395
rect 3065 24361 3099 24395
rect 3099 24361 3108 24395
rect 3056 24352 3108 24361
rect 4804 24216 4856 24268
rect 32404 24216 32456 24268
rect 1860 24123 1912 24132
rect 1860 24089 1869 24123
rect 1869 24089 1903 24123
rect 1903 24089 1912 24123
rect 1860 24080 1912 24089
rect 2872 24191 2924 24200
rect 2872 24157 2881 24191
rect 2881 24157 2915 24191
rect 2915 24157 2924 24191
rect 2872 24148 2924 24157
rect 30840 24148 30892 24200
rect 12164 24080 12216 24132
rect 13728 24080 13780 24132
rect 26700 24080 26752 24132
rect 26976 24080 27028 24132
rect 54944 24080 54996 24132
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 12808 23783 12860 23792
rect 12808 23749 12817 23783
rect 12817 23749 12851 23783
rect 12851 23749 12860 23783
rect 12808 23740 12860 23749
rect 13728 23672 13780 23724
rect 46296 23536 46348 23588
rect 47860 23536 47912 23588
rect 49516 23536 49568 23588
rect 57520 23536 57572 23588
rect 32496 23468 32548 23520
rect 33140 23468 33192 23520
rect 43628 23468 43680 23520
rect 47584 23468 47636 23520
rect 47676 23468 47728 23520
rect 48596 23468 48648 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 12164 23307 12216 23316
rect 12164 23273 12173 23307
rect 12173 23273 12207 23307
rect 12207 23273 12216 23307
rect 12164 23264 12216 23273
rect 26700 23264 26752 23316
rect 29644 23264 29696 23316
rect 18788 23196 18840 23248
rect 1860 23035 1912 23044
rect 1860 23001 1869 23035
rect 1869 23001 1903 23035
rect 1903 23001 1912 23035
rect 1860 22992 1912 23001
rect 10140 23060 10192 23112
rect 10692 23060 10744 23112
rect 10876 23103 10928 23112
rect 10876 23069 10885 23103
rect 10885 23069 10919 23103
rect 10919 23069 10928 23103
rect 10876 23060 10928 23069
rect 23388 23128 23440 23180
rect 26608 23128 26660 23180
rect 58164 23171 58216 23180
rect 58164 23137 58173 23171
rect 58173 23137 58207 23171
rect 58207 23137 58216 23171
rect 58164 23128 58216 23137
rect 10876 22924 10928 22976
rect 12808 23060 12860 23112
rect 17868 23060 17920 23112
rect 44088 23060 44140 23112
rect 18236 23035 18288 23044
rect 18236 23001 18245 23035
rect 18245 23001 18279 23035
rect 18279 23001 18288 23035
rect 18236 22992 18288 23001
rect 31300 22992 31352 23044
rect 39672 22992 39724 23044
rect 17960 22924 18012 22976
rect 22560 22924 22612 22976
rect 44824 22924 44876 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 18236 22720 18288 22772
rect 9680 22584 9732 22636
rect 1768 22559 1820 22568
rect 1768 22525 1777 22559
rect 1777 22525 1811 22559
rect 1811 22525 1820 22559
rect 1768 22516 1820 22525
rect 16672 22516 16724 22568
rect 17868 22652 17920 22704
rect 24952 22720 25004 22772
rect 17960 22584 18012 22636
rect 18144 22627 18196 22636
rect 18144 22593 18153 22627
rect 18153 22593 18187 22627
rect 18187 22593 18196 22627
rect 18144 22584 18196 22593
rect 18328 22584 18380 22636
rect 21640 22652 21692 22704
rect 48688 22720 48740 22772
rect 58164 22695 58216 22704
rect 58164 22661 58173 22695
rect 58173 22661 58207 22695
rect 58207 22661 58216 22695
rect 58164 22652 58216 22661
rect 24584 22584 24636 22636
rect 16764 22380 16816 22432
rect 25596 22516 25648 22568
rect 19340 22448 19392 22500
rect 20812 22448 20864 22500
rect 24676 22448 24728 22500
rect 20260 22380 20312 22432
rect 24860 22380 24912 22432
rect 41972 22380 42024 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 9680 22219 9732 22228
rect 9680 22185 9689 22219
rect 9689 22185 9723 22219
rect 9723 22185 9732 22219
rect 9680 22176 9732 22185
rect 7288 21972 7340 22024
rect 10140 22040 10192 22092
rect 11060 21972 11112 22024
rect 15936 21972 15988 22024
rect 17132 21972 17184 22024
rect 20996 22108 21048 22160
rect 37280 22108 37332 22160
rect 42432 22108 42484 22160
rect 26148 22083 26200 22092
rect 26148 22049 26157 22083
rect 26157 22049 26191 22083
rect 26191 22049 26200 22083
rect 26148 22040 26200 22049
rect 31208 22040 31260 22092
rect 57336 22040 57388 22092
rect 57704 22040 57756 22092
rect 20996 22015 21048 22024
rect 20996 21981 21005 22015
rect 21005 21981 21039 22015
rect 21039 21981 21048 22015
rect 20996 21972 21048 21981
rect 22008 21972 22060 22024
rect 22100 21972 22152 22024
rect 22836 21972 22888 22024
rect 57060 21972 57112 22024
rect 1860 21947 1912 21956
rect 1860 21913 1869 21947
rect 1869 21913 1903 21947
rect 1903 21913 1912 21947
rect 1860 21904 1912 21913
rect 16396 21904 16448 21956
rect 18144 21904 18196 21956
rect 19432 21904 19484 21956
rect 19708 21904 19760 21956
rect 20260 21904 20312 21956
rect 25044 21904 25096 21956
rect 28632 21904 28684 21956
rect 35992 21904 36044 21956
rect 58164 21947 58216 21956
rect 58164 21913 58173 21947
rect 58173 21913 58207 21947
rect 58207 21913 58216 21947
rect 58164 21904 58216 21913
rect 15384 21836 15436 21888
rect 19800 21879 19852 21888
rect 19800 21845 19809 21879
rect 19809 21845 19843 21879
rect 19843 21845 19852 21879
rect 19800 21836 19852 21845
rect 20168 21879 20220 21888
rect 20168 21845 20177 21879
rect 20177 21845 20211 21879
rect 20211 21845 20220 21879
rect 20168 21836 20220 21845
rect 22100 21836 22152 21888
rect 23848 21836 23900 21888
rect 25872 21836 25924 21888
rect 28540 21836 28592 21888
rect 35808 21836 35860 21888
rect 58992 21836 59044 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 7288 21632 7340 21684
rect 15844 21632 15896 21684
rect 18328 21632 18380 21684
rect 19708 21632 19760 21684
rect 19984 21632 20036 21684
rect 21456 21632 21508 21684
rect 22008 21675 22060 21684
rect 22008 21641 22017 21675
rect 22017 21641 22051 21675
rect 22051 21641 22060 21675
rect 22008 21632 22060 21641
rect 22284 21632 22336 21684
rect 22468 21632 22520 21684
rect 22744 21632 22796 21684
rect 24952 21675 25004 21684
rect 24952 21641 24961 21675
rect 24961 21641 24995 21675
rect 24995 21641 25004 21675
rect 24952 21632 25004 21641
rect 25044 21632 25096 21684
rect 6828 21496 6880 21548
rect 10324 21496 10376 21548
rect 12716 21496 12768 21548
rect 13268 21539 13320 21548
rect 12900 21428 12952 21480
rect 13268 21505 13277 21539
rect 13277 21505 13311 21539
rect 13311 21505 13320 21539
rect 13268 21496 13320 21505
rect 13176 21471 13228 21480
rect 13176 21437 13185 21471
rect 13185 21437 13219 21471
rect 13219 21437 13228 21471
rect 16028 21496 16080 21548
rect 16304 21539 16356 21548
rect 16304 21505 16313 21539
rect 16313 21505 16347 21539
rect 16347 21505 16356 21539
rect 16304 21496 16356 21505
rect 18052 21496 18104 21548
rect 18788 21539 18840 21548
rect 18788 21505 18797 21539
rect 18797 21505 18831 21539
rect 18831 21505 18840 21539
rect 18788 21496 18840 21505
rect 20076 21564 20128 21616
rect 20812 21564 20864 21616
rect 23480 21496 23532 21548
rect 27528 21564 27580 21616
rect 57980 21632 58032 21684
rect 30012 21564 30064 21616
rect 38384 21564 38436 21616
rect 27712 21496 27764 21548
rect 28632 21539 28684 21548
rect 13176 21428 13228 21437
rect 16580 21428 16632 21480
rect 16856 21428 16908 21480
rect 1768 21335 1820 21344
rect 1768 21301 1777 21335
rect 1777 21301 1811 21335
rect 1811 21301 1820 21335
rect 1768 21292 1820 21301
rect 12808 21335 12860 21344
rect 12808 21301 12817 21335
rect 12817 21301 12851 21335
rect 12851 21301 12860 21335
rect 12808 21292 12860 21301
rect 15292 21292 15344 21344
rect 16120 21335 16172 21344
rect 16120 21301 16129 21335
rect 16129 21301 16163 21335
rect 16163 21301 16172 21335
rect 16120 21292 16172 21301
rect 22284 21360 22336 21412
rect 22376 21360 22428 21412
rect 25044 21428 25096 21480
rect 26148 21428 26200 21480
rect 27896 21471 27948 21480
rect 27896 21437 27905 21471
rect 27905 21437 27939 21471
rect 27939 21437 27948 21471
rect 27896 21428 27948 21437
rect 27988 21471 28040 21480
rect 27988 21437 27997 21471
rect 27997 21437 28031 21471
rect 28031 21437 28040 21471
rect 28632 21505 28641 21539
rect 28641 21505 28675 21539
rect 28675 21505 28684 21539
rect 28632 21496 28684 21505
rect 35900 21496 35952 21548
rect 38200 21496 38252 21548
rect 27988 21428 28040 21437
rect 28816 21428 28868 21480
rect 23020 21360 23072 21412
rect 25596 21360 25648 21412
rect 17316 21292 17368 21344
rect 19984 21335 20036 21344
rect 19984 21301 19993 21335
rect 19993 21301 20027 21335
rect 20027 21301 20036 21335
rect 19984 21292 20036 21301
rect 20076 21292 20128 21344
rect 28264 21360 28316 21412
rect 28356 21292 28408 21344
rect 28724 21292 28776 21344
rect 34704 21292 34756 21344
rect 35808 21428 35860 21480
rect 36636 21428 36688 21480
rect 58256 21564 58308 21616
rect 58072 21539 58124 21548
rect 58072 21505 58081 21539
rect 58081 21505 58115 21539
rect 58115 21505 58124 21539
rect 58072 21496 58124 21505
rect 35624 21335 35676 21344
rect 35624 21301 35633 21335
rect 35633 21301 35667 21335
rect 35667 21301 35676 21335
rect 35624 21292 35676 21301
rect 35716 21292 35768 21344
rect 38844 21471 38896 21480
rect 38844 21437 38853 21471
rect 38853 21437 38887 21471
rect 38887 21437 38896 21471
rect 38844 21428 38896 21437
rect 41696 21428 41748 21480
rect 38384 21360 38436 21412
rect 52736 21360 52788 21412
rect 53196 21360 53248 21412
rect 58164 21360 58216 21412
rect 38476 21292 38528 21344
rect 50988 21292 51040 21344
rect 52092 21292 52144 21344
rect 58256 21335 58308 21344
rect 58256 21301 58265 21335
rect 58265 21301 58299 21335
rect 58299 21301 58308 21335
rect 58256 21292 58308 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 15936 21131 15988 21140
rect 15936 21097 15945 21131
rect 15945 21097 15979 21131
rect 15979 21097 15988 21131
rect 15936 21088 15988 21097
rect 16028 21088 16080 21140
rect 12716 21020 12768 21072
rect 11704 20995 11756 21004
rect 11704 20961 11713 20995
rect 11713 20961 11747 20995
rect 11747 20961 11756 20995
rect 11704 20952 11756 20961
rect 12256 20952 12308 21004
rect 11152 20748 11204 20800
rect 12716 20884 12768 20936
rect 13176 20952 13228 21004
rect 13636 20952 13688 21004
rect 16304 21020 16356 21072
rect 27620 21088 27672 21140
rect 27896 21088 27948 21140
rect 28724 21088 28776 21140
rect 32496 21088 32548 21140
rect 58256 21088 58308 21140
rect 15384 20884 15436 20936
rect 16672 20952 16724 21004
rect 17960 20995 18012 21004
rect 17960 20961 17969 20995
rect 17969 20961 18003 20995
rect 18003 20961 18012 20995
rect 17960 20952 18012 20961
rect 19524 20952 19576 21004
rect 15568 20884 15620 20936
rect 15844 20884 15896 20936
rect 16028 20884 16080 20936
rect 16396 20884 16448 20936
rect 16764 20884 16816 20936
rect 17224 20884 17276 20936
rect 20168 20884 20220 20936
rect 22744 20884 22796 20936
rect 23020 20884 23072 20936
rect 23848 20927 23900 20936
rect 23848 20893 23857 20927
rect 23857 20893 23891 20927
rect 23891 20893 23900 20927
rect 23848 20884 23900 20893
rect 26240 20884 26292 20936
rect 27528 20952 27580 21004
rect 27988 20995 28040 21004
rect 27988 20961 27997 20995
rect 27997 20961 28031 20995
rect 28031 20961 28040 20995
rect 27988 20952 28040 20961
rect 28356 20952 28408 21004
rect 13268 20816 13320 20868
rect 12900 20791 12952 20800
rect 12900 20757 12909 20791
rect 12909 20757 12943 20791
rect 12943 20757 12952 20791
rect 12900 20748 12952 20757
rect 13084 20748 13136 20800
rect 15384 20791 15436 20800
rect 15384 20757 15393 20791
rect 15393 20757 15427 20791
rect 15427 20757 15436 20791
rect 15384 20748 15436 20757
rect 19340 20816 19392 20868
rect 18144 20748 18196 20800
rect 20076 20816 20128 20868
rect 19708 20791 19760 20800
rect 19708 20757 19717 20791
rect 19717 20757 19751 20791
rect 19751 20757 19760 20791
rect 19708 20748 19760 20757
rect 20260 20748 20312 20800
rect 23480 20748 23532 20800
rect 25228 20748 25280 20800
rect 25964 20791 26016 20800
rect 25964 20757 25973 20791
rect 25973 20757 26007 20791
rect 26007 20757 26016 20791
rect 25964 20748 26016 20757
rect 26700 20791 26752 20800
rect 26700 20757 26709 20791
rect 26709 20757 26743 20791
rect 26743 20757 26752 20791
rect 26700 20748 26752 20757
rect 26976 20816 27028 20868
rect 27712 20927 27764 20936
rect 27712 20893 27721 20927
rect 27721 20893 27755 20927
rect 27755 20893 27764 20927
rect 27712 20884 27764 20893
rect 29736 20884 29788 20936
rect 53196 21020 53248 21072
rect 30748 20952 30800 21004
rect 31208 20995 31260 21004
rect 31208 20961 31217 20995
rect 31217 20961 31251 20995
rect 31251 20961 31260 20995
rect 31208 20952 31260 20961
rect 35992 20995 36044 21004
rect 35992 20961 36001 20995
rect 36001 20961 36035 20995
rect 36035 20961 36044 20995
rect 35992 20952 36044 20961
rect 37280 20952 37332 21004
rect 41696 20952 41748 21004
rect 52092 20952 52144 21004
rect 34888 20927 34940 20936
rect 34888 20893 34897 20927
rect 34897 20893 34931 20927
rect 34931 20893 34940 20927
rect 34888 20884 34940 20893
rect 38200 20884 38252 20936
rect 38476 20927 38528 20936
rect 38476 20893 38485 20927
rect 38485 20893 38519 20927
rect 38519 20893 38528 20927
rect 38476 20884 38528 20893
rect 41144 20884 41196 20936
rect 42892 20927 42944 20936
rect 42892 20893 42901 20927
rect 42901 20893 42935 20927
rect 42935 20893 42944 20927
rect 42892 20884 42944 20893
rect 42984 20884 43036 20936
rect 44364 20884 44416 20936
rect 47860 20927 47912 20936
rect 47860 20893 47869 20927
rect 47869 20893 47903 20927
rect 47903 20893 47912 20927
rect 47860 20884 47912 20893
rect 52736 20927 52788 20936
rect 52736 20893 52745 20927
rect 52745 20893 52779 20927
rect 52779 20893 52788 20927
rect 52736 20884 52788 20893
rect 53104 20927 53156 20936
rect 36636 20816 36688 20868
rect 38844 20816 38896 20868
rect 42524 20816 42576 20868
rect 28448 20748 28500 20800
rect 28908 20791 28960 20800
rect 28908 20757 28917 20791
rect 28917 20757 28951 20791
rect 28951 20757 28960 20791
rect 28908 20748 28960 20757
rect 30380 20748 30432 20800
rect 31024 20791 31076 20800
rect 31024 20757 31033 20791
rect 31033 20757 31067 20791
rect 31067 20757 31076 20791
rect 31024 20748 31076 20757
rect 31116 20791 31168 20800
rect 31116 20757 31125 20791
rect 31125 20757 31159 20791
rect 31159 20757 31168 20791
rect 31116 20748 31168 20757
rect 31300 20748 31352 20800
rect 32496 20748 32548 20800
rect 38660 20791 38712 20800
rect 38660 20757 38669 20791
rect 38669 20757 38703 20791
rect 38703 20757 38712 20791
rect 38660 20748 38712 20757
rect 41420 20748 41472 20800
rect 41972 20791 42024 20800
rect 41972 20757 41981 20791
rect 41981 20757 42015 20791
rect 42015 20757 42024 20791
rect 43076 20791 43128 20800
rect 41972 20748 42024 20757
rect 43076 20757 43085 20791
rect 43085 20757 43119 20791
rect 43119 20757 43128 20791
rect 43076 20748 43128 20757
rect 43444 20816 43496 20868
rect 47676 20859 47728 20868
rect 47676 20825 47685 20859
rect 47685 20825 47719 20859
rect 47719 20825 47728 20859
rect 47676 20816 47728 20825
rect 49148 20816 49200 20868
rect 50712 20816 50764 20868
rect 53104 20893 53113 20927
rect 53113 20893 53147 20927
rect 53147 20893 53156 20927
rect 53104 20884 53156 20893
rect 54116 20995 54168 21004
rect 54116 20961 54125 20995
rect 54125 20961 54159 20995
rect 54159 20961 54168 20995
rect 54116 20952 54168 20961
rect 55312 20952 55364 21004
rect 54484 20884 54536 20936
rect 54760 20927 54812 20936
rect 54760 20893 54769 20927
rect 54769 20893 54803 20927
rect 54803 20893 54812 20927
rect 54760 20884 54812 20893
rect 54852 20884 54904 20936
rect 56048 20884 56100 20936
rect 48228 20748 48280 20800
rect 55680 20816 55732 20868
rect 58164 20859 58216 20868
rect 58164 20825 58173 20859
rect 58173 20825 58207 20859
rect 58207 20825 58216 20859
rect 58164 20816 58216 20825
rect 55220 20748 55272 20800
rect 56692 20748 56744 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 12900 20544 12952 20596
rect 18880 20544 18932 20596
rect 19340 20544 19392 20596
rect 19800 20544 19852 20596
rect 27712 20544 27764 20596
rect 28172 20544 28224 20596
rect 7380 20408 7432 20460
rect 8024 20451 8076 20460
rect 8024 20417 8033 20451
rect 8033 20417 8067 20451
rect 8067 20417 8076 20451
rect 8024 20408 8076 20417
rect 11704 20476 11756 20528
rect 11152 20451 11204 20460
rect 11152 20417 11161 20451
rect 11161 20417 11195 20451
rect 11195 20417 11204 20451
rect 11152 20408 11204 20417
rect 13360 20408 13412 20460
rect 1768 20383 1820 20392
rect 1768 20349 1777 20383
rect 1777 20349 1811 20383
rect 1811 20349 1820 20383
rect 1768 20340 1820 20349
rect 11888 20340 11940 20392
rect 15384 20408 15436 20460
rect 16672 20408 16724 20460
rect 17868 20451 17920 20460
rect 17868 20417 17877 20451
rect 17877 20417 17911 20451
rect 17911 20417 17920 20451
rect 17868 20408 17920 20417
rect 22100 20476 22152 20528
rect 26700 20476 26752 20528
rect 18512 20451 18564 20460
rect 15844 20340 15896 20392
rect 17224 20340 17276 20392
rect 18512 20417 18521 20451
rect 18521 20417 18555 20451
rect 18555 20417 18564 20451
rect 18512 20408 18564 20417
rect 19340 20408 19392 20460
rect 21456 20451 21508 20460
rect 21456 20417 21465 20451
rect 21465 20417 21499 20451
rect 21499 20417 21508 20451
rect 21456 20408 21508 20417
rect 24308 20451 24360 20460
rect 19432 20340 19484 20392
rect 13636 20272 13688 20324
rect 9404 20247 9456 20256
rect 9404 20213 9413 20247
rect 9413 20213 9447 20247
rect 9447 20213 9456 20247
rect 9404 20204 9456 20213
rect 11060 20247 11112 20256
rect 11060 20213 11069 20247
rect 11069 20213 11103 20247
rect 11103 20213 11112 20247
rect 11060 20204 11112 20213
rect 15200 20247 15252 20256
rect 15200 20213 15209 20247
rect 15209 20213 15243 20247
rect 15243 20213 15252 20247
rect 15200 20204 15252 20213
rect 16580 20204 16632 20256
rect 17592 20272 17644 20324
rect 22008 20383 22060 20392
rect 22008 20349 22017 20383
rect 22017 20349 22051 20383
rect 22051 20349 22060 20383
rect 22008 20340 22060 20349
rect 24308 20417 24317 20451
rect 24317 20417 24351 20451
rect 24351 20417 24360 20451
rect 24308 20408 24360 20417
rect 26240 20408 26292 20460
rect 27160 20451 27212 20460
rect 27160 20417 27169 20451
rect 27169 20417 27203 20451
rect 27203 20417 27212 20451
rect 27160 20408 27212 20417
rect 25320 20340 25372 20392
rect 25504 20340 25556 20392
rect 34888 20476 34940 20528
rect 39948 20544 40000 20596
rect 43904 20544 43956 20596
rect 44088 20587 44140 20596
rect 44088 20553 44097 20587
rect 44097 20553 44131 20587
rect 44131 20553 44140 20587
rect 44088 20544 44140 20553
rect 49148 20544 49200 20596
rect 54484 20587 54536 20596
rect 54484 20553 54493 20587
rect 54493 20553 54527 20587
rect 54527 20553 54536 20587
rect 54484 20544 54536 20553
rect 56600 20544 56652 20596
rect 57888 20544 57940 20596
rect 42524 20476 42576 20528
rect 43076 20476 43128 20528
rect 43536 20476 43588 20528
rect 34612 20408 34664 20460
rect 36084 20408 36136 20460
rect 38752 20408 38804 20460
rect 41420 20451 41472 20460
rect 41420 20417 41429 20451
rect 41429 20417 41463 20451
rect 41463 20417 41472 20451
rect 41420 20408 41472 20417
rect 19800 20204 19852 20256
rect 20076 20204 20128 20256
rect 23204 20204 23256 20256
rect 24216 20204 24268 20256
rect 28264 20272 28316 20324
rect 29736 20204 29788 20256
rect 32496 20272 32548 20324
rect 35348 20340 35400 20392
rect 35808 20340 35860 20392
rect 37280 20340 37332 20392
rect 38660 20383 38712 20392
rect 38660 20349 38669 20383
rect 38669 20349 38703 20383
rect 38703 20349 38712 20383
rect 38660 20340 38712 20349
rect 41144 20340 41196 20392
rect 44364 20408 44416 20460
rect 47032 20451 47084 20460
rect 47032 20417 47041 20451
rect 47041 20417 47075 20451
rect 47075 20417 47084 20451
rect 47032 20408 47084 20417
rect 48412 20451 48464 20460
rect 48412 20417 48446 20451
rect 48446 20417 48464 20451
rect 51448 20476 51500 20528
rect 48412 20408 48464 20417
rect 50528 20451 50580 20460
rect 50528 20417 50562 20451
rect 50562 20417 50580 20451
rect 50528 20408 50580 20417
rect 54116 20408 54168 20460
rect 56508 20476 56560 20528
rect 55220 20451 55272 20460
rect 55220 20417 55254 20451
rect 55254 20417 55272 20451
rect 55220 20408 55272 20417
rect 42708 20383 42760 20392
rect 39672 20272 39724 20324
rect 42708 20349 42717 20383
rect 42717 20349 42751 20383
rect 42751 20349 42760 20383
rect 42708 20340 42760 20349
rect 46848 20383 46900 20392
rect 46848 20349 46857 20383
rect 46857 20349 46891 20383
rect 46891 20349 46900 20383
rect 46848 20340 46900 20349
rect 48136 20383 48188 20392
rect 48136 20349 48145 20383
rect 48145 20349 48179 20383
rect 48179 20349 48188 20383
rect 48136 20340 48188 20349
rect 33692 20247 33744 20256
rect 33692 20213 33701 20247
rect 33701 20213 33735 20247
rect 33735 20213 33744 20247
rect 33692 20204 33744 20213
rect 35900 20204 35952 20256
rect 37832 20247 37884 20256
rect 37832 20213 37841 20247
rect 37841 20213 37875 20247
rect 37875 20213 37884 20247
rect 37832 20204 37884 20213
rect 38200 20204 38252 20256
rect 39764 20247 39816 20256
rect 39764 20213 39773 20247
rect 39773 20213 39807 20247
rect 39807 20213 39816 20247
rect 39764 20204 39816 20213
rect 40224 20204 40276 20256
rect 41604 20247 41656 20256
rect 41604 20213 41613 20247
rect 41613 20213 41647 20247
rect 41647 20213 41656 20247
rect 41604 20204 41656 20213
rect 45284 20272 45336 20324
rect 51632 20315 51684 20324
rect 43444 20204 43496 20256
rect 43812 20204 43864 20256
rect 47216 20247 47268 20256
rect 47216 20213 47225 20247
rect 47225 20213 47259 20247
rect 47259 20213 47268 20247
rect 47216 20204 47268 20213
rect 51632 20281 51641 20315
rect 51641 20281 51675 20315
rect 51675 20281 51684 20315
rect 51632 20272 51684 20281
rect 50988 20204 51040 20256
rect 53104 20204 53156 20256
rect 54392 20204 54444 20256
rect 55864 20204 55916 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 13636 20000 13688 20052
rect 14924 20000 14976 20052
rect 9404 19975 9456 19984
rect 9404 19941 9413 19975
rect 9413 19941 9447 19975
rect 9447 19941 9456 19975
rect 9404 19932 9456 19941
rect 20812 20043 20864 20052
rect 19156 19932 19208 19984
rect 13176 19907 13228 19916
rect 9312 19796 9364 19848
rect 13176 19873 13185 19907
rect 13185 19873 13219 19907
rect 13219 19873 13228 19907
rect 13176 19864 13228 19873
rect 20812 20009 20821 20043
rect 20821 20009 20855 20043
rect 20855 20009 20864 20043
rect 20812 20000 20864 20009
rect 22744 20043 22796 20052
rect 22744 20009 22753 20043
rect 22753 20009 22787 20043
rect 22787 20009 22796 20043
rect 22744 20000 22796 20009
rect 24308 20000 24360 20052
rect 35348 20043 35400 20052
rect 35348 20009 35357 20043
rect 35357 20009 35391 20043
rect 35391 20009 35400 20043
rect 35348 20000 35400 20009
rect 21456 19932 21508 19984
rect 25412 19932 25464 19984
rect 1860 19771 1912 19780
rect 1860 19737 1869 19771
rect 1869 19737 1903 19771
rect 1903 19737 1912 19771
rect 1860 19728 1912 19737
rect 9588 19728 9640 19780
rect 12808 19796 12860 19848
rect 14648 19839 14700 19848
rect 14648 19805 14657 19839
rect 14657 19805 14691 19839
rect 14691 19805 14700 19839
rect 14648 19796 14700 19805
rect 15200 19796 15252 19848
rect 7472 19703 7524 19712
rect 7472 19669 7481 19703
rect 7481 19669 7515 19703
rect 7515 19669 7524 19703
rect 7472 19660 7524 19669
rect 9220 19660 9272 19712
rect 10692 19703 10744 19712
rect 10692 19669 10701 19703
rect 10701 19669 10735 19703
rect 10735 19669 10744 19703
rect 10692 19660 10744 19669
rect 16856 19796 16908 19848
rect 25504 19864 25556 19916
rect 35808 19932 35860 19984
rect 39672 19932 39724 19984
rect 42524 19975 42576 19984
rect 42524 19941 42533 19975
rect 42533 19941 42567 19975
rect 42567 19941 42576 19975
rect 42524 19932 42576 19941
rect 44456 19975 44508 19984
rect 44456 19941 44465 19975
rect 44465 19941 44499 19975
rect 44499 19941 44508 19975
rect 44456 19932 44508 19941
rect 48412 19975 48464 19984
rect 48412 19941 48421 19975
rect 48421 19941 48455 19975
rect 48455 19941 48464 19975
rect 48412 19932 48464 19941
rect 54760 20000 54812 20052
rect 56048 20043 56100 20052
rect 56048 20009 56057 20043
rect 56057 20009 56091 20043
rect 56091 20009 56100 20043
rect 56048 20000 56100 20009
rect 27620 19907 27672 19916
rect 27620 19873 27629 19907
rect 27629 19873 27663 19907
rect 27663 19873 27672 19907
rect 27620 19864 27672 19873
rect 38292 19907 38344 19916
rect 38292 19873 38301 19907
rect 38301 19873 38335 19907
rect 38335 19873 38344 19907
rect 38292 19864 38344 19873
rect 47676 19864 47728 19916
rect 20812 19796 20864 19848
rect 22284 19796 22336 19848
rect 23204 19796 23256 19848
rect 22192 19728 22244 19780
rect 23112 19728 23164 19780
rect 19340 19660 19392 19712
rect 20168 19660 20220 19712
rect 23756 19660 23808 19712
rect 24952 19839 25004 19848
rect 24952 19805 24961 19839
rect 24961 19805 24995 19839
rect 24995 19805 25004 19839
rect 24952 19796 25004 19805
rect 25320 19796 25372 19848
rect 29736 19839 29788 19848
rect 25872 19728 25924 19780
rect 29736 19805 29745 19839
rect 29745 19805 29779 19839
rect 29779 19805 29788 19839
rect 29736 19796 29788 19805
rect 30472 19796 30524 19848
rect 30656 19839 30708 19848
rect 30656 19805 30665 19839
rect 30665 19805 30699 19839
rect 30699 19805 30708 19839
rect 30656 19796 30708 19805
rect 35624 19796 35676 19848
rect 38752 19796 38804 19848
rect 42708 19796 42760 19848
rect 45376 19796 45428 19848
rect 47216 19796 47268 19848
rect 48228 19839 48280 19848
rect 24952 19660 25004 19712
rect 30564 19660 30616 19712
rect 35900 19728 35952 19780
rect 37832 19728 37884 19780
rect 38292 19728 38344 19780
rect 40224 19728 40276 19780
rect 36360 19660 36412 19712
rect 38660 19660 38712 19712
rect 39764 19660 39816 19712
rect 41604 19728 41656 19780
rect 42156 19728 42208 19780
rect 45284 19771 45336 19780
rect 45284 19737 45293 19771
rect 45293 19737 45327 19771
rect 45327 19737 45336 19771
rect 45284 19728 45336 19737
rect 45560 19728 45612 19780
rect 46848 19728 46900 19780
rect 48228 19805 48237 19839
rect 48237 19805 48271 19839
rect 48271 19805 48280 19839
rect 48228 19796 48280 19805
rect 48320 19728 48372 19780
rect 49700 19796 49752 19848
rect 51080 19864 51132 19916
rect 51448 19907 51500 19916
rect 51448 19873 51457 19907
rect 51457 19873 51491 19907
rect 51491 19873 51500 19907
rect 51448 19864 51500 19873
rect 50712 19839 50764 19848
rect 50712 19805 50721 19839
rect 50721 19805 50755 19839
rect 50755 19805 50764 19839
rect 50712 19796 50764 19805
rect 53840 19839 53892 19848
rect 42800 19660 42852 19712
rect 43076 19660 43128 19712
rect 43720 19660 43772 19712
rect 46296 19660 46348 19712
rect 49516 19660 49568 19712
rect 49976 19660 50028 19712
rect 52276 19728 52328 19780
rect 53840 19805 53849 19839
rect 53849 19805 53883 19839
rect 53883 19805 53892 19839
rect 53840 19796 53892 19805
rect 54576 19864 54628 19916
rect 54300 19796 54352 19848
rect 56508 19864 56560 19916
rect 55680 19839 55732 19848
rect 55680 19805 55689 19839
rect 55689 19805 55723 19839
rect 55723 19805 55732 19839
rect 55680 19796 55732 19805
rect 55864 19839 55916 19848
rect 55864 19805 55873 19839
rect 55873 19805 55907 19839
rect 55907 19805 55916 19839
rect 55864 19796 55916 19805
rect 56692 19796 56744 19848
rect 50712 19660 50764 19712
rect 51264 19660 51316 19712
rect 54668 19660 54720 19712
rect 56140 19728 56192 19780
rect 56600 19660 56652 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 7472 19388 7524 19440
rect 30656 19456 30708 19508
rect 33784 19456 33836 19508
rect 34612 19499 34664 19508
rect 1860 19363 1912 19372
rect 1860 19329 1869 19363
rect 1869 19329 1903 19363
rect 1903 19329 1912 19363
rect 1860 19320 1912 19329
rect 6828 19363 6880 19372
rect 6828 19329 6837 19363
rect 6837 19329 6871 19363
rect 6871 19329 6880 19363
rect 6828 19320 6880 19329
rect 10692 19320 10744 19372
rect 11888 19363 11940 19372
rect 11888 19329 11897 19363
rect 11897 19329 11931 19363
rect 11931 19329 11940 19363
rect 11888 19320 11940 19329
rect 12164 19295 12216 19304
rect 12164 19261 12173 19295
rect 12173 19261 12207 19295
rect 12207 19261 12216 19295
rect 12164 19252 12216 19261
rect 15292 19320 15344 19372
rect 16856 19363 16908 19372
rect 16856 19329 16865 19363
rect 16865 19329 16899 19363
rect 16899 19329 16908 19363
rect 16856 19320 16908 19329
rect 17776 19320 17828 19372
rect 19156 19363 19208 19372
rect 19156 19329 19165 19363
rect 19165 19329 19199 19363
rect 19199 19329 19208 19363
rect 19156 19320 19208 19329
rect 20168 19320 20220 19372
rect 22008 19320 22060 19372
rect 24860 19388 24912 19440
rect 25596 19388 25648 19440
rect 30012 19388 30064 19440
rect 24216 19320 24268 19372
rect 24308 19363 24360 19372
rect 24308 19329 24317 19363
rect 24317 19329 24351 19363
rect 24351 19329 24360 19363
rect 24308 19320 24360 19329
rect 26976 19320 27028 19372
rect 30288 19363 30340 19372
rect 14648 19252 14700 19304
rect 17960 19252 18012 19304
rect 20720 19295 20772 19304
rect 20720 19261 20729 19295
rect 20729 19261 20763 19295
rect 20763 19261 20772 19295
rect 20720 19252 20772 19261
rect 25412 19295 25464 19304
rect 25412 19261 25421 19295
rect 25421 19261 25455 19295
rect 25455 19261 25464 19295
rect 25412 19252 25464 19261
rect 2412 19159 2464 19168
rect 2412 19125 2421 19159
rect 2421 19125 2455 19159
rect 2455 19125 2464 19159
rect 2412 19116 2464 19125
rect 10048 19159 10100 19168
rect 10048 19125 10057 19159
rect 10057 19125 10091 19159
rect 10091 19125 10100 19159
rect 10048 19116 10100 19125
rect 15200 19159 15252 19168
rect 15200 19125 15209 19159
rect 15209 19125 15243 19159
rect 15243 19125 15252 19159
rect 15200 19116 15252 19125
rect 16028 19116 16080 19168
rect 21456 19184 21508 19236
rect 17868 19116 17920 19168
rect 23480 19184 23532 19236
rect 23756 19227 23808 19236
rect 23756 19193 23765 19227
rect 23765 19193 23799 19227
rect 23799 19193 23808 19227
rect 23756 19184 23808 19193
rect 30288 19329 30297 19363
rect 30297 19329 30331 19363
rect 30331 19329 30340 19363
rect 30288 19320 30340 19329
rect 30380 19320 30432 19372
rect 33692 19388 33744 19440
rect 34612 19465 34621 19499
rect 34621 19465 34655 19499
rect 34655 19465 34664 19499
rect 34612 19456 34664 19465
rect 35072 19499 35124 19508
rect 35072 19465 35081 19499
rect 35081 19465 35115 19499
rect 35115 19465 35124 19499
rect 35072 19456 35124 19465
rect 36084 19456 36136 19508
rect 36360 19499 36412 19508
rect 36360 19465 36369 19499
rect 36369 19465 36403 19499
rect 36403 19465 36412 19499
rect 36360 19456 36412 19465
rect 36452 19499 36504 19508
rect 36452 19465 36461 19499
rect 36461 19465 36495 19499
rect 36495 19465 36504 19499
rect 36452 19456 36504 19465
rect 59176 19456 59228 19508
rect 32496 19363 32548 19372
rect 32496 19329 32505 19363
rect 32505 19329 32539 19363
rect 32539 19329 32548 19363
rect 32496 19320 32548 19329
rect 33140 19320 33192 19372
rect 39948 19320 40000 19372
rect 40776 19320 40828 19372
rect 43720 19388 43772 19440
rect 43904 19388 43956 19440
rect 51172 19431 51224 19440
rect 42800 19363 42852 19372
rect 42800 19329 42809 19363
rect 42809 19329 42843 19363
rect 42843 19329 42852 19363
rect 42800 19320 42852 19329
rect 34704 19252 34756 19304
rect 35072 19252 35124 19304
rect 36636 19295 36688 19304
rect 36636 19261 36645 19295
rect 36645 19261 36679 19295
rect 36679 19261 36688 19295
rect 36636 19252 36688 19261
rect 37280 19252 37332 19304
rect 31668 19227 31720 19236
rect 23388 19116 23440 19168
rect 26056 19116 26108 19168
rect 28356 19159 28408 19168
rect 28356 19125 28365 19159
rect 28365 19125 28399 19159
rect 28399 19125 28408 19159
rect 28356 19116 28408 19125
rect 31024 19116 31076 19168
rect 31668 19193 31677 19227
rect 31677 19193 31711 19227
rect 31711 19193 31720 19227
rect 31668 19184 31720 19193
rect 33692 19184 33744 19236
rect 42248 19184 42300 19236
rect 35716 19159 35768 19168
rect 35716 19125 35725 19159
rect 35725 19125 35759 19159
rect 35759 19125 35768 19159
rect 35716 19116 35768 19125
rect 36452 19116 36504 19168
rect 41880 19116 41932 19168
rect 42156 19116 42208 19168
rect 43168 19320 43220 19372
rect 45376 19363 45428 19372
rect 45376 19329 45385 19363
rect 45385 19329 45419 19363
rect 45419 19329 45428 19363
rect 45376 19320 45428 19329
rect 45652 19363 45704 19372
rect 45652 19329 45686 19363
rect 45686 19329 45704 19363
rect 45652 19320 45704 19329
rect 47584 19320 47636 19372
rect 47860 19320 47912 19372
rect 48228 19320 48280 19372
rect 50160 19320 50212 19372
rect 50712 19320 50764 19372
rect 51172 19397 51181 19431
rect 51181 19397 51215 19431
rect 51215 19397 51224 19431
rect 51172 19388 51224 19397
rect 51080 19363 51132 19372
rect 51080 19329 51089 19363
rect 51089 19329 51123 19363
rect 51123 19329 51132 19363
rect 51080 19320 51132 19329
rect 52460 19388 52512 19440
rect 54300 19388 54352 19440
rect 44456 19252 44508 19304
rect 48320 19252 48372 19304
rect 51356 19252 51408 19304
rect 46388 19184 46440 19236
rect 52276 19363 52328 19372
rect 52276 19329 52285 19363
rect 52285 19329 52319 19363
rect 52319 19329 52328 19363
rect 52276 19320 52328 19329
rect 51540 19252 51592 19304
rect 43260 19116 43312 19168
rect 43904 19159 43956 19168
rect 43904 19125 43913 19159
rect 43913 19125 43947 19159
rect 43947 19125 43956 19159
rect 43904 19116 43956 19125
rect 46664 19116 46716 19168
rect 46940 19116 46992 19168
rect 47676 19116 47728 19168
rect 50620 19116 50672 19168
rect 58072 19116 58124 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 12164 18912 12216 18964
rect 22100 18912 22152 18964
rect 17592 18844 17644 18896
rect 16396 18776 16448 18828
rect 19432 18844 19484 18896
rect 20812 18844 20864 18896
rect 18052 18819 18104 18828
rect 18052 18785 18061 18819
rect 18061 18785 18095 18819
rect 18095 18785 18104 18819
rect 18052 18776 18104 18785
rect 1860 18683 1912 18692
rect 1860 18649 1869 18683
rect 1869 18649 1903 18683
rect 1903 18649 1912 18683
rect 1860 18640 1912 18649
rect 2412 18683 2464 18692
rect 2412 18649 2421 18683
rect 2421 18649 2455 18683
rect 2455 18649 2464 18683
rect 2412 18640 2464 18649
rect 6828 18708 6880 18760
rect 8208 18708 8260 18760
rect 13728 18708 13780 18760
rect 14556 18708 14608 18760
rect 15200 18708 15252 18760
rect 16580 18751 16632 18760
rect 16580 18717 16589 18751
rect 16589 18717 16623 18751
rect 16623 18717 16632 18751
rect 16580 18708 16632 18717
rect 7012 18640 7064 18692
rect 9680 18640 9732 18692
rect 12348 18640 12400 18692
rect 7104 18572 7156 18624
rect 20996 18640 21048 18692
rect 28356 18912 28408 18964
rect 26700 18844 26752 18896
rect 27068 18844 27120 18896
rect 36452 18912 36504 18964
rect 37004 18912 37056 18964
rect 26056 18776 26108 18828
rect 28264 18776 28316 18828
rect 28356 18819 28408 18828
rect 28356 18785 28365 18819
rect 28365 18785 28399 18819
rect 28399 18785 28408 18819
rect 28356 18776 28408 18785
rect 29460 18776 29512 18828
rect 30288 18819 30340 18828
rect 30288 18785 30297 18819
rect 30297 18785 30331 18819
rect 30331 18785 30340 18819
rect 30288 18776 30340 18785
rect 23480 18708 23532 18760
rect 24768 18751 24820 18760
rect 24768 18717 24777 18751
rect 24777 18717 24811 18751
rect 24811 18717 24820 18751
rect 24768 18708 24820 18717
rect 25780 18751 25832 18760
rect 25780 18717 25789 18751
rect 25789 18717 25823 18751
rect 25823 18717 25832 18751
rect 25780 18708 25832 18717
rect 26516 18751 26568 18760
rect 26516 18717 26525 18751
rect 26525 18717 26559 18751
rect 26559 18717 26568 18751
rect 26516 18708 26568 18717
rect 30012 18708 30064 18760
rect 30564 18751 30616 18760
rect 30564 18717 30598 18751
rect 30598 18717 30616 18751
rect 30564 18708 30616 18717
rect 22008 18640 22060 18692
rect 22192 18640 22244 18692
rect 28356 18640 28408 18692
rect 28632 18640 28684 18692
rect 30656 18640 30708 18692
rect 33692 18844 33744 18896
rect 35716 18887 35768 18896
rect 35716 18853 35725 18887
rect 35725 18853 35759 18887
rect 35759 18853 35768 18887
rect 35716 18844 35768 18853
rect 36360 18887 36412 18896
rect 36360 18853 36369 18887
rect 36369 18853 36403 18887
rect 36403 18853 36412 18887
rect 36360 18844 36412 18853
rect 42616 18844 42668 18896
rect 42892 18844 42944 18896
rect 31484 18776 31536 18828
rect 31760 18776 31812 18828
rect 38292 18776 38344 18828
rect 40040 18776 40092 18828
rect 31668 18708 31720 18760
rect 22284 18572 22336 18624
rect 23388 18572 23440 18624
rect 26792 18572 26844 18624
rect 26884 18572 26936 18624
rect 31392 18640 31444 18692
rect 33692 18640 33744 18692
rect 35900 18708 35952 18760
rect 38844 18751 38896 18760
rect 38844 18717 38853 18751
rect 38853 18717 38887 18751
rect 38887 18717 38896 18751
rect 38844 18708 38896 18717
rect 42248 18776 42300 18828
rect 36728 18640 36780 18692
rect 38384 18640 38436 18692
rect 39212 18640 39264 18692
rect 42892 18711 42902 18738
rect 42902 18711 42936 18738
rect 42936 18711 42944 18738
rect 42892 18686 42944 18711
rect 43260 18844 43312 18896
rect 45284 18844 45336 18896
rect 45652 18912 45704 18964
rect 47032 18912 47084 18964
rect 58072 18955 58124 18964
rect 58072 18921 58081 18955
rect 58081 18921 58115 18955
rect 58115 18921 58124 18955
rect 58072 18912 58124 18921
rect 53840 18844 53892 18896
rect 44088 18776 44140 18828
rect 43628 18708 43680 18760
rect 53932 18776 53984 18828
rect 55036 18776 55088 18828
rect 31208 18572 31260 18624
rect 33048 18572 33100 18624
rect 34520 18572 34572 18624
rect 35440 18572 35492 18624
rect 37188 18572 37240 18624
rect 39028 18615 39080 18624
rect 39028 18581 39037 18615
rect 39037 18581 39071 18615
rect 39071 18581 39080 18615
rect 39028 18572 39080 18581
rect 40592 18615 40644 18624
rect 40592 18581 40601 18615
rect 40601 18581 40635 18615
rect 40635 18581 40644 18615
rect 40592 18572 40644 18581
rect 40960 18615 41012 18624
rect 40960 18581 40969 18615
rect 40969 18581 41003 18615
rect 41003 18581 41012 18615
rect 40960 18572 41012 18581
rect 41880 18572 41932 18624
rect 43168 18640 43220 18692
rect 43720 18640 43772 18692
rect 45928 18708 45980 18760
rect 46020 18751 46072 18760
rect 46020 18717 46029 18751
rect 46029 18717 46063 18751
rect 46063 18717 46072 18751
rect 46296 18751 46348 18760
rect 46020 18708 46072 18717
rect 46296 18717 46305 18751
rect 46305 18717 46339 18751
rect 46339 18717 46348 18751
rect 46296 18708 46348 18717
rect 46388 18751 46440 18760
rect 46388 18717 46397 18751
rect 46397 18717 46431 18751
rect 46431 18717 46440 18751
rect 46388 18708 46440 18717
rect 47860 18708 47912 18760
rect 48320 18751 48372 18760
rect 48320 18717 48329 18751
rect 48329 18717 48363 18751
rect 48363 18717 48372 18751
rect 48320 18708 48372 18717
rect 48504 18751 48556 18760
rect 48504 18717 48513 18751
rect 48513 18717 48547 18751
rect 48547 18717 48556 18751
rect 48504 18708 48556 18717
rect 51356 18708 51408 18760
rect 55312 18708 55364 18760
rect 45560 18640 45612 18692
rect 45284 18572 45336 18624
rect 46756 18640 46808 18692
rect 46848 18640 46900 18692
rect 47584 18640 47636 18692
rect 45836 18572 45888 18624
rect 49700 18640 49752 18692
rect 53840 18640 53892 18692
rect 58440 18776 58492 18828
rect 56600 18708 56652 18760
rect 57980 18751 58032 18760
rect 57980 18717 57989 18751
rect 57989 18717 58023 18751
rect 58023 18717 58032 18751
rect 57980 18708 58032 18717
rect 57244 18683 57296 18692
rect 57244 18649 57253 18683
rect 57253 18649 57287 18683
rect 57287 18649 57296 18683
rect 57244 18640 57296 18649
rect 48780 18572 48832 18624
rect 55864 18615 55916 18624
rect 55864 18581 55873 18615
rect 55873 18581 55907 18615
rect 55907 18581 55916 18615
rect 55864 18572 55916 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 6828 18368 6880 18420
rect 20904 18368 20956 18420
rect 20996 18368 21048 18420
rect 22100 18368 22152 18420
rect 7104 18232 7156 18284
rect 8116 18232 8168 18284
rect 12716 18300 12768 18352
rect 17868 18300 17920 18352
rect 12256 18232 12308 18284
rect 16028 18275 16080 18284
rect 16028 18241 16037 18275
rect 16037 18241 16071 18275
rect 16071 18241 16080 18275
rect 16028 18232 16080 18241
rect 16396 18232 16448 18284
rect 16856 18232 16908 18284
rect 22192 18300 22244 18352
rect 22376 18343 22428 18352
rect 22376 18309 22385 18343
rect 22385 18309 22419 18343
rect 22419 18309 22428 18343
rect 22376 18300 22428 18309
rect 23572 18368 23624 18420
rect 24308 18368 24360 18420
rect 28816 18368 28868 18420
rect 30472 18368 30524 18420
rect 40960 18368 41012 18420
rect 26976 18300 27028 18352
rect 28908 18300 28960 18352
rect 41788 18343 41840 18352
rect 11060 18164 11112 18216
rect 19248 18232 19300 18284
rect 21640 18232 21692 18284
rect 22284 18232 22336 18284
rect 23572 18275 23624 18284
rect 23572 18241 23581 18275
rect 23581 18241 23615 18275
rect 23615 18241 23624 18275
rect 23572 18232 23624 18241
rect 19432 18164 19484 18216
rect 23296 18164 23348 18216
rect 23480 18164 23532 18216
rect 24768 18232 24820 18284
rect 27068 18232 27120 18284
rect 27160 18232 27212 18284
rect 28264 18232 28316 18284
rect 29552 18232 29604 18284
rect 29828 18275 29880 18284
rect 29828 18241 29837 18275
rect 29837 18241 29871 18275
rect 29871 18241 29880 18275
rect 29828 18232 29880 18241
rect 31208 18275 31260 18284
rect 12532 18096 12584 18148
rect 9772 18071 9824 18080
rect 9772 18037 9781 18071
rect 9781 18037 9815 18071
rect 9815 18037 9824 18071
rect 9772 18028 9824 18037
rect 13452 18028 13504 18080
rect 16028 18028 16080 18080
rect 16212 18028 16264 18080
rect 16396 18028 16448 18080
rect 23388 18096 23440 18148
rect 26240 18096 26292 18148
rect 27160 18096 27212 18148
rect 23572 18028 23624 18080
rect 26516 18028 26568 18080
rect 29920 18164 29972 18216
rect 31208 18241 31217 18275
rect 31217 18241 31251 18275
rect 31251 18241 31260 18275
rect 31208 18232 31260 18241
rect 32128 18275 32180 18284
rect 32128 18241 32137 18275
rect 32137 18241 32171 18275
rect 32171 18241 32180 18275
rect 32128 18232 32180 18241
rect 33876 18232 33928 18284
rect 34704 18275 34756 18284
rect 34704 18241 34713 18275
rect 34713 18241 34747 18275
rect 34747 18241 34756 18275
rect 34704 18232 34756 18241
rect 38752 18275 38804 18284
rect 38752 18241 38761 18275
rect 38761 18241 38795 18275
rect 38795 18241 38804 18275
rect 38752 18232 38804 18241
rect 30196 18164 30248 18216
rect 31668 18164 31720 18216
rect 35348 18164 35400 18216
rect 35624 18164 35676 18216
rect 38384 18164 38436 18216
rect 39028 18275 39080 18284
rect 39028 18241 39037 18275
rect 39037 18241 39071 18275
rect 39071 18241 39080 18275
rect 39028 18232 39080 18241
rect 33968 18096 34020 18148
rect 28816 18028 28868 18080
rect 29920 18028 29972 18080
rect 30012 18028 30064 18080
rect 33784 18028 33836 18080
rect 34428 18028 34480 18080
rect 36636 18028 36688 18080
rect 39028 18028 39080 18080
rect 40040 18028 40092 18080
rect 40960 18028 41012 18080
rect 41788 18309 41797 18343
rect 41797 18309 41831 18343
rect 41831 18309 41840 18343
rect 41788 18300 41840 18309
rect 42432 18300 42484 18352
rect 42616 18368 42668 18420
rect 45836 18368 45888 18420
rect 45928 18368 45980 18420
rect 46572 18368 46624 18420
rect 53840 18368 53892 18420
rect 53932 18368 53984 18420
rect 42800 18300 42852 18352
rect 45284 18300 45336 18352
rect 46664 18300 46716 18352
rect 46940 18300 46992 18352
rect 50068 18300 50120 18352
rect 42708 18275 42760 18284
rect 42708 18241 42718 18275
rect 42718 18241 42752 18275
rect 42752 18241 42760 18275
rect 42708 18232 42760 18241
rect 42892 18275 42944 18284
rect 42892 18241 42901 18275
rect 42901 18241 42935 18275
rect 42935 18241 42944 18275
rect 42892 18232 42944 18241
rect 43076 18275 43128 18284
rect 43076 18241 43090 18275
rect 43090 18241 43124 18275
rect 43124 18241 43128 18275
rect 43076 18232 43128 18241
rect 43352 18232 43404 18284
rect 44180 18232 44232 18284
rect 46388 18232 46440 18284
rect 48780 18275 48832 18284
rect 48780 18241 48814 18275
rect 48814 18241 48832 18275
rect 48780 18232 48832 18241
rect 49608 18232 49660 18284
rect 42156 18164 42208 18216
rect 42248 18164 42300 18216
rect 43168 18164 43220 18216
rect 48136 18164 48188 18216
rect 49608 18028 49660 18080
rect 52184 18028 52236 18080
rect 55036 18368 55088 18420
rect 57152 18411 57204 18420
rect 57152 18377 57161 18411
rect 57161 18377 57195 18411
rect 57195 18377 57204 18411
rect 57152 18368 57204 18377
rect 54576 18275 54628 18284
rect 54576 18241 54585 18275
rect 54585 18241 54619 18275
rect 54619 18241 54628 18275
rect 54576 18232 54628 18241
rect 56508 18300 56560 18352
rect 55864 18232 55916 18284
rect 54392 18096 54444 18148
rect 57612 18028 57664 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 8024 17867 8076 17876
rect 8024 17833 8033 17867
rect 8033 17833 8067 17867
rect 8067 17833 8076 17867
rect 8024 17824 8076 17833
rect 8116 17756 8168 17808
rect 9128 17824 9180 17876
rect 9680 17824 9732 17876
rect 13360 17867 13412 17876
rect 13360 17833 13369 17867
rect 13369 17833 13403 17867
rect 13403 17833 13412 17867
rect 13360 17824 13412 17833
rect 14832 17824 14884 17876
rect 15568 17824 15620 17876
rect 16672 17824 16724 17876
rect 17316 17867 17368 17876
rect 17316 17833 17325 17867
rect 17325 17833 17359 17867
rect 17359 17833 17368 17867
rect 17316 17824 17368 17833
rect 19340 17824 19392 17876
rect 19708 17824 19760 17876
rect 23388 17824 23440 17876
rect 24584 17867 24636 17876
rect 24584 17833 24593 17867
rect 24593 17833 24627 17867
rect 24627 17833 24636 17867
rect 24584 17824 24636 17833
rect 28632 17867 28684 17876
rect 9496 17756 9548 17808
rect 12992 17756 13044 17808
rect 13176 17799 13228 17808
rect 13176 17765 13185 17799
rect 13185 17765 13219 17799
rect 13219 17765 13228 17799
rect 13176 17756 13228 17765
rect 1584 17663 1636 17672
rect 1584 17629 1593 17663
rect 1593 17629 1627 17663
rect 1627 17629 1636 17663
rect 1584 17620 1636 17629
rect 1860 17595 1912 17604
rect 1860 17561 1869 17595
rect 1869 17561 1903 17595
rect 1903 17561 1912 17595
rect 1860 17552 1912 17561
rect 9220 17620 9272 17672
rect 9496 17663 9548 17672
rect 9496 17629 9505 17663
rect 9505 17629 9539 17663
rect 9539 17629 9548 17663
rect 9496 17620 9548 17629
rect 10048 17620 10100 17672
rect 13084 17620 13136 17672
rect 22652 17688 22704 17740
rect 23204 17731 23256 17740
rect 23204 17697 23213 17731
rect 23213 17697 23247 17731
rect 23247 17697 23256 17731
rect 23204 17688 23256 17697
rect 14832 17663 14884 17672
rect 14832 17629 14841 17663
rect 14841 17629 14875 17663
rect 14875 17629 14884 17663
rect 14832 17620 14884 17629
rect 9404 17595 9456 17604
rect 9404 17561 9413 17595
rect 9413 17561 9447 17595
rect 9447 17561 9456 17595
rect 9404 17552 9456 17561
rect 9588 17484 9640 17536
rect 15936 17552 15988 17604
rect 15384 17484 15436 17536
rect 15844 17484 15896 17536
rect 19524 17620 19576 17672
rect 19984 17620 20036 17672
rect 24584 17688 24636 17740
rect 25044 17688 25096 17740
rect 26056 17688 26108 17740
rect 28632 17833 28641 17867
rect 28641 17833 28675 17867
rect 28675 17833 28684 17867
rect 28632 17824 28684 17833
rect 27344 17756 27396 17808
rect 30656 17824 30708 17876
rect 30380 17756 30432 17808
rect 38844 17824 38896 17876
rect 46020 17824 46072 17876
rect 48504 17824 48556 17876
rect 16304 17552 16356 17604
rect 19708 17552 19760 17604
rect 17776 17484 17828 17536
rect 23480 17620 23532 17672
rect 24952 17663 25004 17672
rect 24952 17629 24961 17663
rect 24961 17629 24995 17663
rect 24995 17629 25004 17663
rect 24952 17620 25004 17629
rect 26240 17620 26292 17672
rect 26700 17620 26752 17672
rect 23664 17552 23716 17604
rect 27896 17620 27948 17672
rect 28080 17663 28132 17672
rect 28080 17629 28089 17663
rect 28089 17629 28123 17663
rect 28123 17629 28132 17663
rect 28080 17620 28132 17629
rect 28172 17620 28224 17672
rect 30472 17688 30524 17740
rect 27252 17552 27304 17604
rect 31208 17620 31260 17672
rect 31392 17663 31444 17672
rect 31392 17629 31401 17663
rect 31401 17629 31435 17663
rect 31435 17629 31444 17663
rect 31392 17620 31444 17629
rect 32404 17731 32456 17740
rect 32404 17697 32413 17731
rect 32413 17697 32447 17731
rect 32447 17697 32456 17731
rect 32404 17688 32456 17697
rect 33048 17688 33100 17740
rect 33784 17688 33836 17740
rect 24860 17484 24912 17536
rect 25044 17527 25096 17536
rect 25044 17493 25053 17527
rect 25053 17493 25087 17527
rect 25087 17493 25096 17527
rect 25044 17484 25096 17493
rect 25780 17484 25832 17536
rect 27620 17484 27672 17536
rect 30472 17552 30524 17604
rect 30656 17552 30708 17604
rect 29920 17484 29972 17536
rect 32128 17552 32180 17604
rect 34428 17620 34480 17672
rect 35164 17688 35216 17740
rect 39120 17688 39172 17740
rect 35256 17663 35308 17672
rect 35256 17629 35265 17663
rect 35265 17629 35299 17663
rect 35299 17629 35308 17663
rect 35256 17620 35308 17629
rect 38936 17620 38988 17672
rect 32864 17552 32916 17604
rect 33048 17595 33100 17604
rect 33048 17561 33057 17595
rect 33057 17561 33091 17595
rect 33091 17561 33100 17595
rect 33048 17552 33100 17561
rect 33876 17552 33928 17604
rect 33232 17484 33284 17536
rect 33692 17527 33744 17536
rect 33692 17493 33701 17527
rect 33701 17493 33735 17527
rect 33735 17493 33744 17527
rect 33692 17484 33744 17493
rect 34336 17484 34388 17536
rect 34520 17552 34572 17604
rect 40592 17663 40644 17672
rect 40592 17629 40626 17663
rect 40626 17629 40644 17663
rect 40592 17620 40644 17629
rect 48228 17663 48280 17672
rect 48228 17629 48237 17663
rect 48237 17629 48271 17663
rect 48271 17629 48280 17663
rect 48228 17620 48280 17629
rect 48320 17620 48372 17672
rect 55588 17824 55640 17876
rect 57060 17824 57112 17876
rect 54576 17756 54628 17808
rect 56508 17688 56560 17740
rect 39120 17527 39172 17536
rect 39120 17493 39129 17527
rect 39129 17493 39163 17527
rect 39163 17493 39172 17527
rect 39120 17484 39172 17493
rect 39672 17484 39724 17536
rect 43076 17552 43128 17604
rect 47676 17552 47728 17604
rect 49608 17552 49660 17604
rect 50620 17595 50672 17604
rect 50620 17561 50629 17595
rect 50629 17561 50663 17595
rect 50663 17561 50672 17595
rect 50620 17552 50672 17561
rect 51080 17620 51132 17672
rect 52460 17620 52512 17672
rect 54576 17620 54628 17672
rect 51724 17595 51776 17604
rect 51724 17561 51758 17595
rect 51758 17561 51776 17595
rect 51724 17552 51776 17561
rect 52368 17552 52420 17604
rect 58900 17620 58952 17672
rect 56140 17552 56192 17604
rect 41880 17484 41932 17536
rect 51540 17484 51592 17536
rect 53104 17484 53156 17536
rect 58348 17484 58400 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 13728 17323 13780 17332
rect 13728 17289 13737 17323
rect 13737 17289 13771 17323
rect 13771 17289 13780 17323
rect 13728 17280 13780 17289
rect 15384 17280 15436 17332
rect 16580 17280 16632 17332
rect 16672 17280 16724 17332
rect 21272 17280 21324 17332
rect 22652 17280 22704 17332
rect 2412 17187 2464 17196
rect 2412 17153 2421 17187
rect 2421 17153 2455 17187
rect 2455 17153 2464 17187
rect 2412 17144 2464 17153
rect 8208 17187 8260 17196
rect 8208 17153 8217 17187
rect 8217 17153 8251 17187
rect 8251 17153 8260 17187
rect 8208 17144 8260 17153
rect 12532 17187 12584 17196
rect 1768 17119 1820 17128
rect 1768 17085 1777 17119
rect 1777 17085 1811 17119
rect 1811 17085 1820 17119
rect 1768 17076 1820 17085
rect 7012 17076 7064 17128
rect 9772 17076 9824 17128
rect 12532 17153 12541 17187
rect 12541 17153 12575 17187
rect 12575 17153 12584 17187
rect 12532 17144 12584 17153
rect 16120 17144 16172 17196
rect 16396 17076 16448 17128
rect 16764 17076 16816 17128
rect 20720 17144 20772 17196
rect 21088 17187 21140 17196
rect 21088 17153 21097 17187
rect 21097 17153 21131 17187
rect 21131 17153 21140 17187
rect 21088 17144 21140 17153
rect 21272 17144 21324 17196
rect 9588 16940 9640 16992
rect 15016 16940 15068 16992
rect 20444 17008 20496 17060
rect 20996 17076 21048 17128
rect 24584 17144 24636 17196
rect 25228 17212 25280 17264
rect 25412 17255 25464 17264
rect 25412 17221 25421 17255
rect 25421 17221 25455 17255
rect 25455 17221 25464 17255
rect 25412 17212 25464 17221
rect 25872 17212 25924 17264
rect 27344 17280 27396 17332
rect 25136 17187 25188 17196
rect 25136 17153 25145 17187
rect 25145 17153 25179 17187
rect 25179 17153 25188 17187
rect 25136 17144 25188 17153
rect 25964 17144 26016 17196
rect 26424 17144 26476 17196
rect 26516 17187 26568 17196
rect 26516 17153 26525 17187
rect 26525 17153 26559 17187
rect 26559 17153 26568 17187
rect 26516 17144 26568 17153
rect 27528 17187 27580 17196
rect 27528 17153 27537 17187
rect 27537 17153 27571 17187
rect 27571 17153 27580 17187
rect 27528 17144 27580 17153
rect 31852 17280 31904 17332
rect 33692 17280 33744 17332
rect 38752 17280 38804 17332
rect 51724 17323 51776 17332
rect 51724 17289 51733 17323
rect 51733 17289 51767 17323
rect 51767 17289 51776 17323
rect 51724 17280 51776 17289
rect 52276 17280 52328 17332
rect 54668 17280 54720 17332
rect 54760 17280 54812 17332
rect 27804 17255 27856 17264
rect 27804 17221 27813 17255
rect 27813 17221 27847 17255
rect 27847 17221 27856 17255
rect 27804 17212 27856 17221
rect 27896 17187 27948 17196
rect 27896 17153 27905 17187
rect 27905 17153 27939 17187
rect 27939 17153 27948 17187
rect 27896 17144 27948 17153
rect 28356 17212 28408 17264
rect 28908 17255 28960 17264
rect 28908 17221 28917 17255
rect 28917 17221 28951 17255
rect 28951 17221 28960 17255
rect 28908 17212 28960 17221
rect 28724 17187 28776 17196
rect 28724 17153 28731 17187
rect 28731 17153 28776 17187
rect 28724 17144 28776 17153
rect 28816 17187 28868 17196
rect 28816 17153 28825 17187
rect 28825 17153 28859 17187
rect 28859 17153 28868 17187
rect 29368 17212 29420 17264
rect 29644 17212 29696 17264
rect 30748 17212 30800 17264
rect 31760 17212 31812 17264
rect 32588 17212 32640 17264
rect 28816 17144 28868 17153
rect 18144 16940 18196 16992
rect 18880 16983 18932 16992
rect 18880 16949 18889 16983
rect 18889 16949 18923 16983
rect 18923 16949 18932 16983
rect 18880 16940 18932 16949
rect 20996 16940 21048 16992
rect 23664 16940 23716 16992
rect 24124 16940 24176 16992
rect 25596 16940 25648 16992
rect 26884 16940 26936 16992
rect 28540 17008 28592 17060
rect 29092 17008 29144 17060
rect 30012 17187 30064 17196
rect 30012 17153 30021 17187
rect 30021 17153 30055 17187
rect 30055 17153 30064 17187
rect 30012 17144 30064 17153
rect 35256 17212 35308 17264
rect 35992 17212 36044 17264
rect 29276 17076 29328 17128
rect 31208 17076 31260 17128
rect 33968 17187 34020 17196
rect 33968 17153 34002 17187
rect 34002 17153 34020 17187
rect 38568 17255 38620 17264
rect 38568 17221 38577 17255
rect 38577 17221 38611 17255
rect 38611 17221 38620 17255
rect 38568 17212 38620 17221
rect 40316 17212 40368 17264
rect 40684 17212 40736 17264
rect 40960 17255 41012 17264
rect 40960 17221 40969 17255
rect 40969 17221 41003 17255
rect 41003 17221 41012 17255
rect 40960 17212 41012 17221
rect 41052 17255 41104 17264
rect 41052 17221 41061 17255
rect 41061 17221 41095 17255
rect 41095 17221 41104 17255
rect 41052 17212 41104 17221
rect 41328 17212 41380 17264
rect 52368 17212 52420 17264
rect 52460 17212 52512 17264
rect 55680 17280 55732 17332
rect 56140 17323 56192 17332
rect 56140 17289 56149 17323
rect 56149 17289 56183 17323
rect 56183 17289 56192 17323
rect 56140 17280 56192 17289
rect 57060 17280 57112 17332
rect 33968 17144 34020 17153
rect 51172 17144 51224 17196
rect 51356 17187 51408 17196
rect 51356 17153 51365 17187
rect 51365 17153 51399 17187
rect 51399 17153 51408 17187
rect 51356 17144 51408 17153
rect 51540 17187 51592 17196
rect 51540 17153 51549 17187
rect 51549 17153 51583 17187
rect 51583 17153 51592 17187
rect 51540 17144 51592 17153
rect 54300 17144 54352 17196
rect 32404 17076 32456 17128
rect 32128 17008 32180 17060
rect 32864 17076 32916 17128
rect 33140 17076 33192 17128
rect 38752 17076 38804 17128
rect 38844 17119 38896 17128
rect 38844 17085 38853 17119
rect 38853 17085 38887 17119
rect 38887 17085 38896 17119
rect 38844 17076 38896 17085
rect 43904 17076 43956 17128
rect 51448 17076 51500 17128
rect 52092 17076 52144 17128
rect 53932 17119 53984 17128
rect 53932 17085 53941 17119
rect 53941 17085 53975 17119
rect 53975 17085 53984 17119
rect 53932 17076 53984 17085
rect 38476 17008 38528 17060
rect 39304 17008 39356 17060
rect 39488 17008 39540 17060
rect 39764 17008 39816 17060
rect 48320 17008 48372 17060
rect 55772 17119 55824 17128
rect 55772 17085 55781 17119
rect 55781 17085 55815 17119
rect 55815 17085 55824 17119
rect 55772 17076 55824 17085
rect 56048 17144 56100 17196
rect 57336 17119 57388 17128
rect 57336 17085 57345 17119
rect 57345 17085 57379 17119
rect 57379 17085 57388 17119
rect 57336 17076 57388 17085
rect 35348 16940 35400 16992
rect 38200 16983 38252 16992
rect 38200 16949 38209 16983
rect 38209 16949 38243 16983
rect 38243 16949 38252 16983
rect 38200 16940 38252 16949
rect 39120 16940 39172 16992
rect 40040 16940 40092 16992
rect 44180 16940 44232 16992
rect 54116 16940 54168 16992
rect 54300 16983 54352 16992
rect 54300 16949 54309 16983
rect 54309 16949 54343 16983
rect 54343 16949 54352 16983
rect 54300 16940 54352 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 1584 16668 1636 16720
rect 7564 16532 7616 16584
rect 9128 16575 9180 16584
rect 9128 16541 9137 16575
rect 9137 16541 9171 16575
rect 9171 16541 9180 16575
rect 9128 16532 9180 16541
rect 9404 16600 9456 16652
rect 14280 16736 14332 16788
rect 16764 16668 16816 16720
rect 17132 16668 17184 16720
rect 17408 16668 17460 16720
rect 12808 16532 12860 16584
rect 13360 16575 13412 16584
rect 1860 16507 1912 16516
rect 1860 16473 1869 16507
rect 1869 16473 1903 16507
rect 1903 16473 1912 16507
rect 1860 16464 1912 16473
rect 12900 16464 12952 16516
rect 13360 16541 13369 16575
rect 13369 16541 13403 16575
rect 13403 16541 13412 16575
rect 13360 16532 13412 16541
rect 13728 16532 13780 16584
rect 14280 16532 14332 16584
rect 16580 16575 16632 16584
rect 15016 16507 15068 16516
rect 15016 16473 15050 16507
rect 15050 16473 15068 16507
rect 15016 16464 15068 16473
rect 16580 16541 16589 16575
rect 16589 16541 16623 16575
rect 16623 16541 16632 16575
rect 16580 16532 16632 16541
rect 22468 16600 22520 16652
rect 23388 16643 23440 16652
rect 23388 16609 23397 16643
rect 23397 16609 23431 16643
rect 23431 16609 23440 16643
rect 23388 16600 23440 16609
rect 23572 16600 23624 16652
rect 24768 16668 24820 16720
rect 16856 16464 16908 16516
rect 20076 16532 20128 16584
rect 22192 16532 22244 16584
rect 22836 16575 22888 16584
rect 22836 16541 22878 16575
rect 22878 16541 22888 16575
rect 22836 16532 22888 16541
rect 21088 16464 21140 16516
rect 23204 16532 23256 16584
rect 23848 16575 23900 16584
rect 23848 16541 23857 16575
rect 23857 16541 23891 16575
rect 23891 16541 23900 16575
rect 23848 16532 23900 16541
rect 24492 16532 24544 16584
rect 24860 16532 24912 16584
rect 9312 16439 9364 16448
rect 9312 16405 9321 16439
rect 9321 16405 9355 16439
rect 9355 16405 9364 16439
rect 9312 16396 9364 16405
rect 16396 16396 16448 16448
rect 16580 16396 16632 16448
rect 16948 16396 17000 16448
rect 17960 16439 18012 16448
rect 17960 16405 17969 16439
rect 17969 16405 18003 16439
rect 18003 16405 18012 16439
rect 17960 16396 18012 16405
rect 18052 16396 18104 16448
rect 22284 16396 22336 16448
rect 23388 16396 23440 16448
rect 24860 16439 24912 16448
rect 24860 16405 24869 16439
rect 24869 16405 24903 16439
rect 24903 16405 24912 16439
rect 24860 16396 24912 16405
rect 25044 16396 25096 16448
rect 25412 16396 25464 16448
rect 26332 16736 26384 16788
rect 26884 16736 26936 16788
rect 28632 16736 28684 16788
rect 31668 16668 31720 16720
rect 27068 16600 27120 16652
rect 28264 16600 28316 16652
rect 28448 16600 28500 16652
rect 30012 16600 30064 16652
rect 33140 16736 33192 16788
rect 33600 16736 33652 16788
rect 35348 16736 35400 16788
rect 26792 16532 26844 16584
rect 27896 16575 27948 16584
rect 27896 16541 27905 16575
rect 27905 16541 27939 16575
rect 27939 16541 27948 16575
rect 27896 16532 27948 16541
rect 28908 16575 28960 16584
rect 28908 16541 28917 16575
rect 28917 16541 28951 16575
rect 28951 16541 28960 16575
rect 28908 16532 28960 16541
rect 36084 16600 36136 16652
rect 36728 16643 36780 16652
rect 36728 16609 36737 16643
rect 36737 16609 36771 16643
rect 36771 16609 36780 16643
rect 36728 16600 36780 16609
rect 39672 16736 39724 16788
rect 52276 16736 52328 16788
rect 52460 16736 52512 16788
rect 38936 16668 38988 16720
rect 39488 16668 39540 16720
rect 33048 16532 33100 16584
rect 33232 16575 33284 16584
rect 33232 16541 33266 16575
rect 33266 16541 33284 16575
rect 33232 16532 33284 16541
rect 36360 16532 36412 16584
rect 38752 16600 38804 16652
rect 38200 16532 38252 16584
rect 26240 16396 26292 16448
rect 27068 16439 27120 16448
rect 27068 16405 27077 16439
rect 27077 16405 27111 16439
rect 27111 16405 27120 16439
rect 27068 16396 27120 16405
rect 30380 16464 30432 16516
rect 32220 16464 32272 16516
rect 32496 16464 32548 16516
rect 36544 16507 36596 16516
rect 36544 16473 36553 16507
rect 36553 16473 36587 16507
rect 36587 16473 36596 16507
rect 36544 16464 36596 16473
rect 28264 16396 28316 16448
rect 28724 16396 28776 16448
rect 29092 16439 29144 16448
rect 29092 16405 29101 16439
rect 29101 16405 29135 16439
rect 29135 16405 29144 16439
rect 29092 16396 29144 16405
rect 34336 16439 34388 16448
rect 34336 16405 34345 16439
rect 34345 16405 34379 16439
rect 34379 16405 34388 16439
rect 34336 16396 34388 16405
rect 36452 16396 36504 16448
rect 36728 16396 36780 16448
rect 38384 16396 38436 16448
rect 38660 16396 38712 16448
rect 40868 16532 40920 16584
rect 41052 16575 41104 16584
rect 41052 16541 41061 16575
rect 41061 16541 41095 16575
rect 41095 16541 41104 16575
rect 42892 16668 42944 16720
rect 41052 16532 41104 16541
rect 41236 16464 41288 16516
rect 41328 16464 41380 16516
rect 41420 16464 41472 16516
rect 42064 16575 42116 16584
rect 42064 16541 42073 16575
rect 42073 16541 42107 16575
rect 42107 16541 42116 16575
rect 42708 16600 42760 16652
rect 44732 16600 44784 16652
rect 45192 16643 45244 16652
rect 45192 16609 45201 16643
rect 45201 16609 45235 16643
rect 45235 16609 45244 16643
rect 45192 16600 45244 16609
rect 50620 16600 50672 16652
rect 50988 16600 51040 16652
rect 56508 16736 56560 16788
rect 54668 16668 54720 16720
rect 58532 16668 58584 16720
rect 42064 16532 42116 16541
rect 47124 16532 47176 16584
rect 51356 16575 51408 16584
rect 51356 16541 51365 16575
rect 51365 16541 51399 16575
rect 51399 16541 51408 16575
rect 51356 16532 51408 16541
rect 51540 16575 51592 16584
rect 51540 16541 51549 16575
rect 51549 16541 51583 16575
rect 51583 16541 51592 16575
rect 51540 16532 51592 16541
rect 43168 16464 43220 16516
rect 46388 16464 46440 16516
rect 47584 16464 47636 16516
rect 40868 16396 40920 16448
rect 46572 16439 46624 16448
rect 46572 16405 46581 16439
rect 46581 16405 46615 16439
rect 46615 16405 46624 16439
rect 46572 16396 46624 16405
rect 51724 16439 51776 16448
rect 51724 16405 51733 16439
rect 51733 16405 51767 16439
rect 51767 16405 51776 16439
rect 51724 16396 51776 16405
rect 53104 16575 53156 16584
rect 53104 16541 53113 16575
rect 53113 16541 53147 16575
rect 53147 16541 53156 16575
rect 53104 16532 53156 16541
rect 54300 16532 54352 16584
rect 57980 16575 58032 16584
rect 57980 16541 57989 16575
rect 57989 16541 58023 16575
rect 58023 16541 58032 16575
rect 57980 16532 58032 16541
rect 54576 16464 54628 16516
rect 57060 16507 57112 16516
rect 55220 16396 55272 16448
rect 56048 16396 56100 16448
rect 57060 16473 57069 16507
rect 57069 16473 57103 16507
rect 57103 16473 57112 16507
rect 57060 16464 57112 16473
rect 56968 16396 57020 16448
rect 57152 16439 57204 16448
rect 57152 16405 57161 16439
rect 57161 16405 57195 16439
rect 57195 16405 57204 16439
rect 57152 16396 57204 16405
rect 58072 16439 58124 16448
rect 58072 16405 58081 16439
rect 58081 16405 58115 16439
rect 58115 16405 58124 16439
rect 58072 16396 58124 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 13636 16192 13688 16244
rect 16672 16192 16724 16244
rect 19432 16192 19484 16244
rect 20444 16192 20496 16244
rect 7564 16124 7616 16176
rect 13084 16124 13136 16176
rect 10140 16099 10192 16108
rect 10140 16065 10149 16099
rect 10149 16065 10183 16099
rect 10183 16065 10192 16099
rect 10140 16056 10192 16065
rect 11888 16099 11940 16108
rect 11888 16065 11897 16099
rect 11897 16065 11931 16099
rect 11931 16065 11940 16099
rect 11888 16056 11940 16065
rect 14280 16124 14332 16176
rect 13452 16099 13504 16108
rect 13452 16065 13486 16099
rect 13486 16065 13504 16099
rect 13452 16056 13504 16065
rect 13728 16056 13780 16108
rect 15384 16099 15436 16108
rect 15384 16065 15393 16099
rect 15393 16065 15427 16099
rect 15427 16065 15436 16099
rect 15384 16056 15436 16065
rect 19340 16124 19392 16176
rect 21824 16192 21876 16244
rect 16120 16099 16172 16108
rect 16120 16065 16129 16099
rect 16129 16065 16163 16099
rect 16163 16065 16172 16099
rect 16120 16056 16172 16065
rect 16304 16099 16356 16108
rect 16304 16065 16313 16099
rect 16313 16065 16347 16099
rect 16347 16065 16356 16099
rect 16304 16056 16356 16065
rect 17684 16099 17736 16108
rect 17684 16065 17693 16099
rect 17693 16065 17727 16099
rect 17727 16065 17736 16099
rect 17684 16056 17736 16065
rect 19248 16056 19300 16108
rect 1768 16031 1820 16040
rect 1768 15997 1777 16031
rect 1777 15997 1811 16031
rect 1811 15997 1820 16031
rect 1768 15988 1820 15997
rect 2412 16031 2464 16040
rect 2412 15997 2421 16031
rect 2421 15997 2455 16031
rect 2455 15997 2464 16031
rect 2412 15988 2464 15997
rect 10048 15988 10100 16040
rect 12624 15988 12676 16040
rect 15568 16031 15620 16040
rect 15568 15997 15577 16031
rect 15577 15997 15611 16031
rect 15611 15997 15620 16031
rect 15568 15988 15620 15997
rect 21180 16056 21232 16108
rect 21456 16099 21508 16108
rect 21456 16065 21465 16099
rect 21465 16065 21499 16099
rect 21499 16065 21508 16099
rect 21456 16056 21508 16065
rect 22836 16124 22888 16176
rect 23572 16124 23624 16176
rect 23388 16056 23440 16108
rect 24124 16192 24176 16244
rect 27068 16192 27120 16244
rect 28908 16192 28960 16244
rect 30380 16192 30432 16244
rect 37188 16192 37240 16244
rect 24216 16124 24268 16176
rect 26792 16124 26844 16176
rect 27896 16124 27948 16176
rect 28264 16056 28316 16108
rect 29276 16124 29328 16176
rect 29460 16124 29512 16176
rect 30472 16167 30524 16176
rect 30472 16133 30481 16167
rect 30481 16133 30515 16167
rect 30515 16133 30524 16167
rect 30472 16124 30524 16133
rect 39488 16192 39540 16244
rect 41052 16192 41104 16244
rect 42064 16192 42116 16244
rect 43168 16235 43220 16244
rect 38752 16124 38804 16176
rect 38844 16124 38896 16176
rect 40132 16167 40184 16176
rect 40132 16133 40141 16167
rect 40141 16133 40175 16167
rect 40175 16133 40184 16167
rect 40132 16124 40184 16133
rect 29736 16056 29788 16108
rect 30380 16056 30432 16108
rect 32404 16099 32456 16108
rect 32404 16065 32413 16099
rect 32413 16065 32447 16099
rect 32447 16065 32456 16099
rect 32404 16056 32456 16065
rect 32588 16099 32640 16108
rect 32588 16065 32597 16099
rect 32597 16065 32631 16099
rect 32631 16065 32640 16099
rect 32588 16056 32640 16065
rect 32680 16099 32732 16108
rect 32680 16065 32689 16099
rect 32689 16065 32723 16099
rect 32723 16065 32732 16099
rect 32680 16056 32732 16065
rect 19432 15988 19484 16040
rect 21824 15988 21876 16040
rect 22008 16031 22060 16040
rect 22008 15997 22017 16031
rect 22017 15997 22051 16031
rect 22051 15997 22060 16031
rect 22008 15988 22060 15997
rect 24860 15988 24912 16040
rect 27712 15988 27764 16040
rect 27988 15988 28040 16040
rect 29552 15988 29604 16040
rect 31300 15988 31352 16040
rect 33048 16056 33100 16108
rect 39764 16056 39816 16108
rect 37004 15988 37056 16040
rect 38844 15988 38896 16040
rect 40592 16056 40644 16108
rect 41696 16056 41748 16108
rect 42156 16124 42208 16176
rect 42892 16167 42944 16176
rect 42892 16133 42901 16167
rect 42901 16133 42935 16167
rect 42935 16133 42944 16167
rect 42892 16124 42944 16133
rect 43168 16201 43177 16235
rect 43177 16201 43211 16235
rect 43211 16201 43220 16235
rect 43168 16192 43220 16201
rect 45376 16192 45428 16244
rect 46388 16235 46440 16244
rect 46388 16201 46397 16235
rect 46397 16201 46431 16235
rect 46431 16201 46440 16235
rect 46388 16192 46440 16201
rect 46572 16192 46624 16244
rect 53748 16192 53800 16244
rect 54116 16235 54168 16244
rect 54116 16201 54125 16235
rect 54125 16201 54159 16235
rect 54159 16201 54168 16235
rect 54116 16192 54168 16201
rect 54760 16235 54812 16244
rect 54760 16201 54769 16235
rect 54769 16201 54803 16235
rect 54803 16201 54812 16235
rect 54760 16192 54812 16201
rect 44180 16099 44232 16108
rect 41604 16031 41656 16040
rect 41604 15997 41613 16031
rect 41613 15997 41647 16031
rect 41647 15997 41656 16031
rect 41604 15988 41656 15997
rect 42524 15988 42576 16040
rect 9864 15852 9916 15904
rect 12256 15895 12308 15904
rect 12256 15861 12265 15895
rect 12265 15861 12299 15895
rect 12299 15861 12308 15895
rect 12256 15852 12308 15861
rect 13360 15852 13412 15904
rect 14924 15852 14976 15904
rect 16856 15920 16908 15972
rect 20904 15920 20956 15972
rect 21088 15920 21140 15972
rect 17868 15852 17920 15904
rect 19616 15852 19668 15904
rect 20076 15852 20128 15904
rect 23480 15920 23532 15972
rect 24032 15920 24084 15972
rect 29460 15920 29512 15972
rect 42064 15920 42116 15972
rect 23572 15852 23624 15904
rect 27712 15852 27764 15904
rect 30012 15852 30064 15904
rect 31024 15852 31076 15904
rect 35992 15852 36044 15904
rect 37188 15852 37240 15904
rect 40960 15895 41012 15904
rect 40960 15861 40969 15895
rect 40969 15861 41003 15895
rect 41003 15861 41012 15895
rect 40960 15852 41012 15861
rect 42892 15988 42944 16040
rect 44180 16065 44189 16099
rect 44189 16065 44223 16099
rect 44223 16065 44232 16099
rect 44180 16056 44232 16065
rect 46756 16099 46808 16108
rect 46756 16065 46765 16099
rect 46765 16065 46799 16099
rect 46799 16065 46808 16099
rect 46756 16056 46808 16065
rect 43260 15988 43312 16040
rect 46572 15988 46624 16040
rect 48228 16031 48280 16040
rect 48228 15997 48237 16031
rect 48237 15997 48271 16031
rect 48271 15997 48280 16031
rect 48228 15988 48280 15997
rect 51080 16056 51132 16108
rect 51724 16124 51776 16176
rect 55220 16124 55272 16176
rect 53932 16099 53984 16108
rect 53932 16065 53941 16099
rect 53941 16065 53975 16099
rect 53975 16065 53984 16099
rect 53932 16056 53984 16065
rect 54392 16056 54444 16108
rect 54576 16099 54628 16108
rect 54576 16065 54585 16099
rect 54585 16065 54619 16099
rect 54619 16065 54628 16099
rect 54576 16056 54628 16065
rect 48136 15920 48188 15972
rect 54760 15988 54812 16040
rect 47216 15852 47268 15904
rect 47768 15895 47820 15904
rect 47768 15861 47777 15895
rect 47777 15861 47811 15895
rect 47811 15861 47820 15895
rect 47768 15852 47820 15861
rect 51172 15852 51224 15904
rect 52368 15895 52420 15904
rect 52368 15861 52377 15895
rect 52377 15861 52411 15895
rect 52411 15861 52420 15895
rect 52368 15852 52420 15861
rect 53748 15852 53800 15904
rect 58624 15852 58676 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 13084 15648 13136 15700
rect 13360 15555 13412 15564
rect 13360 15521 13369 15555
rect 13369 15521 13403 15555
rect 13403 15521 13412 15555
rect 13360 15512 13412 15521
rect 24860 15648 24912 15700
rect 29460 15648 29512 15700
rect 29736 15691 29788 15700
rect 29736 15657 29745 15691
rect 29745 15657 29779 15691
rect 29779 15657 29788 15691
rect 29736 15648 29788 15657
rect 16304 15580 16356 15632
rect 9864 15487 9916 15496
rect 9864 15453 9873 15487
rect 9873 15453 9907 15487
rect 9907 15453 9916 15487
rect 9864 15444 9916 15453
rect 11612 15444 11664 15496
rect 13728 15512 13780 15564
rect 14280 15555 14332 15564
rect 14280 15521 14289 15555
rect 14289 15521 14323 15555
rect 14323 15521 14332 15555
rect 14280 15512 14332 15521
rect 14648 15512 14700 15564
rect 15568 15512 15620 15564
rect 18052 15512 18104 15564
rect 20260 15580 20312 15632
rect 21456 15580 21508 15632
rect 23480 15580 23532 15632
rect 23572 15512 23624 15564
rect 12716 15376 12768 15428
rect 15200 15444 15252 15496
rect 16672 15444 16724 15496
rect 19248 15376 19300 15428
rect 19616 15487 19668 15496
rect 19616 15453 19625 15487
rect 19625 15453 19659 15487
rect 19659 15453 19668 15487
rect 19616 15444 19668 15453
rect 20168 15444 20220 15496
rect 21088 15487 21140 15496
rect 21088 15453 21097 15487
rect 21097 15453 21131 15487
rect 21131 15453 21140 15487
rect 21088 15444 21140 15453
rect 24492 15444 24544 15496
rect 23204 15376 23256 15428
rect 24952 15487 25004 15496
rect 24952 15453 24966 15487
rect 24966 15453 25000 15487
rect 25000 15453 25004 15487
rect 24952 15444 25004 15453
rect 24768 15419 24820 15428
rect 24768 15385 24777 15419
rect 24777 15385 24811 15419
rect 24811 15385 24820 15419
rect 24768 15376 24820 15385
rect 10232 15308 10284 15360
rect 11888 15308 11940 15360
rect 17224 15308 17276 15360
rect 18420 15308 18472 15360
rect 19156 15308 19208 15360
rect 20076 15308 20128 15360
rect 22652 15308 22704 15360
rect 23388 15308 23440 15360
rect 23480 15308 23532 15360
rect 25136 15308 25188 15360
rect 28448 15580 28500 15632
rect 31668 15648 31720 15700
rect 41328 15648 41380 15700
rect 41696 15691 41748 15700
rect 41696 15657 41705 15691
rect 41705 15657 41739 15691
rect 41739 15657 41748 15691
rect 41696 15648 41748 15657
rect 42524 15648 42576 15700
rect 47400 15648 47452 15700
rect 51540 15691 51592 15700
rect 51540 15657 51549 15691
rect 51549 15657 51583 15691
rect 51583 15657 51592 15691
rect 51540 15648 51592 15657
rect 26332 15512 26384 15564
rect 27344 15555 27396 15564
rect 27344 15521 27353 15555
rect 27353 15521 27387 15555
rect 27387 15521 27396 15555
rect 27344 15512 27396 15521
rect 28724 15512 28776 15564
rect 28908 15512 28960 15564
rect 25320 15376 25372 15428
rect 25964 15419 26016 15428
rect 25964 15385 25973 15419
rect 25973 15385 26007 15419
rect 26007 15385 26016 15419
rect 25964 15376 26016 15385
rect 31668 15444 31720 15496
rect 32128 15487 32180 15496
rect 32128 15453 32137 15487
rect 32137 15453 32171 15487
rect 32171 15453 32180 15487
rect 32128 15444 32180 15453
rect 46756 15580 46808 15632
rect 58808 15580 58860 15632
rect 41420 15512 41472 15564
rect 34152 15444 34204 15496
rect 36360 15487 36412 15496
rect 36360 15453 36369 15487
rect 36369 15453 36403 15487
rect 36403 15453 36412 15487
rect 36360 15444 36412 15453
rect 36452 15444 36504 15496
rect 41052 15487 41104 15496
rect 41052 15453 41061 15487
rect 41061 15453 41095 15487
rect 41095 15453 41104 15487
rect 41052 15444 41104 15453
rect 29092 15376 29144 15428
rect 29276 15376 29328 15428
rect 29736 15376 29788 15428
rect 30012 15376 30064 15428
rect 27528 15308 27580 15360
rect 28264 15308 28316 15360
rect 31116 15376 31168 15428
rect 30472 15308 30524 15360
rect 34336 15376 34388 15428
rect 40132 15376 40184 15428
rect 41236 15444 41288 15496
rect 41788 15376 41840 15428
rect 36728 15308 36780 15360
rect 40592 15308 40644 15360
rect 42432 15444 42484 15496
rect 44180 15444 44232 15496
rect 51172 15487 51224 15496
rect 51172 15453 51181 15487
rect 51181 15453 51215 15487
rect 51215 15453 51224 15487
rect 51172 15444 51224 15453
rect 53932 15512 53984 15564
rect 52368 15444 52420 15496
rect 58164 15419 58216 15428
rect 58164 15385 58173 15419
rect 58173 15385 58207 15419
rect 58207 15385 58216 15419
rect 58164 15376 58216 15385
rect 48136 15351 48188 15360
rect 48136 15317 48145 15351
rect 48145 15317 48179 15351
rect 48179 15317 48188 15351
rect 48136 15308 48188 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 12900 15104 12952 15156
rect 14556 15036 14608 15088
rect 14740 15036 14792 15088
rect 15844 15036 15896 15088
rect 16396 15036 16448 15088
rect 9772 14968 9824 15020
rect 12256 15011 12308 15020
rect 12256 14977 12265 15011
rect 12265 14977 12299 15011
rect 12299 14977 12308 15011
rect 12256 14968 12308 14977
rect 12624 14968 12676 15020
rect 16028 15011 16080 15020
rect 16028 14977 16037 15011
rect 16037 14977 16071 15011
rect 16071 14977 16080 15011
rect 16028 14968 16080 14977
rect 1768 14943 1820 14952
rect 1768 14909 1777 14943
rect 1777 14909 1811 14943
rect 1811 14909 1820 14943
rect 1768 14900 1820 14909
rect 15936 14943 15988 14952
rect 15936 14909 15945 14943
rect 15945 14909 15979 14943
rect 15979 14909 15988 14943
rect 16672 14968 16724 15020
rect 16856 15011 16908 15020
rect 16856 14977 16865 15011
rect 16865 14977 16899 15011
rect 16899 14977 16908 15011
rect 16856 14968 16908 14977
rect 17960 15036 18012 15088
rect 18144 15104 18196 15156
rect 22008 15104 22060 15156
rect 18328 15036 18380 15088
rect 20076 15036 20128 15088
rect 25504 15104 25556 15156
rect 26056 15104 26108 15156
rect 26332 15036 26384 15088
rect 27528 15036 27580 15088
rect 28264 15104 28316 15156
rect 28908 15104 28960 15156
rect 29828 15104 29880 15156
rect 15936 14900 15988 14909
rect 16764 14900 16816 14952
rect 24308 14968 24360 15020
rect 24768 15011 24820 15020
rect 24768 14977 24777 15011
rect 24777 14977 24811 15011
rect 24811 14977 24820 15011
rect 24768 14968 24820 14977
rect 27620 14968 27672 15020
rect 27896 15011 27948 15020
rect 27896 14977 27905 15011
rect 27905 14977 27939 15011
rect 27939 14977 27948 15011
rect 27896 14968 27948 14977
rect 29276 15036 29328 15088
rect 30472 15104 30524 15156
rect 32588 15104 32640 15156
rect 32680 15104 32732 15156
rect 28632 14968 28684 15020
rect 29828 14968 29880 15020
rect 19248 14900 19300 14952
rect 25872 14900 25924 14952
rect 27712 14900 27764 14952
rect 27988 14900 28040 14952
rect 30104 14968 30156 15020
rect 30012 14900 30064 14952
rect 31944 15036 31996 15088
rect 32036 14968 32088 15020
rect 36360 15036 36412 15088
rect 38936 15104 38988 15156
rect 57704 15036 57756 15088
rect 34704 15011 34756 15020
rect 34704 14977 34738 15011
rect 34738 14977 34756 15011
rect 34704 14968 34756 14977
rect 40316 14968 40368 15020
rect 43536 14968 43588 15020
rect 31760 14900 31812 14952
rect 33232 14900 33284 14952
rect 38752 14900 38804 14952
rect 41144 14900 41196 14952
rect 43168 14900 43220 14952
rect 44364 14900 44416 14952
rect 54852 14900 54904 14952
rect 1584 14832 1636 14884
rect 15660 14832 15712 14884
rect 19432 14832 19484 14884
rect 31024 14832 31076 14884
rect 33508 14832 33560 14884
rect 9680 14764 9732 14816
rect 15936 14764 15988 14816
rect 18420 14764 18472 14816
rect 19524 14764 19576 14816
rect 20628 14764 20680 14816
rect 24032 14764 24084 14816
rect 24952 14764 25004 14816
rect 25412 14764 25464 14816
rect 25964 14764 26016 14816
rect 26332 14764 26384 14816
rect 28908 14764 28960 14816
rect 29092 14764 29144 14816
rect 29644 14764 29696 14816
rect 32588 14764 32640 14816
rect 34336 14764 34388 14816
rect 35900 14764 35952 14816
rect 38476 14807 38528 14816
rect 38476 14773 38485 14807
rect 38485 14773 38519 14807
rect 38519 14773 38528 14807
rect 38476 14764 38528 14773
rect 38568 14764 38620 14816
rect 39488 14832 39540 14884
rect 48320 14832 48372 14884
rect 41052 14764 41104 14816
rect 41604 14764 41656 14816
rect 52460 14764 52512 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 14556 14560 14608 14612
rect 19432 14560 19484 14612
rect 27620 14603 27672 14612
rect 19524 14492 19576 14544
rect 20812 14492 20864 14544
rect 24400 14492 24452 14544
rect 2412 14467 2464 14476
rect 2412 14433 2421 14467
rect 2421 14433 2455 14467
rect 2455 14433 2464 14467
rect 2412 14424 2464 14433
rect 8300 14424 8352 14476
rect 9312 14467 9364 14476
rect 9312 14433 9321 14467
rect 9321 14433 9355 14467
rect 9355 14433 9364 14467
rect 9312 14424 9364 14433
rect 10232 14424 10284 14476
rect 14280 14467 14332 14476
rect 14280 14433 14289 14467
rect 14289 14433 14323 14467
rect 14323 14433 14332 14467
rect 14280 14424 14332 14433
rect 15660 14424 15712 14476
rect 19248 14424 19300 14476
rect 11152 14356 11204 14408
rect 15384 14356 15436 14408
rect 18052 14356 18104 14408
rect 19800 14356 19852 14408
rect 21824 14424 21876 14476
rect 22008 14424 22060 14476
rect 21640 14399 21692 14408
rect 21640 14365 21649 14399
rect 21649 14365 21683 14399
rect 21683 14365 21692 14399
rect 27620 14569 27629 14603
rect 27629 14569 27663 14603
rect 27663 14569 27672 14603
rect 27620 14560 27672 14569
rect 27712 14560 27764 14612
rect 29276 14560 29328 14612
rect 31116 14603 31168 14612
rect 31116 14569 31125 14603
rect 31125 14569 31159 14603
rect 31159 14569 31168 14603
rect 31116 14560 31168 14569
rect 32036 14560 32088 14612
rect 35256 14560 35308 14612
rect 24860 14424 24912 14476
rect 26148 14424 26200 14476
rect 21640 14356 21692 14365
rect 1860 14331 1912 14340
rect 1860 14297 1869 14331
rect 1869 14297 1903 14331
rect 1903 14297 1912 14331
rect 1860 14288 1912 14297
rect 12440 14288 12492 14340
rect 16764 14288 16816 14340
rect 17592 14288 17644 14340
rect 19616 14288 19668 14340
rect 11980 14220 12032 14272
rect 15660 14263 15712 14272
rect 15660 14229 15669 14263
rect 15669 14229 15703 14263
rect 15703 14229 15712 14263
rect 15660 14220 15712 14229
rect 17776 14263 17828 14272
rect 17776 14229 17785 14263
rect 17785 14229 17819 14263
rect 17819 14229 17828 14263
rect 17776 14220 17828 14229
rect 21456 14288 21508 14340
rect 23848 14288 23900 14340
rect 24308 14288 24360 14340
rect 25412 14331 25464 14340
rect 25412 14297 25421 14331
rect 25421 14297 25455 14331
rect 25455 14297 25464 14331
rect 25412 14288 25464 14297
rect 20904 14220 20956 14272
rect 21088 14263 21140 14272
rect 21088 14229 21097 14263
rect 21097 14229 21131 14263
rect 21131 14229 21140 14263
rect 21088 14220 21140 14229
rect 22928 14220 22980 14272
rect 25872 14356 25924 14408
rect 26424 14424 26476 14476
rect 27160 14424 27212 14476
rect 29644 14492 29696 14544
rect 30748 14492 30800 14544
rect 26608 14399 26660 14408
rect 26608 14365 26617 14399
rect 26617 14365 26651 14399
rect 26651 14365 26660 14399
rect 27252 14399 27304 14408
rect 26608 14356 26660 14365
rect 27252 14365 27261 14399
rect 27261 14365 27295 14399
rect 27295 14365 27304 14399
rect 27252 14356 27304 14365
rect 29092 14424 29144 14476
rect 29276 14356 29328 14408
rect 29736 14399 29788 14408
rect 29736 14365 29745 14399
rect 29745 14365 29779 14399
rect 29779 14365 29788 14399
rect 29736 14356 29788 14365
rect 32680 14399 32732 14408
rect 26332 14288 26384 14340
rect 27988 14288 28040 14340
rect 30196 14288 30248 14340
rect 32680 14365 32689 14399
rect 32689 14365 32723 14399
rect 32723 14365 32732 14399
rect 32680 14356 32732 14365
rect 33416 14424 33468 14476
rect 33048 14356 33100 14408
rect 35992 14492 36044 14544
rect 39488 14560 39540 14612
rect 40224 14560 40276 14612
rect 40316 14560 40368 14612
rect 44364 14560 44416 14612
rect 44548 14603 44600 14612
rect 44548 14569 44557 14603
rect 44557 14569 44591 14603
rect 44591 14569 44600 14603
rect 44548 14560 44600 14569
rect 48228 14560 48280 14612
rect 48320 14560 48372 14612
rect 56600 14560 56652 14612
rect 56784 14492 56836 14544
rect 34612 14424 34664 14476
rect 35072 14424 35124 14476
rect 35164 14424 35216 14476
rect 35624 14424 35676 14476
rect 37372 14399 37424 14408
rect 25688 14220 25740 14272
rect 27160 14220 27212 14272
rect 31668 14220 31720 14272
rect 31760 14220 31812 14272
rect 33508 14220 33560 14272
rect 33600 14220 33652 14272
rect 37372 14365 37381 14399
rect 37381 14365 37415 14399
rect 37415 14365 37424 14399
rect 37372 14356 37424 14365
rect 41052 14424 41104 14476
rect 39948 14356 40000 14408
rect 43076 14356 43128 14408
rect 43260 14399 43312 14408
rect 43260 14365 43269 14399
rect 43269 14365 43303 14399
rect 43303 14365 43312 14399
rect 43260 14356 43312 14365
rect 34888 14263 34940 14272
rect 34888 14229 34897 14263
rect 34897 14229 34931 14263
rect 34931 14229 34940 14263
rect 34888 14220 34940 14229
rect 35072 14220 35124 14272
rect 35900 14220 35952 14272
rect 39120 14288 39172 14340
rect 41788 14220 41840 14272
rect 48136 14356 48188 14408
rect 57980 14399 58032 14408
rect 57980 14365 57989 14399
rect 57989 14365 58023 14399
rect 58023 14365 58032 14399
rect 57980 14356 58032 14365
rect 47768 14288 47820 14340
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 10048 14059 10100 14068
rect 10048 14025 10057 14059
rect 10057 14025 10091 14059
rect 10091 14025 10100 14059
rect 10048 14016 10100 14025
rect 1584 13923 1636 13932
rect 1584 13889 1593 13923
rect 1593 13889 1627 13923
rect 1627 13889 1636 13923
rect 1584 13880 1636 13889
rect 8852 13923 8904 13932
rect 8852 13889 8861 13923
rect 8861 13889 8895 13923
rect 8895 13889 8904 13923
rect 8852 13880 8904 13889
rect 9312 13880 9364 13932
rect 14280 13948 14332 14000
rect 17776 13948 17828 14000
rect 21088 14016 21140 14068
rect 24400 14016 24452 14068
rect 26424 14016 26476 14068
rect 28080 14016 28132 14068
rect 29276 14059 29328 14068
rect 29276 14025 29285 14059
rect 29285 14025 29319 14059
rect 29319 14025 29328 14059
rect 29276 14016 29328 14025
rect 21640 13948 21692 14000
rect 11980 13923 12032 13932
rect 11980 13889 12014 13923
rect 12014 13889 12032 13923
rect 11980 13880 12032 13889
rect 13728 13923 13780 13932
rect 13728 13889 13737 13923
rect 13737 13889 13771 13923
rect 13771 13889 13780 13923
rect 13728 13880 13780 13889
rect 16856 13923 16908 13932
rect 16856 13889 16865 13923
rect 16865 13889 16899 13923
rect 16899 13889 16908 13923
rect 16856 13880 16908 13889
rect 20720 13880 20772 13932
rect 21456 13923 21508 13932
rect 21456 13889 21465 13923
rect 21465 13889 21499 13923
rect 21499 13889 21508 13923
rect 21456 13880 21508 13889
rect 21824 13923 21876 13932
rect 21824 13889 21833 13923
rect 21833 13889 21867 13923
rect 21867 13889 21876 13923
rect 21824 13880 21876 13889
rect 22376 13880 22428 13932
rect 1768 13855 1820 13864
rect 1768 13821 1777 13855
rect 1777 13821 1811 13855
rect 1811 13821 1820 13855
rect 1768 13812 1820 13821
rect 15200 13855 15252 13864
rect 15200 13821 15209 13855
rect 15209 13821 15243 13855
rect 15243 13821 15252 13855
rect 15200 13812 15252 13821
rect 18236 13812 18288 13864
rect 20812 13812 20864 13864
rect 1584 13676 1636 13728
rect 21824 13744 21876 13796
rect 17960 13676 18012 13728
rect 19432 13676 19484 13728
rect 22192 13676 22244 13728
rect 23020 13948 23072 14000
rect 23940 13948 23992 14000
rect 31760 14016 31812 14068
rect 32128 14016 32180 14068
rect 33048 14016 33100 14068
rect 34520 14016 34572 14068
rect 35624 14016 35676 14068
rect 37372 14016 37424 14068
rect 23572 13923 23624 13932
rect 23572 13889 23581 13923
rect 23581 13889 23615 13923
rect 23615 13889 23624 13923
rect 23572 13880 23624 13889
rect 23020 13812 23072 13864
rect 24952 13880 25004 13932
rect 23204 13787 23256 13796
rect 23204 13753 23213 13787
rect 23213 13753 23247 13787
rect 23247 13753 23256 13787
rect 23204 13744 23256 13753
rect 24400 13812 24452 13864
rect 24860 13812 24912 13864
rect 25688 13923 25740 13932
rect 25688 13889 25697 13923
rect 25697 13889 25731 13923
rect 25731 13889 25740 13923
rect 25688 13880 25740 13889
rect 25964 13744 26016 13796
rect 26516 13880 26568 13932
rect 27528 13923 27580 13932
rect 27528 13889 27537 13923
rect 27537 13889 27571 13923
rect 27571 13889 27580 13923
rect 27528 13880 27580 13889
rect 29644 13923 29696 13932
rect 29644 13889 29653 13923
rect 29653 13889 29687 13923
rect 29687 13889 29696 13923
rect 29644 13880 29696 13889
rect 32036 13948 32088 14000
rect 33416 13948 33468 14000
rect 38936 14016 38988 14068
rect 39120 14059 39172 14068
rect 39120 14025 39129 14059
rect 39129 14025 39163 14059
rect 39163 14025 39172 14059
rect 39120 14016 39172 14025
rect 42800 14016 42852 14068
rect 44088 14016 44140 14068
rect 31300 13880 31352 13932
rect 31484 13923 31536 13932
rect 31484 13889 31493 13923
rect 31493 13889 31527 13923
rect 31527 13889 31536 13923
rect 31484 13880 31536 13889
rect 31852 13880 31904 13932
rect 31944 13880 31996 13932
rect 32680 13880 32732 13932
rect 26424 13855 26476 13864
rect 26424 13821 26433 13855
rect 26433 13821 26467 13855
rect 26467 13821 26476 13855
rect 26424 13812 26476 13821
rect 27252 13812 27304 13864
rect 29368 13812 29420 13864
rect 28632 13744 28684 13796
rect 29000 13744 29052 13796
rect 30012 13812 30064 13864
rect 32404 13812 32456 13864
rect 35716 13880 35768 13932
rect 36820 13880 36872 13932
rect 37372 13880 37424 13932
rect 39488 13948 39540 14000
rect 38476 13880 38528 13932
rect 41604 13948 41656 14000
rect 41512 13923 41564 13932
rect 41512 13889 41521 13923
rect 41521 13889 41555 13923
rect 41555 13889 41564 13923
rect 41512 13880 41564 13889
rect 41696 13923 41748 13932
rect 41696 13889 41705 13923
rect 41705 13889 41739 13923
rect 41739 13889 41748 13923
rect 41696 13880 41748 13889
rect 42800 13880 42852 13932
rect 43076 13923 43128 13932
rect 43076 13889 43085 13923
rect 43085 13889 43119 13923
rect 43119 13889 43128 13923
rect 43076 13880 43128 13889
rect 34612 13812 34664 13864
rect 35164 13855 35216 13864
rect 35164 13821 35173 13855
rect 35173 13821 35207 13855
rect 35207 13821 35216 13855
rect 35164 13812 35216 13821
rect 38660 13812 38712 13864
rect 43352 13855 43404 13864
rect 43352 13821 43361 13855
rect 43361 13821 43395 13855
rect 43395 13821 43404 13855
rect 43352 13812 43404 13821
rect 57244 13812 57296 13864
rect 30656 13744 30708 13796
rect 26240 13676 26292 13728
rect 34520 13719 34572 13728
rect 34520 13685 34529 13719
rect 34529 13685 34563 13719
rect 34563 13685 34572 13719
rect 34520 13676 34572 13685
rect 34704 13676 34756 13728
rect 42064 13719 42116 13728
rect 42064 13685 42073 13719
rect 42073 13685 42107 13719
rect 42107 13685 42116 13719
rect 42064 13676 42116 13685
rect 49056 13744 49108 13796
rect 55220 13744 55272 13796
rect 43536 13676 43588 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 16028 13472 16080 13524
rect 17316 13472 17368 13524
rect 17868 13472 17920 13524
rect 18880 13472 18932 13524
rect 19340 13472 19392 13524
rect 19800 13472 19852 13524
rect 18420 13404 18472 13456
rect 20720 13472 20772 13524
rect 23940 13472 23992 13524
rect 26424 13472 26476 13524
rect 27344 13515 27396 13524
rect 27344 13481 27353 13515
rect 27353 13481 27387 13515
rect 27387 13481 27396 13515
rect 27344 13472 27396 13481
rect 27896 13472 27948 13524
rect 31576 13472 31628 13524
rect 38200 13472 38252 13524
rect 38292 13472 38344 13524
rect 9312 13379 9364 13388
rect 9312 13345 9321 13379
rect 9321 13345 9355 13379
rect 9355 13345 9364 13379
rect 9312 13336 9364 13345
rect 9680 13336 9732 13388
rect 14280 13379 14332 13388
rect 14280 13345 14289 13379
rect 14289 13345 14323 13379
rect 14323 13345 14332 13379
rect 14280 13336 14332 13345
rect 16304 13336 16356 13388
rect 1584 13311 1636 13320
rect 1584 13277 1593 13311
rect 1593 13277 1627 13311
rect 1627 13277 1636 13311
rect 1584 13268 1636 13277
rect 11428 13311 11480 13320
rect 11428 13277 11437 13311
rect 11437 13277 11471 13311
rect 11471 13277 11480 13311
rect 11428 13268 11480 13277
rect 13544 13268 13596 13320
rect 16764 13268 16816 13320
rect 17224 13336 17276 13388
rect 17868 13336 17920 13388
rect 18144 13379 18196 13388
rect 18144 13345 18153 13379
rect 18153 13345 18187 13379
rect 18187 13345 18196 13379
rect 18144 13336 18196 13345
rect 20076 13336 20128 13388
rect 35808 13404 35860 13456
rect 38936 13404 38988 13456
rect 23480 13336 23532 13388
rect 25044 13379 25096 13388
rect 25044 13345 25053 13379
rect 25053 13345 25087 13379
rect 25087 13345 25096 13379
rect 25044 13336 25096 13345
rect 1860 13243 1912 13252
rect 1860 13209 1869 13243
rect 1869 13209 1903 13243
rect 1903 13209 1912 13243
rect 1860 13200 1912 13209
rect 11244 13132 11296 13184
rect 19432 13200 19484 13252
rect 21088 13268 21140 13320
rect 23848 13311 23900 13320
rect 23848 13277 23857 13311
rect 23857 13277 23891 13311
rect 23891 13277 23900 13311
rect 23848 13268 23900 13277
rect 24032 13311 24084 13320
rect 24032 13277 24041 13311
rect 24041 13277 24075 13311
rect 24075 13277 24084 13311
rect 24032 13268 24084 13277
rect 15568 13132 15620 13184
rect 15936 13132 15988 13184
rect 19800 13132 19852 13184
rect 19984 13175 20036 13184
rect 19984 13141 19993 13175
rect 19993 13141 20027 13175
rect 20027 13141 20036 13175
rect 19984 13132 20036 13141
rect 23388 13200 23440 13252
rect 21088 13132 21140 13184
rect 22008 13132 22060 13184
rect 24676 13268 24728 13320
rect 24952 13268 25004 13320
rect 25136 13311 25188 13320
rect 25136 13277 25145 13311
rect 25145 13277 25179 13311
rect 25179 13277 25188 13311
rect 25136 13268 25188 13277
rect 31576 13336 31628 13388
rect 28264 13311 28316 13320
rect 28264 13277 28273 13311
rect 28273 13277 28307 13311
rect 28307 13277 28316 13311
rect 28264 13268 28316 13277
rect 29092 13268 29144 13320
rect 28632 13200 28684 13252
rect 31576 13200 31628 13252
rect 32496 13268 32548 13320
rect 41604 13336 41656 13388
rect 43260 13472 43312 13524
rect 48412 13404 48464 13456
rect 58164 13379 58216 13388
rect 36268 13311 36320 13320
rect 36268 13277 36277 13311
rect 36277 13277 36311 13311
rect 36311 13277 36320 13311
rect 36268 13268 36320 13277
rect 36360 13268 36412 13320
rect 24952 13132 25004 13184
rect 29552 13132 29604 13184
rect 32128 13243 32180 13252
rect 32128 13209 32137 13243
rect 32137 13209 32171 13243
rect 32171 13209 32180 13243
rect 32128 13200 32180 13209
rect 32588 13200 32640 13252
rect 35992 13200 36044 13252
rect 32496 13132 32548 13184
rect 32864 13132 32916 13184
rect 34704 13132 34756 13184
rect 36636 13175 36688 13184
rect 36636 13141 36645 13175
rect 36645 13141 36679 13175
rect 36679 13141 36688 13175
rect 36636 13132 36688 13141
rect 37096 13132 37148 13184
rect 37280 13175 37332 13184
rect 37280 13141 37289 13175
rect 37289 13141 37323 13175
rect 37323 13141 37332 13175
rect 37832 13268 37884 13320
rect 38660 13311 38712 13320
rect 38660 13277 38669 13311
rect 38669 13277 38703 13311
rect 38703 13277 38712 13311
rect 38660 13268 38712 13277
rect 41420 13268 41472 13320
rect 42616 13311 42668 13320
rect 42616 13277 42625 13311
rect 42625 13277 42659 13311
rect 42659 13277 42668 13311
rect 42616 13268 42668 13277
rect 43168 13268 43220 13320
rect 58164 13345 58173 13379
rect 58173 13345 58207 13379
rect 58207 13345 58216 13379
rect 58164 13336 58216 13345
rect 56968 13311 57020 13320
rect 56968 13277 56977 13311
rect 56977 13277 57011 13311
rect 57011 13277 57020 13311
rect 56968 13268 57020 13277
rect 57888 13311 57940 13320
rect 57888 13277 57897 13311
rect 57897 13277 57931 13311
rect 57931 13277 57940 13311
rect 57888 13268 57940 13277
rect 38476 13200 38528 13252
rect 39304 13200 39356 13252
rect 37280 13132 37332 13141
rect 41696 13132 41748 13184
rect 44548 13200 44600 13252
rect 55864 13200 55916 13252
rect 42616 13132 42668 13184
rect 43720 13132 43772 13184
rect 44456 13132 44508 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 9772 12928 9824 12980
rect 11152 12971 11204 12980
rect 11152 12937 11161 12971
rect 11161 12937 11195 12971
rect 11195 12937 11204 12971
rect 11152 12928 11204 12937
rect 13544 12971 13596 12980
rect 13544 12937 13553 12971
rect 13553 12937 13587 12971
rect 13587 12937 13596 12971
rect 13544 12928 13596 12937
rect 15384 12971 15436 12980
rect 15384 12937 15393 12971
rect 15393 12937 15427 12971
rect 15427 12937 15436 12971
rect 15384 12928 15436 12937
rect 17224 12971 17276 12980
rect 17224 12937 17233 12971
rect 17233 12937 17267 12971
rect 17267 12937 17276 12971
rect 17224 12928 17276 12937
rect 17776 12928 17828 12980
rect 18144 12928 18196 12980
rect 11888 12903 11940 12912
rect 11888 12869 11897 12903
rect 11897 12869 11931 12903
rect 11931 12869 11940 12903
rect 11888 12860 11940 12869
rect 11980 12860 12032 12912
rect 12072 12835 12124 12844
rect 12072 12801 12081 12835
rect 12081 12801 12115 12835
rect 12115 12801 12124 12835
rect 12072 12792 12124 12801
rect 12624 12835 12676 12844
rect 12624 12801 12633 12835
rect 12633 12801 12667 12835
rect 12667 12801 12676 12835
rect 12624 12792 12676 12801
rect 8852 12724 8904 12776
rect 9496 12767 9548 12776
rect 9496 12733 9505 12767
rect 9505 12733 9539 12767
rect 9539 12733 9548 12767
rect 9496 12724 9548 12733
rect 15200 12860 15252 12912
rect 15936 12860 15988 12912
rect 14004 12835 14056 12844
rect 14004 12801 14013 12835
rect 14013 12801 14047 12835
rect 14047 12801 14056 12835
rect 14004 12792 14056 12801
rect 17316 12835 17368 12844
rect 13084 12767 13136 12776
rect 13084 12733 13093 12767
rect 13093 12733 13127 12767
rect 13127 12733 13136 12767
rect 13084 12724 13136 12733
rect 11244 12656 11296 12708
rect 16672 12656 16724 12708
rect 17316 12801 17325 12835
rect 17325 12801 17359 12835
rect 17359 12801 17368 12835
rect 17316 12792 17368 12801
rect 17868 12860 17920 12912
rect 19616 12860 19668 12912
rect 23020 12928 23072 12980
rect 23480 12928 23532 12980
rect 25136 12928 25188 12980
rect 26148 12928 26200 12980
rect 26240 12928 26292 12980
rect 28540 12928 28592 12980
rect 37188 12928 37240 12980
rect 40868 12928 40920 12980
rect 42800 12928 42852 12980
rect 43352 12928 43404 12980
rect 46664 12928 46716 12980
rect 57888 12928 57940 12980
rect 27804 12860 27856 12912
rect 28632 12903 28684 12912
rect 28632 12869 28641 12903
rect 28641 12869 28675 12903
rect 28675 12869 28684 12903
rect 28632 12860 28684 12869
rect 29736 12860 29788 12912
rect 33232 12860 33284 12912
rect 35992 12903 36044 12912
rect 22560 12792 22612 12844
rect 23020 12792 23072 12844
rect 24768 12835 24820 12844
rect 24768 12801 24777 12835
rect 24777 12801 24811 12835
rect 24811 12801 24820 12835
rect 24768 12792 24820 12801
rect 25412 12792 25464 12844
rect 26148 12792 26200 12844
rect 17408 12724 17460 12776
rect 20812 12767 20864 12776
rect 20812 12733 20821 12767
rect 20821 12733 20855 12767
rect 20855 12733 20864 12767
rect 20812 12724 20864 12733
rect 20904 12724 20956 12776
rect 27436 12835 27488 12844
rect 27436 12801 27445 12835
rect 27445 12801 27479 12835
rect 27479 12801 27488 12835
rect 27436 12792 27488 12801
rect 27620 12792 27672 12844
rect 30380 12792 30432 12844
rect 30932 12835 30984 12844
rect 30932 12801 30941 12835
rect 30941 12801 30975 12835
rect 30975 12801 30984 12835
rect 30932 12792 30984 12801
rect 31116 12835 31168 12844
rect 31116 12801 31125 12835
rect 31125 12801 31159 12835
rect 31159 12801 31168 12835
rect 31116 12792 31168 12801
rect 31392 12792 31444 12844
rect 32680 12835 32732 12844
rect 32680 12801 32689 12835
rect 32689 12801 32723 12835
rect 32723 12801 32732 12835
rect 32680 12792 32732 12801
rect 32956 12835 33008 12844
rect 32956 12801 32965 12835
rect 32965 12801 32999 12835
rect 32999 12801 33008 12835
rect 32956 12792 33008 12801
rect 35992 12869 36001 12903
rect 36001 12869 36035 12903
rect 36035 12869 36044 12903
rect 35992 12860 36044 12869
rect 38016 12860 38068 12912
rect 38200 12860 38252 12912
rect 43536 12860 43588 12912
rect 33968 12792 34020 12844
rect 34520 12792 34572 12844
rect 34704 12792 34756 12844
rect 35808 12835 35860 12844
rect 19432 12656 19484 12708
rect 19524 12656 19576 12708
rect 15016 12588 15068 12640
rect 21456 12588 21508 12640
rect 27068 12656 27120 12708
rect 28264 12656 28316 12708
rect 32864 12724 32916 12776
rect 33416 12767 33468 12776
rect 33416 12733 33425 12767
rect 33425 12733 33459 12767
rect 33459 12733 33468 12767
rect 33416 12724 33468 12733
rect 35808 12801 35817 12835
rect 35817 12801 35851 12835
rect 35851 12801 35860 12835
rect 35808 12792 35860 12801
rect 36268 12792 36320 12844
rect 36452 12792 36504 12844
rect 37832 12792 37884 12844
rect 41788 12835 41840 12844
rect 41788 12801 41797 12835
rect 41797 12801 41831 12835
rect 41831 12801 41840 12835
rect 41788 12792 41840 12801
rect 42064 12792 42116 12844
rect 37096 12724 37148 12776
rect 41144 12724 41196 12776
rect 43168 12724 43220 12776
rect 25504 12588 25556 12640
rect 25872 12588 25924 12640
rect 26608 12588 26660 12640
rect 27712 12631 27764 12640
rect 27712 12597 27721 12631
rect 27721 12597 27755 12631
rect 27755 12597 27764 12631
rect 27712 12588 27764 12597
rect 28172 12588 28224 12640
rect 28540 12588 28592 12640
rect 31024 12588 31076 12640
rect 31944 12656 31996 12708
rect 36360 12699 36412 12708
rect 36360 12665 36369 12699
rect 36369 12665 36403 12699
rect 36403 12665 36412 12699
rect 36360 12656 36412 12665
rect 31852 12588 31904 12640
rect 33232 12588 33284 12640
rect 33508 12588 33560 12640
rect 34520 12588 34572 12640
rect 37096 12588 37148 12640
rect 43444 12656 43496 12708
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 2228 12427 2280 12436
rect 2228 12393 2237 12427
rect 2237 12393 2271 12427
rect 2271 12393 2280 12427
rect 2228 12384 2280 12393
rect 10140 12384 10192 12436
rect 11428 12384 11480 12436
rect 11980 12384 12032 12436
rect 12256 12384 12308 12436
rect 13084 12384 13136 12436
rect 16120 12384 16172 12436
rect 16396 12384 16448 12436
rect 16672 12384 16724 12436
rect 19156 12384 19208 12436
rect 23480 12384 23532 12436
rect 25044 12384 25096 12436
rect 25412 12427 25464 12436
rect 25412 12393 25421 12427
rect 25421 12393 25455 12427
rect 25455 12393 25464 12427
rect 25412 12384 25464 12393
rect 25504 12384 25556 12436
rect 13728 12359 13780 12368
rect 10324 12248 10376 12300
rect 13728 12325 13737 12359
rect 13737 12325 13771 12359
rect 13771 12325 13780 12359
rect 13728 12316 13780 12325
rect 18512 12316 18564 12368
rect 18696 12316 18748 12368
rect 19432 12316 19484 12368
rect 23020 12316 23072 12368
rect 23388 12316 23440 12368
rect 24768 12316 24820 12368
rect 26516 12316 26568 12368
rect 28356 12384 28408 12436
rect 29828 12316 29880 12368
rect 32312 12384 32364 12436
rect 32680 12384 32732 12436
rect 32956 12384 33008 12436
rect 40776 12384 40828 12436
rect 10508 12223 10560 12232
rect 10508 12189 10517 12223
rect 10517 12189 10551 12223
rect 10551 12189 10560 12223
rect 10508 12180 10560 12189
rect 12072 12223 12124 12232
rect 12072 12189 12081 12223
rect 12081 12189 12115 12223
rect 12115 12189 12124 12223
rect 12072 12180 12124 12189
rect 11060 12112 11112 12164
rect 11888 12112 11940 12164
rect 12532 12180 12584 12232
rect 14924 12291 14976 12300
rect 14924 12257 14933 12291
rect 14933 12257 14967 12291
rect 14967 12257 14976 12291
rect 14924 12248 14976 12257
rect 15384 12180 15436 12232
rect 15660 12180 15712 12232
rect 15936 12223 15988 12232
rect 15936 12189 15945 12223
rect 15945 12189 15979 12223
rect 15979 12189 15988 12223
rect 15936 12180 15988 12189
rect 18144 12180 18196 12232
rect 18696 12223 18748 12232
rect 18696 12189 18705 12223
rect 18705 12189 18739 12223
rect 18739 12189 18748 12223
rect 18696 12180 18748 12189
rect 18880 12223 18932 12232
rect 18880 12189 18889 12223
rect 18889 12189 18923 12223
rect 18923 12189 18932 12223
rect 18880 12180 18932 12189
rect 19432 12223 19484 12232
rect 19432 12189 19441 12223
rect 19441 12189 19475 12223
rect 19475 12189 19484 12223
rect 19432 12180 19484 12189
rect 19616 12223 19668 12232
rect 19616 12189 19625 12223
rect 19625 12189 19659 12223
rect 19659 12189 19668 12223
rect 19616 12180 19668 12189
rect 16120 12112 16172 12164
rect 19984 12112 20036 12164
rect 11244 12044 11296 12096
rect 14740 12044 14792 12096
rect 15660 12044 15712 12096
rect 17868 12044 17920 12096
rect 18972 12044 19024 12096
rect 20536 12248 20588 12300
rect 23296 12248 23348 12300
rect 24860 12248 24912 12300
rect 25228 12248 25280 12300
rect 20904 12180 20956 12232
rect 23204 12180 23256 12232
rect 23756 12180 23808 12232
rect 24584 12223 24636 12232
rect 24584 12189 24593 12223
rect 24593 12189 24627 12223
rect 24627 12189 24636 12223
rect 24584 12180 24636 12189
rect 24768 12223 24820 12232
rect 24768 12189 24777 12223
rect 24777 12189 24811 12223
rect 24811 12189 24820 12223
rect 24768 12180 24820 12189
rect 25044 12180 25096 12232
rect 25872 12223 25924 12232
rect 25872 12189 25881 12223
rect 25881 12189 25915 12223
rect 25915 12189 25924 12223
rect 25872 12180 25924 12189
rect 26976 12248 27028 12300
rect 29092 12248 29144 12300
rect 28908 12180 28960 12232
rect 31484 12248 31536 12300
rect 31300 12223 31352 12232
rect 25412 12112 25464 12164
rect 26792 12112 26844 12164
rect 29184 12112 29236 12164
rect 31300 12189 31309 12223
rect 31309 12189 31343 12223
rect 31343 12189 31352 12223
rect 31300 12180 31352 12189
rect 31852 12248 31904 12300
rect 32496 12291 32548 12300
rect 32496 12257 32505 12291
rect 32505 12257 32539 12291
rect 32539 12257 32548 12291
rect 32496 12248 32548 12257
rect 35532 12248 35584 12300
rect 36636 12291 36688 12300
rect 31944 12223 31996 12232
rect 31944 12189 31953 12223
rect 31953 12189 31987 12223
rect 31987 12189 31996 12223
rect 31944 12180 31996 12189
rect 30472 12112 30524 12164
rect 20904 12044 20956 12096
rect 23020 12087 23072 12096
rect 23020 12053 23029 12087
rect 23029 12053 23063 12087
rect 23063 12053 23072 12087
rect 23020 12044 23072 12053
rect 23296 12044 23348 12096
rect 24308 12044 24360 12096
rect 24860 12044 24912 12096
rect 25504 12044 25556 12096
rect 26884 12044 26936 12096
rect 28448 12087 28500 12096
rect 28448 12053 28457 12087
rect 28457 12053 28491 12087
rect 28491 12053 28500 12087
rect 29920 12087 29972 12096
rect 28448 12044 28500 12053
rect 29920 12053 29929 12087
rect 29929 12053 29963 12087
rect 29963 12053 29972 12087
rect 29920 12044 29972 12053
rect 30840 12087 30892 12096
rect 30840 12053 30849 12087
rect 30849 12053 30883 12087
rect 30883 12053 30892 12087
rect 30840 12044 30892 12053
rect 31208 12087 31260 12096
rect 31208 12053 31217 12087
rect 31217 12053 31251 12087
rect 31251 12053 31260 12087
rect 31208 12044 31260 12053
rect 31392 12044 31444 12096
rect 32588 12180 32640 12232
rect 32956 12180 33008 12232
rect 34244 12180 34296 12232
rect 35348 12223 35400 12232
rect 35348 12189 35357 12223
rect 35357 12189 35391 12223
rect 35391 12189 35400 12223
rect 35348 12180 35400 12189
rect 35808 12180 35860 12232
rect 35900 12180 35952 12232
rect 36636 12257 36645 12291
rect 36645 12257 36679 12291
rect 36679 12257 36688 12291
rect 36636 12248 36688 12257
rect 41236 12316 41288 12368
rect 42340 12384 42392 12436
rect 40040 12223 40092 12232
rect 40040 12189 40049 12223
rect 40049 12189 40083 12223
rect 40083 12189 40092 12223
rect 40040 12180 40092 12189
rect 40132 12223 40184 12232
rect 40132 12189 40142 12223
rect 40142 12189 40176 12223
rect 40176 12189 40184 12223
rect 40132 12180 40184 12189
rect 33876 12112 33928 12164
rect 38016 12155 38068 12164
rect 38016 12121 38025 12155
rect 38025 12121 38059 12155
rect 38059 12121 38068 12155
rect 38016 12112 38068 12121
rect 40592 12180 40644 12232
rect 41236 12180 41288 12232
rect 37924 12044 37976 12096
rect 41420 12112 41472 12164
rect 42064 12180 42116 12232
rect 44640 12316 44692 12368
rect 57888 12223 57940 12232
rect 42248 12112 42300 12164
rect 57888 12189 57897 12223
rect 57897 12189 57931 12223
rect 57931 12189 57940 12223
rect 57888 12180 57940 12189
rect 43352 12112 43404 12164
rect 43720 12112 43772 12164
rect 58164 12155 58216 12164
rect 58164 12121 58173 12155
rect 58173 12121 58207 12155
rect 58207 12121 58216 12155
rect 58164 12112 58216 12121
rect 43260 12044 43312 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 9496 11840 9548 11892
rect 14004 11840 14056 11892
rect 15936 11840 15988 11892
rect 1860 11815 1912 11824
rect 1860 11781 1869 11815
rect 1869 11781 1903 11815
rect 1903 11781 1912 11815
rect 1860 11772 1912 11781
rect 10508 11747 10560 11756
rect 10508 11713 10517 11747
rect 10517 11713 10551 11747
rect 10551 11713 10560 11747
rect 10508 11704 10560 11713
rect 11060 11772 11112 11824
rect 12256 11772 12308 11824
rect 13268 11772 13320 11824
rect 13636 11772 13688 11824
rect 11888 11747 11940 11756
rect 11888 11713 11897 11747
rect 11897 11713 11931 11747
rect 11931 11713 11940 11747
rect 11888 11704 11940 11713
rect 12348 11704 12400 11756
rect 14924 11704 14976 11756
rect 11796 11568 11848 11620
rect 12164 11679 12216 11688
rect 12164 11645 12173 11679
rect 12173 11645 12207 11679
rect 12207 11645 12216 11679
rect 12164 11636 12216 11645
rect 14832 11636 14884 11688
rect 17408 11840 17460 11892
rect 19432 11840 19484 11892
rect 19892 11840 19944 11892
rect 20076 11840 20128 11892
rect 20904 11840 20956 11892
rect 22376 11883 22428 11892
rect 22376 11849 22385 11883
rect 22385 11849 22419 11883
rect 22419 11849 22428 11883
rect 22376 11840 22428 11849
rect 22744 11840 22796 11892
rect 23480 11840 23532 11892
rect 25228 11840 25280 11892
rect 26792 11840 26844 11892
rect 29920 11840 29972 11892
rect 17776 11772 17828 11824
rect 18880 11772 18932 11824
rect 16672 11704 16724 11756
rect 16856 11747 16908 11756
rect 16856 11713 16865 11747
rect 16865 11713 16899 11747
rect 16899 11713 16908 11747
rect 16856 11704 16908 11713
rect 17408 11704 17460 11756
rect 19800 11704 19852 11756
rect 15292 11679 15344 11688
rect 15292 11645 15301 11679
rect 15301 11645 15335 11679
rect 15335 11645 15344 11679
rect 15292 11636 15344 11645
rect 15660 11636 15712 11688
rect 10324 11500 10376 11552
rect 13176 11500 13228 11552
rect 13360 11543 13412 11552
rect 13360 11509 13369 11543
rect 13369 11509 13403 11543
rect 13403 11509 13412 11543
rect 13360 11500 13412 11509
rect 15660 11500 15712 11552
rect 16396 11500 16448 11552
rect 18880 11568 18932 11620
rect 19156 11636 19208 11688
rect 20536 11704 20588 11756
rect 21088 11772 21140 11824
rect 23020 11704 23072 11756
rect 25412 11772 25464 11824
rect 30288 11772 30340 11824
rect 30840 11772 30892 11824
rect 32864 11772 32916 11824
rect 25228 11747 25280 11756
rect 18696 11500 18748 11552
rect 19248 11568 19300 11620
rect 19708 11568 19760 11620
rect 20076 11568 20128 11620
rect 20352 11568 20404 11620
rect 20812 11568 20864 11620
rect 22284 11636 22336 11688
rect 24676 11636 24728 11688
rect 25228 11713 25237 11747
rect 25237 11713 25271 11747
rect 25271 11713 25280 11747
rect 25228 11704 25280 11713
rect 25504 11704 25556 11756
rect 26240 11747 26292 11756
rect 26240 11713 26249 11747
rect 26249 11713 26283 11747
rect 26283 11713 26292 11747
rect 26240 11704 26292 11713
rect 26424 11747 26476 11756
rect 26424 11713 26433 11747
rect 26433 11713 26467 11747
rect 26467 11713 26476 11747
rect 26424 11704 26476 11713
rect 30472 11747 30524 11756
rect 30472 11713 30481 11747
rect 30481 11713 30515 11747
rect 30515 11713 30524 11747
rect 30472 11704 30524 11713
rect 30932 11704 30984 11756
rect 25412 11679 25464 11688
rect 25412 11645 25421 11679
rect 25421 11645 25455 11679
rect 25455 11645 25464 11679
rect 25412 11636 25464 11645
rect 25596 11679 25648 11688
rect 25596 11645 25605 11679
rect 25605 11645 25639 11679
rect 25639 11645 25648 11679
rect 25596 11636 25648 11645
rect 27344 11636 27396 11688
rect 27436 11636 27488 11688
rect 32312 11704 32364 11756
rect 34152 11772 34204 11824
rect 33140 11704 33192 11756
rect 33968 11704 34020 11756
rect 35900 11772 35952 11824
rect 37188 11840 37240 11892
rect 39120 11772 39172 11824
rect 44180 11840 44232 11892
rect 46296 11840 46348 11892
rect 59084 11840 59136 11892
rect 40592 11772 40644 11824
rect 42892 11772 42944 11824
rect 35348 11704 35400 11756
rect 38752 11747 38804 11756
rect 38752 11713 38761 11747
rect 38761 11713 38795 11747
rect 38795 11713 38804 11747
rect 38752 11704 38804 11713
rect 38936 11704 38988 11756
rect 31484 11636 31536 11688
rect 31852 11636 31904 11688
rect 32772 11636 32824 11688
rect 23756 11568 23808 11620
rect 19524 11500 19576 11552
rect 31208 11568 31260 11620
rect 31944 11568 31996 11620
rect 32404 11568 32456 11620
rect 33140 11568 33192 11620
rect 41236 11636 41288 11688
rect 42064 11704 42116 11756
rect 43076 11704 43128 11756
rect 43260 11747 43312 11756
rect 43260 11713 43269 11747
rect 43269 11713 43303 11747
rect 43303 11713 43312 11747
rect 43260 11704 43312 11713
rect 43996 11772 44048 11824
rect 44272 11772 44324 11824
rect 50712 11772 50764 11824
rect 41420 11636 41472 11688
rect 41512 11636 41564 11688
rect 42708 11636 42760 11688
rect 43720 11679 43772 11688
rect 43720 11645 43729 11679
rect 43729 11645 43763 11679
rect 43763 11645 43772 11679
rect 43720 11636 43772 11645
rect 45192 11704 45244 11756
rect 45468 11747 45520 11756
rect 45468 11713 45477 11747
rect 45477 11713 45511 11747
rect 45511 11713 45520 11747
rect 45468 11704 45520 11713
rect 45560 11704 45612 11756
rect 46112 11704 46164 11756
rect 57152 11747 57204 11756
rect 57152 11713 57161 11747
rect 57161 11713 57195 11747
rect 57195 11713 57204 11747
rect 57152 11704 57204 11713
rect 24032 11500 24084 11552
rect 24768 11500 24820 11552
rect 26700 11500 26752 11552
rect 31300 11500 31352 11552
rect 32128 11500 32180 11552
rect 32220 11500 32272 11552
rect 38016 11568 38068 11620
rect 35808 11500 35860 11552
rect 39856 11500 39908 11552
rect 42064 11500 42116 11552
rect 42708 11543 42760 11552
rect 42708 11509 42717 11543
rect 42717 11509 42751 11543
rect 42751 11509 42760 11543
rect 42708 11500 42760 11509
rect 43168 11500 43220 11552
rect 57428 11568 57480 11620
rect 46848 11543 46900 11552
rect 46848 11509 46857 11543
rect 46857 11509 46891 11543
rect 46891 11509 46900 11543
rect 46848 11500 46900 11509
rect 48320 11500 48372 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 1768 11203 1820 11212
rect 1768 11169 1777 11203
rect 1777 11169 1811 11203
rect 1811 11169 1820 11203
rect 1768 11160 1820 11169
rect 11888 11296 11940 11348
rect 16764 11296 16816 11348
rect 18052 11339 18104 11348
rect 18052 11305 18061 11339
rect 18061 11305 18095 11339
rect 18095 11305 18104 11339
rect 18052 11296 18104 11305
rect 19340 11296 19392 11348
rect 20260 11296 20312 11348
rect 20352 11296 20404 11348
rect 21088 11296 21140 11348
rect 11704 11160 11756 11212
rect 13176 11203 13228 11212
rect 13176 11169 13185 11203
rect 13185 11169 13219 11203
rect 13219 11169 13228 11203
rect 13176 11160 13228 11169
rect 14832 11203 14884 11212
rect 14832 11169 14841 11203
rect 14841 11169 14875 11203
rect 14875 11169 14884 11203
rect 14832 11160 14884 11169
rect 20628 11228 20680 11280
rect 17868 11203 17920 11212
rect 2872 11024 2924 11076
rect 8576 11024 8628 11076
rect 11428 11135 11480 11144
rect 11428 11101 11437 11135
rect 11437 11101 11471 11135
rect 11471 11101 11480 11135
rect 11428 11092 11480 11101
rect 15016 11135 15068 11144
rect 15016 11101 15025 11135
rect 15025 11101 15059 11135
rect 15059 11101 15068 11135
rect 15016 11092 15068 11101
rect 16396 11135 16448 11144
rect 16396 11101 16405 11135
rect 16405 11101 16439 11135
rect 16439 11101 16448 11135
rect 16396 11092 16448 11101
rect 16580 11135 16632 11144
rect 16580 11101 16589 11135
rect 16589 11101 16623 11135
rect 16623 11101 16632 11135
rect 16580 11092 16632 11101
rect 16672 11092 16724 11144
rect 17868 11169 17877 11203
rect 17877 11169 17911 11203
rect 17911 11169 17920 11203
rect 17868 11160 17920 11169
rect 17960 11160 18012 11212
rect 19524 11160 19576 11212
rect 23848 11228 23900 11280
rect 25228 11296 25280 11348
rect 24308 11228 24360 11280
rect 24584 11228 24636 11280
rect 25688 11228 25740 11280
rect 26148 11296 26200 11348
rect 27804 11296 27856 11348
rect 29000 11296 29052 11348
rect 30472 11296 30524 11348
rect 35348 11339 35400 11348
rect 35348 11305 35357 11339
rect 35357 11305 35391 11339
rect 35391 11305 35400 11339
rect 35348 11296 35400 11305
rect 36544 11296 36596 11348
rect 26056 11228 26108 11280
rect 29736 11228 29788 11280
rect 29828 11228 29880 11280
rect 30288 11160 30340 11212
rect 30748 11203 30800 11212
rect 30748 11169 30757 11203
rect 30757 11169 30791 11203
rect 30791 11169 30800 11203
rect 30748 11160 30800 11169
rect 32404 11228 32456 11280
rect 36084 11228 36136 11280
rect 39856 11228 39908 11280
rect 1584 10956 1636 11008
rect 15752 10999 15804 11008
rect 15752 10965 15761 10999
rect 15761 10965 15795 10999
rect 15795 10965 15804 10999
rect 15752 10956 15804 10965
rect 17132 11024 17184 11076
rect 17592 11092 17644 11144
rect 19432 11092 19484 11144
rect 19892 11135 19944 11144
rect 19892 11101 19915 11135
rect 19915 11101 19944 11135
rect 19892 11092 19944 11101
rect 23020 11135 23072 11144
rect 23020 11101 23029 11135
rect 23029 11101 23063 11135
rect 23063 11101 23072 11135
rect 23020 11092 23072 11101
rect 23112 11092 23164 11144
rect 23756 11135 23808 11144
rect 23756 11101 23765 11135
rect 23765 11101 23799 11135
rect 23799 11101 23808 11135
rect 23756 11092 23808 11101
rect 24492 11092 24544 11144
rect 22744 11024 22796 11076
rect 23940 11024 23992 11076
rect 24676 11092 24728 11144
rect 26056 11135 26108 11144
rect 26056 11101 26065 11135
rect 26065 11101 26099 11135
rect 26099 11101 26108 11135
rect 26056 11092 26108 11101
rect 26148 11092 26200 11144
rect 28908 11092 28960 11144
rect 29000 11092 29052 11144
rect 31116 11092 31168 11144
rect 31484 11092 31536 11144
rect 31852 11160 31904 11212
rect 32496 11160 32548 11212
rect 35808 11203 35860 11212
rect 32128 11135 32180 11144
rect 32128 11101 32137 11135
rect 32137 11101 32171 11135
rect 32171 11101 32180 11135
rect 32128 11092 32180 11101
rect 32312 11092 32364 11144
rect 25688 11024 25740 11076
rect 27712 11024 27764 11076
rect 35808 11169 35817 11203
rect 35817 11169 35851 11203
rect 35851 11169 35860 11203
rect 35808 11160 35860 11169
rect 35992 11203 36044 11212
rect 35992 11169 36001 11203
rect 36001 11169 36035 11203
rect 36035 11169 36044 11203
rect 35992 11160 36044 11169
rect 33784 11135 33836 11144
rect 33784 11101 33793 11135
rect 33793 11101 33827 11135
rect 33827 11101 33836 11135
rect 33784 11092 33836 11101
rect 34060 11135 34112 11144
rect 34060 11101 34069 11135
rect 34069 11101 34103 11135
rect 34103 11101 34112 11135
rect 34060 11092 34112 11101
rect 34428 11092 34480 11144
rect 35716 11135 35768 11144
rect 35716 11101 35725 11135
rect 35725 11101 35759 11135
rect 35759 11101 35768 11135
rect 35716 11092 35768 11101
rect 33876 11024 33928 11076
rect 38936 11160 38988 11212
rect 41328 11296 41380 11348
rect 46112 11339 46164 11348
rect 42064 11228 42116 11280
rect 43076 11271 43128 11280
rect 38384 11092 38436 11144
rect 39948 11092 40000 11144
rect 42248 11160 42300 11212
rect 42432 11135 42484 11144
rect 36360 11024 36412 11076
rect 37096 11024 37148 11076
rect 38660 11024 38712 11076
rect 41144 11024 41196 11076
rect 42432 11101 42441 11135
rect 42441 11101 42475 11135
rect 42475 11101 42484 11135
rect 42432 11092 42484 11101
rect 42616 11135 42668 11144
rect 42616 11101 42623 11135
rect 42623 11101 42668 11135
rect 42616 11092 42668 11101
rect 43076 11237 43085 11271
rect 43085 11237 43119 11271
rect 43119 11237 43128 11271
rect 43076 11228 43128 11237
rect 46112 11305 46121 11339
rect 46121 11305 46155 11339
rect 46155 11305 46164 11339
rect 46112 11296 46164 11305
rect 42892 11135 42944 11144
rect 46572 11228 46624 11280
rect 42892 11101 42906 11135
rect 42906 11101 42940 11135
rect 42940 11101 42944 11135
rect 42892 11092 42944 11101
rect 44456 11135 44508 11144
rect 44456 11101 44465 11135
rect 44465 11101 44499 11135
rect 44499 11101 44508 11135
rect 44456 11092 44508 11101
rect 45100 11092 45152 11144
rect 46296 11092 46348 11144
rect 46756 11092 46808 11144
rect 57888 11228 57940 11280
rect 56876 11135 56928 11144
rect 56876 11101 56885 11135
rect 56885 11101 56919 11135
rect 56919 11101 56928 11135
rect 56876 11092 56928 11101
rect 46848 11024 46900 11076
rect 56140 11067 56192 11076
rect 56140 11033 56149 11067
rect 56149 11033 56183 11067
rect 56183 11033 56192 11067
rect 56140 11024 56192 11033
rect 56968 11024 57020 11076
rect 24584 10956 24636 11008
rect 24676 10956 24728 11008
rect 31300 10956 31352 11008
rect 31484 10956 31536 11008
rect 32772 10956 32824 11008
rect 34060 10956 34112 11008
rect 34336 10999 34388 11008
rect 34336 10965 34345 10999
rect 34345 10965 34379 10999
rect 34379 10965 34388 10999
rect 34336 10956 34388 10965
rect 36084 10956 36136 11008
rect 40960 10956 41012 11008
rect 42064 10956 42116 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 1676 10752 1728 10804
rect 1860 10727 1912 10736
rect 1860 10693 1869 10727
rect 1869 10693 1903 10727
rect 1903 10693 1912 10727
rect 1860 10684 1912 10693
rect 7380 10752 7432 10804
rect 12164 10795 12216 10804
rect 12164 10761 12173 10795
rect 12173 10761 12207 10795
rect 12207 10761 12216 10795
rect 12164 10752 12216 10761
rect 1584 10659 1636 10668
rect 1584 10625 1593 10659
rect 1593 10625 1627 10659
rect 1627 10625 1636 10659
rect 1584 10616 1636 10625
rect 12716 10616 12768 10668
rect 12900 10659 12952 10668
rect 12900 10625 12909 10659
rect 12909 10625 12943 10659
rect 12943 10625 12952 10659
rect 12900 10616 12952 10625
rect 13360 10616 13412 10668
rect 15292 10616 15344 10668
rect 9496 10591 9548 10600
rect 9496 10557 9505 10591
rect 9505 10557 9539 10591
rect 9539 10557 9548 10591
rect 9496 10548 9548 10557
rect 9680 10591 9732 10600
rect 9680 10557 9689 10591
rect 9689 10557 9723 10591
rect 9723 10557 9732 10591
rect 11704 10591 11756 10600
rect 9680 10548 9732 10557
rect 11704 10557 11713 10591
rect 11713 10557 11747 10591
rect 11747 10557 11756 10591
rect 11704 10548 11756 10557
rect 12256 10548 12308 10600
rect 25044 10752 25096 10804
rect 15844 10684 15896 10736
rect 16212 10684 16264 10736
rect 16488 10684 16540 10736
rect 17040 10727 17092 10736
rect 17040 10693 17049 10727
rect 17049 10693 17083 10727
rect 17083 10693 17092 10727
rect 17040 10684 17092 10693
rect 17960 10684 18012 10736
rect 15660 10616 15712 10668
rect 17316 10616 17368 10668
rect 16212 10591 16264 10600
rect 11152 10480 11204 10532
rect 13176 10480 13228 10532
rect 15200 10523 15252 10532
rect 15200 10489 15209 10523
rect 15209 10489 15243 10523
rect 15243 10489 15252 10523
rect 15200 10480 15252 10489
rect 12164 10412 12216 10464
rect 16212 10557 16221 10591
rect 16221 10557 16255 10591
rect 16255 10557 16264 10591
rect 16212 10548 16264 10557
rect 16488 10548 16540 10600
rect 17132 10548 17184 10600
rect 20628 10684 20680 10736
rect 18972 10591 19024 10600
rect 18972 10557 18981 10591
rect 18981 10557 19015 10591
rect 19015 10557 19024 10591
rect 20536 10616 20588 10668
rect 18972 10548 19024 10557
rect 19432 10548 19484 10600
rect 23388 10684 23440 10736
rect 26424 10752 26476 10804
rect 28448 10752 28500 10804
rect 29092 10752 29144 10804
rect 30288 10752 30340 10804
rect 32128 10752 32180 10804
rect 27620 10684 27672 10736
rect 29828 10684 29880 10736
rect 25872 10659 25924 10668
rect 23480 10548 23532 10600
rect 19524 10480 19576 10532
rect 21916 10480 21968 10532
rect 24952 10480 25004 10532
rect 25320 10523 25372 10532
rect 25320 10489 25329 10523
rect 25329 10489 25363 10523
rect 25363 10489 25372 10523
rect 25320 10480 25372 10489
rect 25872 10625 25881 10659
rect 25881 10625 25915 10659
rect 25915 10625 25924 10659
rect 25872 10616 25924 10625
rect 25964 10591 26016 10600
rect 25964 10557 25973 10591
rect 25973 10557 26007 10591
rect 26007 10557 26016 10591
rect 25964 10548 26016 10557
rect 26056 10480 26108 10532
rect 27252 10480 27304 10532
rect 21180 10412 21232 10464
rect 22100 10412 22152 10464
rect 23664 10412 23716 10464
rect 24308 10412 24360 10464
rect 24492 10455 24544 10464
rect 24492 10421 24501 10455
rect 24501 10421 24535 10455
rect 24535 10421 24544 10455
rect 24492 10412 24544 10421
rect 24676 10412 24728 10464
rect 28448 10616 28500 10668
rect 29920 10616 29972 10668
rect 31024 10616 31076 10668
rect 31484 10616 31536 10668
rect 34336 10684 34388 10736
rect 34980 10752 35032 10804
rect 39396 10752 39448 10804
rect 41144 10795 41196 10804
rect 41144 10761 41153 10795
rect 41153 10761 41187 10795
rect 41187 10761 41196 10795
rect 41144 10752 41196 10761
rect 49424 10752 49476 10804
rect 27804 10591 27856 10600
rect 27804 10557 27813 10591
rect 27813 10557 27847 10591
rect 27847 10557 27856 10591
rect 27804 10548 27856 10557
rect 28172 10548 28224 10600
rect 29092 10548 29144 10600
rect 31760 10591 31812 10600
rect 31760 10557 31769 10591
rect 31769 10557 31803 10591
rect 31803 10557 31812 10591
rect 31760 10548 31812 10557
rect 32588 10548 32640 10600
rect 34796 10548 34848 10600
rect 35256 10616 35308 10668
rect 35532 10616 35584 10668
rect 42064 10684 42116 10736
rect 42892 10684 42944 10736
rect 54024 10752 54076 10804
rect 56968 10752 57020 10804
rect 53380 10727 53432 10736
rect 37740 10591 37792 10600
rect 37740 10557 37749 10591
rect 37749 10557 37783 10591
rect 37783 10557 37792 10591
rect 37740 10548 37792 10557
rect 38016 10548 38068 10600
rect 38660 10548 38712 10600
rect 38752 10548 38804 10600
rect 39120 10548 39172 10600
rect 41972 10616 42024 10668
rect 44180 10659 44232 10668
rect 44180 10625 44189 10659
rect 44189 10625 44223 10659
rect 44223 10625 44232 10659
rect 44180 10616 44232 10625
rect 46848 10616 46900 10668
rect 53380 10693 53389 10727
rect 53389 10693 53423 10727
rect 53423 10693 53432 10727
rect 53380 10684 53432 10693
rect 53472 10659 53524 10668
rect 46572 10548 46624 10600
rect 53472 10625 53481 10659
rect 53481 10625 53515 10659
rect 53515 10625 53524 10659
rect 53472 10616 53524 10625
rect 54300 10616 54352 10668
rect 57060 10616 57112 10668
rect 57888 10616 57940 10668
rect 54208 10548 54260 10600
rect 28356 10480 28408 10532
rect 27804 10412 27856 10464
rect 29184 10412 29236 10464
rect 29736 10412 29788 10464
rect 30288 10455 30340 10464
rect 30288 10421 30297 10455
rect 30297 10421 30331 10455
rect 30331 10421 30340 10455
rect 30288 10412 30340 10421
rect 33324 10480 33376 10532
rect 34980 10412 35032 10464
rect 35348 10412 35400 10464
rect 38108 10412 38160 10464
rect 44824 10412 44876 10464
rect 45192 10412 45244 10464
rect 45652 10412 45704 10464
rect 53472 10412 53524 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 11428 10208 11480 10260
rect 11336 10183 11388 10192
rect 11336 10149 11345 10183
rect 11345 10149 11379 10183
rect 11379 10149 11388 10183
rect 11336 10140 11388 10149
rect 1768 10115 1820 10124
rect 1768 10081 1777 10115
rect 1777 10081 1811 10115
rect 1811 10081 1820 10115
rect 1768 10072 1820 10081
rect 2596 10072 2648 10124
rect 13176 10140 13228 10192
rect 13820 10208 13872 10260
rect 16212 10140 16264 10192
rect 17684 10140 17736 10192
rect 17868 10140 17920 10192
rect 19340 10140 19392 10192
rect 19524 10208 19576 10260
rect 21088 10208 21140 10260
rect 23664 10208 23716 10260
rect 24492 10208 24544 10260
rect 19800 10140 19852 10192
rect 21640 10183 21692 10192
rect 21640 10149 21649 10183
rect 21649 10149 21683 10183
rect 21683 10149 21692 10183
rect 21640 10140 21692 10149
rect 23480 10183 23532 10192
rect 23480 10149 23489 10183
rect 23489 10149 23523 10183
rect 23523 10149 23532 10183
rect 23480 10140 23532 10149
rect 11704 9936 11756 9988
rect 13452 10004 13504 10056
rect 15108 10072 15160 10124
rect 15292 10072 15344 10124
rect 12900 9936 12952 9988
rect 13360 9936 13412 9988
rect 15660 10004 15712 10056
rect 18696 10072 18748 10124
rect 18788 10115 18840 10124
rect 18788 10081 18797 10115
rect 18797 10081 18831 10115
rect 18831 10081 18840 10115
rect 18788 10072 18840 10081
rect 21824 10072 21876 10124
rect 22284 10072 22336 10124
rect 25136 10208 25188 10260
rect 15292 9936 15344 9988
rect 1952 9868 2004 9920
rect 14188 9868 14240 9920
rect 16488 10004 16540 10056
rect 16672 10047 16724 10056
rect 16672 10013 16681 10047
rect 16681 10013 16715 10047
rect 16715 10013 16724 10047
rect 16672 10004 16724 10013
rect 17408 10004 17460 10056
rect 19156 10004 19208 10056
rect 19432 10004 19484 10056
rect 20996 10004 21048 10056
rect 19616 9936 19668 9988
rect 21640 9936 21692 9988
rect 21824 9936 21876 9988
rect 24584 10047 24636 10056
rect 24584 10013 24593 10047
rect 24593 10013 24627 10047
rect 24627 10013 24636 10047
rect 24584 10004 24636 10013
rect 23664 9979 23716 9988
rect 23664 9945 23673 9979
rect 23673 9945 23707 9979
rect 23707 9945 23716 9979
rect 23664 9936 23716 9945
rect 24768 10140 24820 10192
rect 26516 10208 26568 10260
rect 28172 10251 28224 10260
rect 28172 10217 28181 10251
rect 28181 10217 28215 10251
rect 28215 10217 28224 10251
rect 28172 10208 28224 10217
rect 25320 10140 25372 10192
rect 31484 10208 31536 10260
rect 32220 10208 32272 10260
rect 34428 10208 34480 10260
rect 35532 10208 35584 10260
rect 36912 10208 36964 10260
rect 38752 10208 38804 10260
rect 45468 10208 45520 10260
rect 48780 10208 48832 10260
rect 28816 10140 28868 10192
rect 30656 10140 30708 10192
rect 30748 10140 30800 10192
rect 33876 10140 33928 10192
rect 37740 10140 37792 10192
rect 38614 10140 38666 10192
rect 26240 10072 26292 10124
rect 26884 10072 26936 10124
rect 25136 10047 25188 10056
rect 25136 10013 25145 10047
rect 25145 10013 25179 10047
rect 25179 10013 25188 10047
rect 25136 10004 25188 10013
rect 27252 10047 27304 10056
rect 27252 10013 27261 10047
rect 27261 10013 27295 10047
rect 27295 10013 27304 10047
rect 27252 10004 27304 10013
rect 27988 10047 28040 10056
rect 27988 10013 27997 10047
rect 27997 10013 28031 10047
rect 28031 10013 28040 10047
rect 27988 10004 28040 10013
rect 28816 10047 28868 10056
rect 28816 10013 28825 10047
rect 28825 10013 28859 10047
rect 28859 10013 28868 10047
rect 28816 10004 28868 10013
rect 28908 10004 28960 10056
rect 30012 10047 30064 10056
rect 30012 10013 30021 10047
rect 30021 10013 30055 10047
rect 30055 10013 30064 10047
rect 30196 10047 30248 10056
rect 30012 10004 30064 10013
rect 30196 10013 30205 10047
rect 30205 10013 30239 10047
rect 30239 10013 30248 10047
rect 30196 10004 30248 10013
rect 30472 10004 30524 10056
rect 32036 10072 32088 10124
rect 32956 10072 33008 10124
rect 32128 10047 32180 10056
rect 32128 10013 32137 10047
rect 32137 10013 32171 10047
rect 32171 10013 32180 10047
rect 32128 10004 32180 10013
rect 32404 10047 32456 10056
rect 32404 10013 32413 10047
rect 32413 10013 32447 10047
rect 32447 10013 32456 10047
rect 32404 10004 32456 10013
rect 33324 10047 33376 10056
rect 33324 10013 33333 10047
rect 33333 10013 33367 10047
rect 33367 10013 33376 10047
rect 33324 10004 33376 10013
rect 33416 10047 33468 10056
rect 33416 10013 33426 10047
rect 33426 10013 33460 10047
rect 33460 10013 33468 10047
rect 34244 10072 34296 10124
rect 34796 10072 34848 10124
rect 35348 10072 35400 10124
rect 36636 10072 36688 10124
rect 33416 10004 33468 10013
rect 24952 9979 25004 9988
rect 18972 9868 19024 9920
rect 20536 9868 20588 9920
rect 24952 9945 24979 9979
rect 24979 9945 25004 9979
rect 25596 9979 25648 9988
rect 24952 9936 25004 9945
rect 25596 9945 25605 9979
rect 25605 9945 25639 9979
rect 25639 9945 25648 9979
rect 25596 9936 25648 9945
rect 25780 9936 25832 9988
rect 27620 9936 27672 9988
rect 29828 9936 29880 9988
rect 30104 9936 30156 9988
rect 31116 9936 31168 9988
rect 33692 9979 33744 9988
rect 33692 9945 33701 9979
rect 33701 9945 33735 9979
rect 33735 9945 33744 9979
rect 33692 9936 33744 9945
rect 29552 9868 29604 9920
rect 31208 9868 31260 9920
rect 32220 9868 32272 9920
rect 34152 9936 34204 9988
rect 36912 10004 36964 10056
rect 37372 10047 37424 10056
rect 37372 10013 37381 10047
rect 37381 10013 37415 10047
rect 37415 10013 37424 10047
rect 37372 10004 37424 10013
rect 37464 10047 37516 10056
rect 37464 10013 37473 10047
rect 37473 10013 37507 10047
rect 37507 10013 37516 10047
rect 41236 10072 41288 10124
rect 37464 10004 37516 10013
rect 35164 9979 35216 9988
rect 35164 9945 35173 9979
rect 35173 9945 35207 9979
rect 35207 9945 35216 9979
rect 35164 9936 35216 9945
rect 35348 9979 35400 9988
rect 35348 9945 35357 9979
rect 35357 9945 35391 9979
rect 35391 9945 35400 9979
rect 35348 9936 35400 9945
rect 37740 9936 37792 9988
rect 38384 10047 38436 10056
rect 38384 10013 38393 10047
rect 38393 10013 38427 10047
rect 38427 10013 38436 10047
rect 38384 10004 38436 10013
rect 38568 10004 38620 10056
rect 41052 10004 41104 10056
rect 44088 10047 44140 10056
rect 44088 10013 44097 10047
rect 44097 10013 44131 10047
rect 44131 10013 44140 10047
rect 44088 10004 44140 10013
rect 44548 10140 44600 10192
rect 44824 10072 44876 10124
rect 45652 10072 45704 10124
rect 46664 10072 46716 10124
rect 39396 9936 39448 9988
rect 46112 10004 46164 10056
rect 46848 10047 46900 10056
rect 46848 10013 46857 10047
rect 46857 10013 46891 10047
rect 46891 10013 46900 10047
rect 46848 10004 46900 10013
rect 36176 9868 36228 9920
rect 37464 9868 37516 9920
rect 38568 9868 38620 9920
rect 40316 9868 40368 9920
rect 40776 9868 40828 9920
rect 45468 9868 45520 9920
rect 46296 9868 46348 9920
rect 58164 10115 58216 10124
rect 58164 10081 58173 10115
rect 58173 10081 58207 10115
rect 58207 10081 58216 10115
rect 58164 10072 58216 10081
rect 56508 10004 56560 10056
rect 57060 9979 57112 9988
rect 57060 9945 57069 9979
rect 57069 9945 57103 9979
rect 57103 9945 57112 9979
rect 57060 9936 57112 9945
rect 51724 9868 51776 9920
rect 57152 9911 57204 9920
rect 57152 9877 57161 9911
rect 57161 9877 57195 9911
rect 57195 9877 57204 9911
rect 57152 9868 57204 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 11244 9596 11296 9648
rect 13544 9596 13596 9648
rect 1584 9571 1636 9580
rect 1584 9537 1593 9571
rect 1593 9537 1627 9571
rect 1627 9537 1636 9571
rect 1584 9528 1636 9537
rect 13360 9571 13412 9580
rect 13360 9537 13369 9571
rect 13369 9537 13403 9571
rect 13403 9537 13412 9571
rect 13360 9528 13412 9537
rect 13452 9571 13504 9580
rect 13452 9537 13461 9571
rect 13461 9537 13495 9571
rect 13495 9537 13504 9571
rect 15108 9596 15160 9648
rect 16396 9664 16448 9716
rect 17408 9664 17460 9716
rect 18604 9664 18656 9716
rect 18788 9664 18840 9716
rect 13452 9528 13504 9537
rect 14188 9571 14240 9580
rect 14188 9537 14197 9571
rect 14197 9537 14231 9571
rect 14231 9537 14240 9571
rect 14188 9528 14240 9537
rect 1768 9503 1820 9512
rect 1768 9469 1777 9503
rect 1777 9469 1811 9503
rect 1811 9469 1820 9503
rect 1768 9460 1820 9469
rect 8760 9503 8812 9512
rect 8760 9469 8769 9503
rect 8769 9469 8803 9503
rect 8803 9469 8812 9503
rect 8760 9460 8812 9469
rect 9680 9460 9732 9512
rect 13268 9460 13320 9512
rect 14280 9503 14332 9512
rect 14280 9469 14289 9503
rect 14289 9469 14323 9503
rect 14323 9469 14332 9503
rect 14280 9460 14332 9469
rect 7196 9392 7248 9444
rect 12716 9324 12768 9376
rect 13176 9367 13228 9376
rect 13176 9333 13185 9367
rect 13185 9333 13219 9367
rect 13219 9333 13228 9367
rect 13176 9324 13228 9333
rect 13636 9324 13688 9376
rect 15568 9571 15620 9580
rect 15568 9537 15577 9571
rect 15577 9537 15611 9571
rect 15611 9537 15620 9571
rect 15568 9528 15620 9537
rect 15936 9571 15988 9580
rect 15936 9537 15945 9571
rect 15945 9537 15979 9571
rect 15979 9537 15988 9571
rect 15936 9528 15988 9537
rect 16212 9571 16264 9580
rect 16212 9537 16221 9571
rect 16221 9537 16255 9571
rect 16255 9537 16264 9571
rect 16212 9528 16264 9537
rect 17592 9528 17644 9580
rect 17500 9460 17552 9512
rect 23020 9664 23072 9716
rect 24676 9664 24728 9716
rect 24952 9664 25004 9716
rect 28172 9664 28224 9716
rect 28448 9664 28500 9716
rect 29460 9707 29512 9716
rect 29460 9673 29469 9707
rect 29469 9673 29503 9707
rect 29503 9673 29512 9707
rect 29460 9664 29512 9673
rect 29552 9707 29604 9716
rect 29552 9673 29561 9707
rect 29561 9673 29595 9707
rect 29595 9673 29604 9707
rect 29552 9664 29604 9673
rect 23572 9596 23624 9648
rect 28356 9639 28408 9648
rect 21180 9528 21232 9580
rect 21732 9528 21784 9580
rect 18788 9460 18840 9512
rect 19156 9503 19208 9512
rect 19156 9469 19165 9503
rect 19165 9469 19199 9503
rect 19199 9469 19208 9503
rect 19156 9460 19208 9469
rect 19432 9460 19484 9512
rect 21088 9460 21140 9512
rect 23940 9528 23992 9580
rect 23480 9503 23532 9512
rect 23480 9469 23489 9503
rect 23489 9469 23523 9503
rect 23523 9469 23532 9503
rect 23480 9460 23532 9469
rect 25044 9528 25096 9580
rect 25412 9571 25464 9580
rect 25412 9537 25421 9571
rect 25421 9537 25455 9571
rect 25455 9537 25464 9571
rect 25412 9528 25464 9537
rect 25504 9528 25556 9580
rect 25872 9571 25924 9580
rect 25872 9537 25881 9571
rect 25881 9537 25915 9571
rect 25915 9537 25924 9571
rect 25872 9528 25924 9537
rect 25964 9528 26016 9580
rect 24308 9460 24360 9512
rect 26608 9460 26660 9512
rect 15200 9392 15252 9444
rect 16304 9392 16356 9444
rect 16488 9392 16540 9444
rect 15660 9324 15712 9376
rect 28356 9605 28365 9639
rect 28365 9605 28399 9639
rect 28399 9605 28408 9639
rect 28356 9596 28408 9605
rect 29736 9639 29788 9648
rect 29736 9605 29745 9639
rect 29745 9605 29779 9639
rect 29779 9605 29788 9639
rect 29736 9596 29788 9605
rect 31944 9664 31996 9716
rect 32128 9664 32180 9716
rect 32680 9664 32732 9716
rect 32956 9664 33008 9716
rect 33324 9707 33376 9716
rect 33324 9673 33339 9707
rect 33339 9673 33373 9707
rect 33373 9673 33376 9707
rect 33324 9664 33376 9673
rect 33692 9664 33744 9716
rect 38384 9664 38436 9716
rect 46664 9664 46716 9716
rect 31300 9596 31352 9648
rect 33968 9596 34020 9648
rect 39212 9596 39264 9648
rect 44272 9596 44324 9648
rect 45468 9639 45520 9648
rect 45468 9605 45502 9639
rect 45502 9605 45520 9639
rect 45468 9596 45520 9605
rect 27620 9528 27672 9580
rect 27528 9392 27580 9444
rect 21088 9324 21140 9376
rect 23020 9324 23072 9376
rect 23940 9324 23992 9376
rect 24768 9324 24820 9376
rect 28448 9571 28500 9580
rect 28448 9537 28457 9571
rect 28457 9537 28491 9571
rect 28491 9537 28500 9571
rect 28448 9528 28500 9537
rect 29276 9528 29328 9580
rect 28816 9460 28868 9512
rect 29092 9460 29144 9512
rect 30288 9528 30340 9580
rect 31024 9571 31076 9580
rect 31024 9537 31033 9571
rect 31033 9537 31067 9571
rect 31067 9537 31076 9571
rect 31024 9528 31076 9537
rect 31760 9528 31812 9580
rect 32680 9528 32732 9580
rect 33416 9571 33468 9580
rect 33140 9460 33192 9512
rect 33416 9537 33425 9571
rect 33425 9537 33459 9571
rect 33459 9537 33468 9571
rect 33416 9528 33468 9537
rect 33692 9528 33744 9580
rect 35992 9571 36044 9580
rect 35992 9537 36001 9571
rect 36001 9537 36035 9571
rect 36035 9537 36044 9571
rect 35992 9528 36044 9537
rect 36544 9528 36596 9580
rect 37464 9571 37516 9580
rect 37464 9537 37473 9571
rect 37473 9537 37507 9571
rect 37507 9537 37516 9571
rect 37464 9528 37516 9537
rect 33876 9460 33928 9512
rect 37832 9571 37884 9580
rect 37832 9537 37841 9571
rect 37841 9537 37875 9571
rect 37875 9537 37884 9571
rect 37832 9528 37884 9537
rect 38108 9528 38160 9580
rect 38568 9571 38620 9580
rect 38568 9537 38577 9571
rect 38577 9537 38611 9571
rect 38611 9537 38620 9571
rect 38568 9528 38620 9537
rect 38660 9571 38712 9580
rect 38660 9537 38670 9571
rect 38670 9537 38704 9571
rect 38704 9537 38712 9571
rect 38844 9571 38896 9580
rect 38660 9528 38712 9537
rect 38844 9537 38853 9571
rect 38853 9537 38887 9571
rect 38887 9537 38896 9571
rect 38844 9528 38896 9537
rect 40592 9528 40644 9580
rect 40776 9528 40828 9580
rect 42432 9528 42484 9580
rect 43996 9460 44048 9512
rect 44180 9571 44232 9580
rect 44180 9537 44189 9571
rect 44189 9537 44223 9571
rect 44223 9537 44232 9571
rect 45192 9571 45244 9580
rect 44180 9528 44232 9537
rect 45192 9537 45201 9571
rect 45201 9537 45235 9571
rect 45235 9537 45244 9571
rect 45192 9528 45244 9537
rect 46296 9528 46348 9580
rect 56968 9571 57020 9580
rect 56968 9537 56977 9571
rect 56977 9537 57011 9571
rect 57011 9537 57020 9571
rect 56968 9528 57020 9537
rect 57060 9528 57112 9580
rect 31668 9392 31720 9444
rect 34520 9392 34572 9444
rect 35164 9392 35216 9444
rect 29000 9324 29052 9376
rect 29828 9324 29880 9376
rect 31024 9324 31076 9376
rect 31576 9324 31628 9376
rect 32588 9324 32640 9376
rect 35900 9324 35952 9376
rect 36268 9324 36320 9376
rect 37556 9324 37608 9376
rect 38844 9392 38896 9444
rect 39304 9392 39356 9444
rect 44456 9392 44508 9444
rect 40316 9324 40368 9376
rect 56324 9324 56376 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 13820 9120 13872 9172
rect 13268 9095 13320 9104
rect 13268 9061 13277 9095
rect 13277 9061 13311 9095
rect 13311 9061 13320 9095
rect 13268 9052 13320 9061
rect 15200 9120 15252 9172
rect 16212 9120 16264 9172
rect 21088 9120 21140 9172
rect 21272 9163 21324 9172
rect 21272 9129 21281 9163
rect 21281 9129 21315 9163
rect 21315 9129 21324 9163
rect 21272 9120 21324 9129
rect 23664 9120 23716 9172
rect 27068 9120 27120 9172
rect 27988 9120 28040 9172
rect 10692 8984 10744 9036
rect 23572 9052 23624 9104
rect 24032 9052 24084 9104
rect 24400 9052 24452 9104
rect 13544 8984 13596 9036
rect 8300 8916 8352 8968
rect 14280 8916 14332 8968
rect 17592 8984 17644 9036
rect 1860 8891 1912 8900
rect 1860 8857 1869 8891
rect 1869 8857 1903 8891
rect 1903 8857 1912 8891
rect 1860 8848 1912 8857
rect 12440 8848 12492 8900
rect 13636 8848 13688 8900
rect 14924 8891 14976 8900
rect 14924 8857 14933 8891
rect 14933 8857 14967 8891
rect 14967 8857 14976 8891
rect 14924 8848 14976 8857
rect 17040 8916 17092 8968
rect 17500 8891 17552 8900
rect 13452 8780 13504 8832
rect 15108 8823 15160 8832
rect 15108 8789 15117 8823
rect 15117 8789 15151 8823
rect 15151 8789 15160 8823
rect 17500 8857 17509 8891
rect 17509 8857 17543 8891
rect 17543 8857 17552 8891
rect 17500 8848 17552 8857
rect 18052 8925 18061 8934
rect 18061 8925 18095 8934
rect 18095 8925 18104 8934
rect 18052 8882 18104 8925
rect 18788 8984 18840 9036
rect 25872 9052 25924 9104
rect 28172 9052 28224 9104
rect 30288 9120 30340 9172
rect 29736 9052 29788 9104
rect 30656 9052 30708 9104
rect 21548 8848 21600 8900
rect 22468 8916 22520 8968
rect 23664 8959 23716 8968
rect 23664 8925 23673 8959
rect 23673 8925 23707 8959
rect 23707 8925 23716 8959
rect 23664 8916 23716 8925
rect 23388 8848 23440 8900
rect 15108 8780 15160 8789
rect 18788 8780 18840 8832
rect 19064 8780 19116 8832
rect 21180 8780 21232 8832
rect 23020 8780 23072 8832
rect 24124 8916 24176 8968
rect 24032 8891 24084 8900
rect 24032 8857 24041 8891
rect 24041 8857 24075 8891
rect 24075 8857 24084 8891
rect 24032 8848 24084 8857
rect 25964 8984 26016 9036
rect 25320 8916 25372 8968
rect 25688 8959 25740 8968
rect 25688 8925 25697 8959
rect 25697 8925 25731 8959
rect 25731 8925 25740 8959
rect 25688 8916 25740 8925
rect 25780 8916 25832 8968
rect 27436 8984 27488 9036
rect 27896 9027 27948 9036
rect 27896 8993 27905 9027
rect 27905 8993 27939 9027
rect 27939 8993 27948 9027
rect 27896 8984 27948 8993
rect 29184 8984 29236 9036
rect 30104 8984 30156 9036
rect 32496 9120 32548 9172
rect 33692 9120 33744 9172
rect 34152 9120 34204 9172
rect 35992 9120 36044 9172
rect 38936 9120 38988 9172
rect 31392 9095 31444 9104
rect 31392 9061 31401 9095
rect 31401 9061 31435 9095
rect 31435 9061 31444 9095
rect 31392 9052 31444 9061
rect 32588 9052 32640 9104
rect 33140 9052 33192 9104
rect 26424 8959 26476 8968
rect 26424 8925 26433 8959
rect 26433 8925 26467 8959
rect 26467 8925 26476 8959
rect 26424 8916 26476 8925
rect 27804 8959 27856 8968
rect 26332 8848 26384 8900
rect 23848 8823 23900 8832
rect 23848 8789 23857 8823
rect 23857 8789 23891 8823
rect 23891 8789 23900 8823
rect 23848 8780 23900 8789
rect 24952 8780 25004 8832
rect 26516 8780 26568 8832
rect 26976 8780 27028 8832
rect 27436 8848 27488 8900
rect 27804 8925 27813 8959
rect 27813 8925 27847 8959
rect 27847 8925 27856 8959
rect 27804 8916 27856 8925
rect 27988 8916 28040 8968
rect 31484 8916 31536 8968
rect 31576 8959 31628 8968
rect 31576 8925 31585 8959
rect 31585 8925 31619 8959
rect 31619 8925 31628 8959
rect 31576 8916 31628 8925
rect 32220 8916 32272 8968
rect 33140 8959 33192 8968
rect 33140 8925 33149 8959
rect 33149 8925 33183 8959
rect 33183 8925 33192 8959
rect 33140 8916 33192 8925
rect 34428 8984 34480 9036
rect 36452 9052 36504 9104
rect 36268 9027 36320 9036
rect 36268 8993 36277 9027
rect 36277 8993 36311 9027
rect 36311 8993 36320 9027
rect 36268 8984 36320 8993
rect 37188 8984 37240 9036
rect 28448 8848 28500 8900
rect 29092 8848 29144 8900
rect 30104 8848 30156 8900
rect 31944 8891 31996 8900
rect 27988 8780 28040 8832
rect 29736 8780 29788 8832
rect 30012 8780 30064 8832
rect 31392 8780 31444 8832
rect 31668 8823 31720 8832
rect 31668 8789 31677 8823
rect 31677 8789 31711 8823
rect 31711 8789 31720 8823
rect 31668 8780 31720 8789
rect 31944 8857 31953 8891
rect 31953 8857 31987 8891
rect 31987 8857 31996 8891
rect 31944 8848 31996 8857
rect 34244 8916 34296 8968
rect 35900 8916 35952 8968
rect 37096 8916 37148 8968
rect 37740 8959 37792 8968
rect 37740 8925 37749 8959
rect 37749 8925 37783 8959
rect 37783 8925 37792 8959
rect 37740 8916 37792 8925
rect 38568 8984 38620 9036
rect 39304 8984 39356 9036
rect 33692 8848 33744 8900
rect 37464 8848 37516 8900
rect 38476 8916 38528 8968
rect 41328 9120 41380 9172
rect 46756 9120 46808 9172
rect 40040 9095 40092 9104
rect 40040 9061 40049 9095
rect 40049 9061 40083 9095
rect 40083 9061 40092 9095
rect 40040 9052 40092 9061
rect 41788 9052 41840 9104
rect 40224 8916 40276 8968
rect 44088 8984 44140 9036
rect 44456 9027 44508 9036
rect 44456 8993 44465 9027
rect 44465 8993 44499 9027
rect 44499 8993 44508 9027
rect 44456 8984 44508 8993
rect 45008 8984 45060 9036
rect 46204 8984 46256 9036
rect 40868 8916 40920 8968
rect 45100 8916 45152 8968
rect 46112 8959 46164 8968
rect 46112 8925 46121 8959
rect 46121 8925 46155 8959
rect 46155 8925 46164 8959
rect 46112 8916 46164 8925
rect 46296 8959 46348 8968
rect 46296 8925 46305 8959
rect 46305 8925 46339 8959
rect 46339 8925 46348 8959
rect 46296 8916 46348 8925
rect 46848 8916 46900 8968
rect 56876 9027 56928 9036
rect 56140 8959 56192 8968
rect 56140 8925 56149 8959
rect 56149 8925 56183 8959
rect 56183 8925 56192 8959
rect 56140 8916 56192 8925
rect 56324 8959 56376 8968
rect 56324 8925 56333 8959
rect 56333 8925 56367 8959
rect 56367 8925 56376 8959
rect 56324 8916 56376 8925
rect 56876 8993 56885 9027
rect 56885 8993 56919 9027
rect 56919 8993 56928 9027
rect 56876 8984 56928 8993
rect 38016 8891 38068 8900
rect 38016 8857 38025 8891
rect 38025 8857 38059 8891
rect 38059 8857 38068 8891
rect 38016 8848 38068 8857
rect 32588 8780 32640 8832
rect 33140 8780 33192 8832
rect 35992 8823 36044 8832
rect 35992 8789 36001 8823
rect 36001 8789 36035 8823
rect 36035 8789 36044 8823
rect 35992 8780 36044 8789
rect 37280 8780 37332 8832
rect 41236 8848 41288 8900
rect 41328 8848 41380 8900
rect 43444 8848 43496 8900
rect 43720 8891 43772 8900
rect 43720 8857 43729 8891
rect 43729 8857 43763 8891
rect 43763 8857 43772 8891
rect 43720 8848 43772 8857
rect 44088 8848 44140 8900
rect 38384 8823 38436 8832
rect 38384 8789 38393 8823
rect 38393 8789 38427 8823
rect 38427 8789 38436 8823
rect 38384 8780 38436 8789
rect 40960 8780 41012 8832
rect 57060 8780 57112 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 13452 8576 13504 8628
rect 14924 8576 14976 8628
rect 16580 8576 16632 8628
rect 17224 8576 17276 8628
rect 15108 8508 15160 8560
rect 17040 8551 17092 8560
rect 10600 8440 10652 8492
rect 14004 8483 14056 8492
rect 14004 8449 14013 8483
rect 14013 8449 14047 8483
rect 14047 8449 14056 8483
rect 14004 8440 14056 8449
rect 15292 8440 15344 8492
rect 17040 8517 17049 8551
rect 17049 8517 17083 8551
rect 17083 8517 17092 8551
rect 17040 8508 17092 8517
rect 19156 8576 19208 8628
rect 19248 8576 19300 8628
rect 19892 8576 19944 8628
rect 22744 8576 22796 8628
rect 15476 8440 15528 8492
rect 16672 8440 16724 8492
rect 17132 8440 17184 8492
rect 17960 8508 18012 8560
rect 23296 8576 23348 8628
rect 23848 8576 23900 8628
rect 25136 8576 25188 8628
rect 28356 8576 28408 8628
rect 28724 8576 28776 8628
rect 31576 8576 31628 8628
rect 34244 8576 34296 8628
rect 1768 8415 1820 8424
rect 1768 8381 1777 8415
rect 1777 8381 1811 8415
rect 1811 8381 1820 8415
rect 1768 8372 1820 8381
rect 17316 8372 17368 8424
rect 17868 8440 17920 8492
rect 29552 8508 29604 8560
rect 20352 8440 20404 8492
rect 22376 8483 22428 8492
rect 22376 8449 22385 8483
rect 22385 8449 22419 8483
rect 22419 8449 22428 8483
rect 22376 8440 22428 8449
rect 24124 8483 24176 8492
rect 19984 8372 20036 8424
rect 22284 8372 22336 8424
rect 13360 8304 13412 8356
rect 15660 8236 15712 8288
rect 17408 8236 17460 8288
rect 17868 8304 17920 8356
rect 18972 8304 19024 8356
rect 19892 8304 19944 8356
rect 20260 8304 20312 8356
rect 24124 8449 24133 8483
rect 24133 8449 24167 8483
rect 24167 8449 24176 8483
rect 24124 8440 24176 8449
rect 27160 8483 27212 8492
rect 27160 8449 27169 8483
rect 27169 8449 27203 8483
rect 27203 8449 27212 8483
rect 27160 8440 27212 8449
rect 27528 8440 27580 8492
rect 29000 8440 29052 8492
rect 29460 8483 29512 8492
rect 29460 8449 29469 8483
rect 29469 8449 29503 8483
rect 29503 8449 29512 8483
rect 29460 8440 29512 8449
rect 23940 8372 23992 8424
rect 25412 8372 25464 8424
rect 25780 8372 25832 8424
rect 27712 8372 27764 8424
rect 28540 8372 28592 8424
rect 31024 8508 31076 8560
rect 33508 8508 33560 8560
rect 29736 8372 29788 8424
rect 24492 8304 24544 8356
rect 30196 8440 30248 8492
rect 30656 8440 30708 8492
rect 32772 8483 32824 8492
rect 32772 8449 32781 8483
rect 32781 8449 32815 8483
rect 32815 8449 32824 8483
rect 32772 8440 32824 8449
rect 33140 8483 33192 8492
rect 30104 8415 30156 8424
rect 30104 8381 30113 8415
rect 30113 8381 30147 8415
rect 30147 8381 30156 8415
rect 31300 8415 31352 8424
rect 30104 8372 30156 8381
rect 31300 8381 31309 8415
rect 31309 8381 31343 8415
rect 31343 8381 31352 8415
rect 31300 8372 31352 8381
rect 31760 8372 31812 8424
rect 33140 8449 33149 8483
rect 33149 8449 33183 8483
rect 33183 8449 33192 8483
rect 33140 8440 33192 8449
rect 33692 8440 33744 8492
rect 33876 8483 33928 8492
rect 33876 8449 33885 8483
rect 33885 8449 33919 8483
rect 33919 8449 33928 8483
rect 33876 8440 33928 8449
rect 30196 8304 30248 8356
rect 30472 8304 30524 8356
rect 31208 8347 31260 8356
rect 31208 8313 31217 8347
rect 31217 8313 31251 8347
rect 31251 8313 31260 8347
rect 31208 8304 31260 8313
rect 33416 8304 33468 8356
rect 35348 8576 35400 8628
rect 40960 8576 41012 8628
rect 46112 8576 46164 8628
rect 46204 8576 46256 8628
rect 18512 8236 18564 8288
rect 19064 8236 19116 8288
rect 19248 8236 19300 8288
rect 20812 8236 20864 8288
rect 23020 8236 23072 8288
rect 23572 8236 23624 8288
rect 27620 8236 27672 8288
rect 29092 8236 29144 8288
rect 31300 8236 31352 8288
rect 33968 8236 34020 8288
rect 34428 8440 34480 8492
rect 35900 8483 35952 8492
rect 35900 8449 35909 8483
rect 35909 8449 35943 8483
rect 35943 8449 35952 8483
rect 35900 8440 35952 8449
rect 36728 8483 36780 8492
rect 36728 8449 36737 8483
rect 36737 8449 36771 8483
rect 36771 8449 36780 8483
rect 36728 8440 36780 8449
rect 35808 8415 35860 8424
rect 35808 8381 35817 8415
rect 35817 8381 35851 8415
rect 35851 8381 35860 8415
rect 35808 8372 35860 8381
rect 37280 8440 37332 8492
rect 37648 8508 37700 8560
rect 37556 8483 37608 8492
rect 37556 8449 37565 8483
rect 37565 8449 37599 8483
rect 37599 8449 37608 8483
rect 37556 8440 37608 8449
rect 37096 8372 37148 8424
rect 39948 8508 40000 8560
rect 45192 8508 45244 8560
rect 39212 8440 39264 8492
rect 42984 8440 43036 8492
rect 44272 8440 44324 8492
rect 44548 8483 44600 8492
rect 44548 8449 44557 8483
rect 44557 8449 44591 8483
rect 44591 8449 44600 8483
rect 44548 8440 44600 8449
rect 38016 8372 38068 8424
rect 39120 8415 39172 8424
rect 39120 8381 39129 8415
rect 39129 8381 39163 8415
rect 39163 8381 39172 8415
rect 39120 8372 39172 8381
rect 42524 8372 42576 8424
rect 43904 8372 43956 8424
rect 44824 8483 44876 8492
rect 44824 8449 44833 8483
rect 44833 8449 44867 8483
rect 44867 8449 44876 8483
rect 53104 8508 53156 8560
rect 57336 8551 57388 8560
rect 57336 8517 57345 8551
rect 57345 8517 57379 8551
rect 57379 8517 57388 8551
rect 57336 8508 57388 8517
rect 44824 8440 44876 8449
rect 46388 8483 46440 8492
rect 46388 8449 46397 8483
rect 46397 8449 46431 8483
rect 46431 8449 46440 8483
rect 46388 8440 46440 8449
rect 56232 8483 56284 8492
rect 56232 8449 56241 8483
rect 56241 8449 56275 8483
rect 56275 8449 56284 8483
rect 56232 8440 56284 8449
rect 57060 8483 57112 8492
rect 57060 8449 57069 8483
rect 57069 8449 57103 8483
rect 57103 8449 57112 8483
rect 57060 8440 57112 8449
rect 45376 8372 45428 8424
rect 45468 8415 45520 8424
rect 45468 8381 45477 8415
rect 45477 8381 45511 8415
rect 45511 8381 45520 8415
rect 46572 8415 46624 8424
rect 45468 8372 45520 8381
rect 46572 8381 46581 8415
rect 46581 8381 46615 8415
rect 46615 8381 46624 8415
rect 46572 8372 46624 8381
rect 34428 8236 34480 8288
rect 40868 8304 40920 8356
rect 56508 8304 56560 8356
rect 36912 8279 36964 8288
rect 36912 8245 36921 8279
rect 36921 8245 36955 8279
rect 36955 8245 36964 8279
rect 36912 8236 36964 8245
rect 38844 8236 38896 8288
rect 43168 8236 43220 8288
rect 43444 8236 43496 8288
rect 44824 8236 44876 8288
rect 45468 8236 45520 8288
rect 55496 8236 55548 8288
rect 56968 8236 57020 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 2688 8032 2740 8084
rect 10048 8032 10100 8084
rect 26240 8032 26292 8084
rect 12716 7964 12768 8016
rect 14004 7964 14056 8016
rect 15200 7964 15252 8016
rect 16488 7964 16540 8016
rect 16672 7964 16724 8016
rect 17500 7964 17552 8016
rect 17592 7964 17644 8016
rect 17776 7964 17828 8016
rect 18696 7964 18748 8016
rect 19156 7964 19208 8016
rect 20812 8007 20864 8016
rect 20812 7973 20821 8007
rect 20821 7973 20855 8007
rect 20855 7973 20864 8007
rect 20812 7964 20864 7973
rect 1584 7871 1636 7880
rect 1584 7837 1593 7871
rect 1593 7837 1627 7871
rect 1627 7837 1636 7871
rect 1584 7828 1636 7837
rect 6000 7828 6052 7880
rect 7932 7871 7984 7880
rect 7932 7837 7941 7871
rect 7941 7837 7975 7871
rect 7975 7837 7984 7871
rect 7932 7828 7984 7837
rect 8760 7828 8812 7880
rect 10048 7828 10100 7880
rect 16304 7896 16356 7948
rect 15016 7828 15068 7880
rect 15200 7871 15252 7880
rect 15200 7837 15209 7871
rect 15209 7837 15243 7871
rect 15243 7837 15252 7871
rect 15200 7828 15252 7837
rect 15476 7871 15528 7880
rect 15476 7837 15485 7871
rect 15485 7837 15519 7871
rect 15519 7837 15528 7871
rect 15476 7828 15528 7837
rect 16028 7828 16080 7880
rect 17316 7896 17368 7948
rect 19432 7939 19484 7948
rect 19432 7905 19441 7939
rect 19441 7905 19475 7939
rect 19475 7905 19484 7939
rect 19432 7896 19484 7905
rect 20720 7896 20772 7948
rect 23756 7896 23808 7948
rect 32404 8032 32456 8084
rect 33968 8032 34020 8084
rect 35808 8032 35860 8084
rect 27344 7964 27396 8016
rect 30472 7964 30524 8016
rect 30932 8007 30984 8016
rect 30932 7973 30941 8007
rect 30941 7973 30975 8007
rect 30975 7973 30984 8007
rect 30932 7964 30984 7973
rect 31300 7964 31352 8016
rect 31668 7964 31720 8016
rect 31852 7964 31904 8016
rect 32496 7964 32548 8016
rect 33140 7964 33192 8016
rect 33324 7964 33376 8016
rect 34612 7964 34664 8016
rect 35624 7964 35676 8016
rect 35716 7964 35768 8016
rect 37740 8032 37792 8084
rect 39212 8032 39264 8084
rect 43720 8032 43772 8084
rect 46388 8032 46440 8084
rect 37280 7964 37332 8016
rect 38844 7964 38896 8016
rect 38936 8007 38988 8016
rect 38936 7973 38945 8007
rect 38945 7973 38979 8007
rect 38979 7973 38988 8007
rect 38936 7964 38988 7973
rect 43168 7964 43220 8016
rect 55956 7964 56008 8016
rect 28724 7939 28776 7948
rect 28724 7905 28733 7939
rect 28733 7905 28767 7939
rect 28767 7905 28776 7939
rect 28724 7896 28776 7905
rect 29828 7939 29880 7948
rect 29828 7905 29837 7939
rect 29837 7905 29871 7939
rect 29871 7905 29880 7939
rect 29828 7896 29880 7905
rect 17224 7871 17276 7880
rect 17224 7837 17233 7871
rect 17233 7837 17267 7871
rect 17267 7837 17276 7871
rect 17224 7828 17276 7837
rect 17408 7828 17460 7880
rect 17960 7871 18012 7880
rect 17960 7837 17969 7871
rect 17969 7837 18003 7871
rect 18003 7837 18012 7871
rect 17960 7828 18012 7837
rect 19064 7828 19116 7880
rect 1860 7803 1912 7812
rect 1860 7769 1869 7803
rect 1869 7769 1903 7803
rect 1903 7769 1912 7803
rect 1860 7760 1912 7769
rect 8576 7803 8628 7812
rect 8576 7769 8585 7803
rect 8585 7769 8619 7803
rect 8619 7769 8628 7803
rect 8576 7760 8628 7769
rect 9772 7803 9824 7812
rect 9772 7769 9781 7803
rect 9781 7769 9815 7803
rect 9815 7769 9824 7803
rect 9772 7760 9824 7769
rect 12440 7760 12492 7812
rect 15752 7760 15804 7812
rect 19984 7828 20036 7880
rect 24032 7828 24084 7880
rect 24952 7871 25004 7880
rect 24952 7837 24961 7871
rect 24961 7837 24995 7871
rect 24995 7837 25004 7871
rect 24952 7828 25004 7837
rect 28264 7828 28316 7880
rect 29460 7828 29512 7880
rect 30012 7871 30064 7880
rect 30012 7837 30021 7871
rect 30021 7837 30055 7871
rect 30055 7837 30064 7871
rect 30012 7828 30064 7837
rect 31024 7828 31076 7880
rect 9956 7692 10008 7744
rect 15292 7692 15344 7744
rect 16028 7692 16080 7744
rect 16764 7692 16816 7744
rect 17960 7692 18012 7744
rect 18512 7692 18564 7744
rect 19340 7692 19392 7744
rect 28724 7760 28776 7812
rect 31208 7760 31260 7812
rect 32220 7828 32272 7880
rect 20168 7692 20220 7744
rect 20352 7692 20404 7744
rect 21456 7692 21508 7744
rect 22284 7692 22336 7744
rect 23020 7735 23072 7744
rect 23020 7701 23029 7735
rect 23029 7701 23063 7735
rect 23063 7701 23072 7735
rect 23020 7692 23072 7701
rect 23112 7735 23164 7744
rect 23112 7701 23121 7735
rect 23121 7701 23155 7735
rect 23155 7701 23164 7735
rect 23112 7692 23164 7701
rect 23480 7692 23532 7744
rect 31116 7692 31168 7744
rect 31852 7735 31904 7744
rect 31852 7701 31861 7735
rect 31861 7701 31895 7735
rect 31895 7701 31904 7735
rect 31852 7692 31904 7701
rect 33600 7828 33652 7880
rect 34152 7871 34204 7880
rect 34152 7837 34161 7871
rect 34161 7837 34195 7871
rect 34195 7837 34204 7871
rect 34152 7828 34204 7837
rect 33140 7803 33192 7812
rect 33140 7769 33149 7803
rect 33149 7769 33183 7803
rect 33183 7769 33192 7803
rect 33140 7760 33192 7769
rect 35164 7828 35216 7880
rect 34704 7760 34756 7812
rect 38384 7896 38436 7948
rect 38660 7896 38712 7948
rect 39396 7896 39448 7948
rect 39672 7896 39724 7948
rect 36912 7828 36964 7880
rect 38660 7760 38712 7812
rect 38835 7837 38862 7846
rect 38862 7837 38887 7846
rect 38835 7794 38887 7837
rect 39212 7828 39264 7880
rect 40040 7828 40092 7880
rect 42524 7828 42576 7880
rect 43444 7828 43496 7880
rect 43996 7871 44048 7880
rect 43996 7837 44005 7871
rect 44005 7837 44039 7871
rect 44039 7837 44048 7871
rect 43996 7828 44048 7837
rect 44180 7828 44232 7880
rect 45284 7871 45336 7880
rect 45284 7837 45293 7871
rect 45293 7837 45327 7871
rect 45327 7837 45336 7871
rect 45284 7828 45336 7837
rect 45376 7828 45428 7880
rect 46572 7896 46624 7948
rect 46664 7939 46716 7948
rect 46664 7905 46673 7939
rect 46673 7905 46707 7939
rect 46707 7905 46716 7939
rect 57796 8032 57848 8084
rect 56876 7939 56928 7948
rect 46664 7896 46716 7905
rect 55496 7871 55548 7880
rect 55496 7837 55505 7871
rect 55505 7837 55539 7871
rect 55539 7837 55548 7871
rect 55496 7828 55548 7837
rect 55772 7828 55824 7880
rect 56876 7905 56885 7939
rect 56885 7905 56919 7939
rect 56919 7905 56928 7939
rect 56876 7896 56928 7905
rect 43904 7803 43956 7812
rect 43904 7769 43913 7803
rect 43913 7769 43947 7803
rect 43947 7769 43956 7803
rect 43904 7760 43956 7769
rect 44456 7803 44508 7812
rect 44456 7769 44465 7803
rect 44465 7769 44499 7803
rect 44499 7769 44508 7803
rect 44456 7760 44508 7769
rect 46756 7760 46808 7812
rect 56140 7803 56192 7812
rect 56140 7769 56149 7803
rect 56149 7769 56183 7803
rect 56183 7769 56192 7803
rect 56140 7760 56192 7769
rect 33048 7692 33100 7744
rect 34152 7692 34204 7744
rect 36544 7692 36596 7744
rect 37740 7692 37792 7744
rect 39672 7692 39724 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 10600 7531 10652 7540
rect 10600 7497 10609 7531
rect 10609 7497 10643 7531
rect 10643 7497 10652 7531
rect 10600 7488 10652 7497
rect 15016 7488 15068 7540
rect 16764 7488 16816 7540
rect 1584 7420 1636 7472
rect 10784 7420 10836 7472
rect 15476 7420 15528 7472
rect 15660 7420 15712 7472
rect 9496 7395 9548 7404
rect 9496 7361 9505 7395
rect 9505 7361 9539 7395
rect 9539 7361 9548 7395
rect 9496 7352 9548 7361
rect 9588 7352 9640 7404
rect 11428 7352 11480 7404
rect 15752 7395 15804 7404
rect 15752 7361 15761 7395
rect 15761 7361 15795 7395
rect 15795 7361 15804 7395
rect 15752 7352 15804 7361
rect 16304 7420 16356 7472
rect 17224 7420 17276 7472
rect 17500 7463 17552 7472
rect 17500 7429 17509 7463
rect 17509 7429 17543 7463
rect 17543 7429 17552 7463
rect 17500 7420 17552 7429
rect 16028 7352 16080 7404
rect 17132 7352 17184 7404
rect 18052 7488 18104 7540
rect 21456 7488 21508 7540
rect 23480 7531 23532 7540
rect 17868 7420 17920 7472
rect 19064 7463 19116 7472
rect 19064 7429 19073 7463
rect 19073 7429 19107 7463
rect 19107 7429 19116 7463
rect 19064 7420 19116 7429
rect 19524 7420 19576 7472
rect 18972 7395 19024 7404
rect 18972 7361 18981 7395
rect 18981 7361 19015 7395
rect 19015 7361 19024 7395
rect 18972 7352 19024 7361
rect 19432 7352 19484 7404
rect 21180 7352 21232 7404
rect 10692 7284 10744 7336
rect 10876 7327 10928 7336
rect 10876 7293 10885 7327
rect 10885 7293 10919 7327
rect 10919 7293 10928 7327
rect 10876 7284 10928 7293
rect 11060 7327 11112 7336
rect 11060 7293 11069 7327
rect 11069 7293 11103 7327
rect 11103 7293 11112 7327
rect 12440 7327 12492 7336
rect 11060 7284 11112 7293
rect 12440 7293 12449 7327
rect 12449 7293 12483 7327
rect 12483 7293 12492 7327
rect 12440 7284 12492 7293
rect 16304 7327 16356 7336
rect 7380 7216 7432 7268
rect 15200 7216 15252 7268
rect 9404 7148 9456 7200
rect 16304 7293 16313 7327
rect 16313 7293 16347 7327
rect 16347 7293 16356 7327
rect 16304 7284 16356 7293
rect 17040 7327 17092 7336
rect 17040 7293 17049 7327
rect 17049 7293 17083 7327
rect 17083 7293 17092 7327
rect 17040 7284 17092 7293
rect 17868 7284 17920 7336
rect 19064 7284 19116 7336
rect 19892 7284 19944 7336
rect 23480 7497 23489 7531
rect 23489 7497 23523 7531
rect 23523 7497 23532 7531
rect 23480 7488 23532 7497
rect 27804 7488 27856 7540
rect 29276 7488 29328 7540
rect 29920 7531 29972 7540
rect 29920 7497 29929 7531
rect 29929 7497 29963 7531
rect 29963 7497 29972 7531
rect 29920 7488 29972 7497
rect 30196 7488 30248 7540
rect 30472 7488 30524 7540
rect 31576 7488 31628 7540
rect 35440 7531 35492 7540
rect 27344 7420 27396 7472
rect 27620 7420 27672 7472
rect 28172 7420 28224 7472
rect 17316 7216 17368 7268
rect 18052 7216 18104 7268
rect 19156 7216 19208 7268
rect 19984 7216 20036 7268
rect 21088 7216 21140 7268
rect 21272 7148 21324 7200
rect 21456 7191 21508 7200
rect 21456 7157 21465 7191
rect 21465 7157 21499 7191
rect 21499 7157 21508 7191
rect 21456 7148 21508 7157
rect 21548 7148 21600 7200
rect 25688 7148 25740 7200
rect 27528 7395 27580 7404
rect 27528 7361 27537 7395
rect 27537 7361 27571 7395
rect 27571 7361 27580 7395
rect 27528 7352 27580 7361
rect 28632 7395 28684 7404
rect 28632 7361 28641 7395
rect 28641 7361 28675 7395
rect 28675 7361 28684 7395
rect 28632 7352 28684 7361
rect 32588 7395 32640 7404
rect 32588 7361 32597 7395
rect 32597 7361 32631 7395
rect 32631 7361 32640 7395
rect 32588 7352 32640 7361
rect 32772 7395 32824 7404
rect 32772 7361 32781 7395
rect 32781 7361 32815 7395
rect 32815 7361 32824 7395
rect 32772 7352 32824 7361
rect 33232 7352 33284 7404
rect 35164 7420 35216 7472
rect 35440 7497 35449 7531
rect 35449 7497 35483 7531
rect 35483 7497 35492 7531
rect 35440 7488 35492 7497
rect 36728 7488 36780 7540
rect 38568 7488 38620 7540
rect 44456 7488 44508 7540
rect 52460 7488 52512 7540
rect 56508 7488 56560 7540
rect 35348 7420 35400 7472
rect 35992 7420 36044 7472
rect 55772 7420 55824 7472
rect 34336 7395 34388 7404
rect 34336 7361 34370 7395
rect 34370 7361 34388 7395
rect 34336 7352 34388 7361
rect 34704 7352 34756 7404
rect 35716 7352 35768 7404
rect 36544 7395 36596 7404
rect 36544 7361 36553 7395
rect 36553 7361 36587 7395
rect 36587 7361 36596 7395
rect 36544 7352 36596 7361
rect 36912 7352 36964 7404
rect 43904 7352 43956 7404
rect 29092 7284 29144 7336
rect 30012 7284 30064 7336
rect 28264 7216 28316 7268
rect 30380 7216 30432 7268
rect 33140 7284 33192 7336
rect 35348 7284 35400 7336
rect 38568 7284 38620 7336
rect 40132 7284 40184 7336
rect 43168 7284 43220 7336
rect 32220 7216 32272 7268
rect 33876 7216 33928 7268
rect 30564 7148 30616 7200
rect 37280 7216 37332 7268
rect 35992 7148 36044 7200
rect 36912 7148 36964 7200
rect 44548 7352 44600 7404
rect 45100 7352 45152 7404
rect 45836 7352 45888 7404
rect 55956 7395 56008 7404
rect 55956 7361 55965 7395
rect 55965 7361 55999 7395
rect 55999 7361 56008 7395
rect 55956 7352 56008 7361
rect 56508 7395 56560 7404
rect 56508 7361 56517 7395
rect 56517 7361 56551 7395
rect 56551 7361 56560 7395
rect 56508 7352 56560 7361
rect 56968 7352 57020 7404
rect 58256 7395 58308 7404
rect 58256 7361 58265 7395
rect 58265 7361 58299 7395
rect 58299 7361 58308 7395
rect 58256 7352 58308 7361
rect 56140 7284 56192 7336
rect 45928 7148 45980 7200
rect 46388 7191 46440 7200
rect 46388 7157 46397 7191
rect 46397 7157 46431 7191
rect 46431 7157 46440 7191
rect 46388 7148 46440 7157
rect 56968 7148 57020 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 10876 6944 10928 6996
rect 20536 6944 20588 6996
rect 21180 6987 21232 6996
rect 21180 6953 21189 6987
rect 21189 6953 21223 6987
rect 21223 6953 21232 6987
rect 21180 6944 21232 6953
rect 21272 6944 21324 6996
rect 27160 6944 27212 6996
rect 27712 6944 27764 6996
rect 27896 6944 27948 6996
rect 31852 6944 31904 6996
rect 34336 6987 34388 6996
rect 18144 6876 18196 6928
rect 20720 6876 20772 6928
rect 23848 6919 23900 6928
rect 23848 6885 23857 6919
rect 23857 6885 23891 6919
rect 23891 6885 23900 6919
rect 23848 6876 23900 6885
rect 30840 6919 30892 6928
rect 8760 6808 8812 6860
rect 10784 6851 10836 6860
rect 9128 6740 9180 6792
rect 10784 6817 10793 6851
rect 10793 6817 10827 6851
rect 10827 6817 10836 6851
rect 10784 6808 10836 6817
rect 10876 6808 10928 6860
rect 18604 6808 18656 6860
rect 9588 6783 9640 6792
rect 9588 6749 9597 6783
rect 9597 6749 9631 6783
rect 9631 6749 9640 6783
rect 9588 6740 9640 6749
rect 10692 6740 10744 6792
rect 1860 6715 1912 6724
rect 1860 6681 1869 6715
rect 1869 6681 1903 6715
rect 1903 6681 1912 6715
rect 1860 6672 1912 6681
rect 9496 6604 9548 6656
rect 9680 6604 9732 6656
rect 11244 6783 11296 6792
rect 11244 6749 11253 6783
rect 11253 6749 11287 6783
rect 11287 6749 11296 6783
rect 11244 6740 11296 6749
rect 17408 6740 17460 6792
rect 17776 6740 17828 6792
rect 17960 6740 18012 6792
rect 18512 6740 18564 6792
rect 18972 6808 19024 6860
rect 21180 6808 21232 6860
rect 21732 6851 21784 6860
rect 21732 6817 21741 6851
rect 21741 6817 21775 6851
rect 21775 6817 21784 6851
rect 21732 6808 21784 6817
rect 26792 6808 26844 6860
rect 27068 6808 27120 6860
rect 11428 6672 11480 6724
rect 17500 6672 17552 6724
rect 19340 6740 19392 6792
rect 19616 6740 19668 6792
rect 24676 6783 24728 6792
rect 24676 6749 24685 6783
rect 24685 6749 24719 6783
rect 24719 6749 24728 6783
rect 24676 6740 24728 6749
rect 30840 6885 30849 6919
rect 30849 6885 30883 6919
rect 30883 6885 30892 6919
rect 30840 6876 30892 6885
rect 31576 6876 31628 6928
rect 34336 6953 34345 6987
rect 34345 6953 34379 6987
rect 34379 6953 34388 6987
rect 34336 6944 34388 6953
rect 27712 6808 27764 6860
rect 28080 6808 28132 6860
rect 28540 6851 28592 6860
rect 28540 6817 28549 6851
rect 28549 6817 28583 6851
rect 28583 6817 28592 6851
rect 28540 6808 28592 6817
rect 29828 6808 29880 6860
rect 31024 6808 31076 6860
rect 31668 6808 31720 6860
rect 33140 6808 33192 6860
rect 21180 6672 21232 6724
rect 16212 6604 16264 6656
rect 18144 6647 18196 6656
rect 18144 6613 18153 6647
rect 18153 6613 18187 6647
rect 18187 6613 18196 6647
rect 18144 6604 18196 6613
rect 18512 6647 18564 6656
rect 18512 6613 18521 6647
rect 18521 6613 18555 6647
rect 18555 6613 18564 6647
rect 18512 6604 18564 6613
rect 18604 6647 18656 6656
rect 18604 6613 18613 6647
rect 18613 6613 18647 6647
rect 18647 6613 18656 6647
rect 18604 6604 18656 6613
rect 20720 6604 20772 6656
rect 21456 6604 21508 6656
rect 22284 6672 22336 6724
rect 23296 6672 23348 6724
rect 24768 6672 24820 6724
rect 25596 6672 25648 6724
rect 26424 6672 26476 6724
rect 27988 6740 28040 6792
rect 28172 6783 28224 6792
rect 28172 6749 28181 6783
rect 28181 6749 28215 6783
rect 28215 6749 28224 6783
rect 28172 6740 28224 6749
rect 27804 6672 27856 6724
rect 22928 6604 22980 6656
rect 25136 6604 25188 6656
rect 26516 6604 26568 6656
rect 31484 6740 31536 6792
rect 31576 6740 31628 6792
rect 32680 6740 32732 6792
rect 30380 6672 30432 6724
rect 30288 6604 30340 6656
rect 32956 6783 33008 6792
rect 32956 6749 32965 6783
rect 32965 6749 32999 6783
rect 32999 6749 33008 6783
rect 32956 6740 33008 6749
rect 33692 6740 33744 6792
rect 34428 6808 34480 6860
rect 35348 6808 35400 6860
rect 45284 6944 45336 6996
rect 45836 6987 45888 6996
rect 45836 6953 45845 6987
rect 45845 6953 45879 6987
rect 45879 6953 45888 6987
rect 45836 6944 45888 6953
rect 45928 6944 45980 6996
rect 58348 6944 58400 6996
rect 37188 6808 37240 6860
rect 38660 6808 38712 6860
rect 46388 6808 46440 6860
rect 46664 6808 46716 6860
rect 48780 6808 48832 6860
rect 36728 6740 36780 6792
rect 44548 6740 44600 6792
rect 45468 6740 45520 6792
rect 33232 6672 33284 6724
rect 35624 6672 35676 6724
rect 35808 6672 35860 6724
rect 48228 6740 48280 6792
rect 56876 6783 56928 6792
rect 56876 6749 56885 6783
rect 56885 6749 56919 6783
rect 56919 6749 56928 6783
rect 56876 6740 56928 6749
rect 56968 6740 57020 6792
rect 58716 6672 58768 6724
rect 33048 6604 33100 6656
rect 35900 6604 35952 6656
rect 36452 6604 36504 6656
rect 36728 6604 36780 6656
rect 57980 6604 58032 6656
rect 58256 6647 58308 6656
rect 58256 6613 58265 6647
rect 58265 6613 58299 6647
rect 58299 6613 58308 6647
rect 58256 6604 58308 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 9128 6443 9180 6452
rect 9128 6409 9137 6443
rect 9137 6409 9171 6443
rect 9171 6409 9180 6443
rect 9128 6400 9180 6409
rect 10876 6332 10928 6384
rect 11704 6332 11756 6384
rect 17868 6400 17920 6452
rect 24676 6443 24728 6452
rect 15384 6375 15436 6384
rect 15384 6341 15393 6375
rect 15393 6341 15427 6375
rect 15427 6341 15436 6375
rect 15384 6332 15436 6341
rect 15660 6332 15712 6384
rect 9128 6264 9180 6316
rect 9312 6307 9364 6316
rect 9312 6273 9321 6307
rect 9321 6273 9355 6307
rect 9355 6273 9364 6307
rect 9312 6264 9364 6273
rect 1768 6239 1820 6248
rect 1768 6205 1777 6239
rect 1777 6205 1811 6239
rect 1811 6205 1820 6239
rect 1768 6196 1820 6205
rect 8944 6196 8996 6248
rect 9496 6239 9548 6248
rect 9496 6205 9505 6239
rect 9505 6205 9539 6239
rect 9539 6205 9548 6239
rect 9496 6196 9548 6205
rect 9588 6239 9640 6248
rect 9588 6205 9597 6239
rect 9597 6205 9631 6239
rect 9631 6205 9640 6239
rect 9588 6196 9640 6205
rect 12440 6128 12492 6180
rect 13728 6171 13780 6180
rect 13728 6137 13737 6171
rect 13737 6137 13771 6171
rect 13771 6137 13780 6171
rect 13728 6128 13780 6137
rect 15200 6264 15252 6316
rect 15476 6264 15528 6316
rect 15752 6307 15804 6316
rect 15752 6273 15761 6307
rect 15761 6273 15795 6307
rect 15795 6273 15804 6307
rect 15752 6264 15804 6273
rect 16212 6264 16264 6316
rect 17776 6332 17828 6384
rect 18512 6332 18564 6384
rect 19524 6332 19576 6384
rect 19800 6332 19852 6384
rect 17040 6264 17092 6316
rect 17960 6264 18012 6316
rect 19248 6264 19300 6316
rect 19340 6264 19392 6316
rect 22652 6264 22704 6316
rect 16396 6196 16448 6248
rect 18512 6196 18564 6248
rect 18788 6196 18840 6248
rect 19432 6239 19484 6248
rect 19432 6205 19441 6239
rect 19441 6205 19475 6239
rect 19475 6205 19484 6239
rect 19432 6196 19484 6205
rect 18696 6128 18748 6180
rect 21364 6128 21416 6180
rect 9404 6060 9456 6112
rect 20720 6060 20772 6112
rect 21456 6060 21508 6112
rect 24676 6409 24685 6443
rect 24685 6409 24719 6443
rect 24719 6409 24728 6443
rect 24676 6400 24728 6409
rect 25596 6443 25648 6452
rect 25596 6409 25605 6443
rect 25605 6409 25639 6443
rect 25639 6409 25648 6443
rect 25596 6400 25648 6409
rect 25688 6400 25740 6452
rect 28264 6400 28316 6452
rect 30564 6400 30616 6452
rect 33784 6400 33836 6452
rect 46756 6443 46808 6452
rect 46756 6409 46765 6443
rect 46765 6409 46799 6443
rect 46799 6409 46808 6443
rect 46756 6400 46808 6409
rect 28632 6332 28684 6384
rect 25044 6264 25096 6316
rect 26240 6264 26292 6316
rect 26608 6264 26660 6316
rect 27160 6307 27212 6316
rect 27160 6273 27169 6307
rect 27169 6273 27203 6307
rect 27203 6273 27212 6307
rect 27160 6264 27212 6273
rect 33692 6332 33744 6384
rect 26056 6239 26108 6248
rect 26056 6205 26065 6239
rect 26065 6205 26099 6239
rect 26099 6205 26108 6239
rect 26056 6196 26108 6205
rect 26424 6196 26476 6248
rect 26884 6196 26936 6248
rect 27528 6196 27580 6248
rect 30564 6264 30616 6316
rect 32128 6264 32180 6316
rect 33876 6307 33928 6316
rect 33876 6273 33885 6307
rect 33885 6273 33919 6307
rect 33919 6273 33928 6307
rect 33876 6264 33928 6273
rect 34612 6264 34664 6316
rect 35440 6264 35492 6316
rect 35900 6307 35952 6316
rect 35900 6273 35909 6307
rect 35909 6273 35943 6307
rect 35943 6273 35952 6307
rect 35900 6264 35952 6273
rect 32772 6128 32824 6180
rect 33140 6196 33192 6248
rect 35808 6196 35860 6248
rect 37280 6264 37332 6316
rect 51356 6332 51408 6384
rect 57152 6375 57204 6384
rect 57152 6341 57161 6375
rect 57161 6341 57195 6375
rect 57195 6341 57204 6375
rect 57152 6332 57204 6341
rect 46848 6264 46900 6316
rect 33324 6128 33376 6180
rect 36268 6128 36320 6180
rect 27528 6103 27580 6112
rect 27528 6069 27537 6103
rect 27537 6069 27571 6103
rect 27571 6069 27580 6103
rect 27528 6060 27580 6069
rect 29092 6060 29144 6112
rect 35440 6060 35492 6112
rect 35900 6060 35952 6112
rect 36912 6128 36964 6180
rect 39304 6060 39356 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 9128 5899 9180 5908
rect 9128 5865 9137 5899
rect 9137 5865 9171 5899
rect 9171 5865 9180 5899
rect 9128 5856 9180 5865
rect 7932 5788 7984 5840
rect 9404 5763 9456 5772
rect 9404 5729 9413 5763
rect 9413 5729 9447 5763
rect 9447 5729 9456 5763
rect 9404 5720 9456 5729
rect 9680 5720 9732 5772
rect 9312 5695 9364 5704
rect 1860 5627 1912 5636
rect 1860 5593 1869 5627
rect 1869 5593 1903 5627
rect 1903 5593 1912 5627
rect 1860 5584 1912 5593
rect 9312 5661 9321 5695
rect 9321 5661 9355 5695
rect 9355 5661 9364 5695
rect 9312 5652 9364 5661
rect 9588 5695 9640 5704
rect 9588 5661 9597 5695
rect 9597 5661 9631 5695
rect 9631 5661 9640 5695
rect 9588 5652 9640 5661
rect 10140 5584 10192 5636
rect 10416 5627 10468 5636
rect 10416 5593 10425 5627
rect 10425 5593 10459 5627
rect 10459 5593 10468 5627
rect 10416 5584 10468 5593
rect 7748 5516 7800 5568
rect 11060 5856 11112 5908
rect 12624 5856 12676 5908
rect 13820 5856 13872 5908
rect 11888 5788 11940 5840
rect 16212 5788 16264 5840
rect 16856 5788 16908 5840
rect 19616 5788 19668 5840
rect 23112 5856 23164 5908
rect 23388 5856 23440 5908
rect 26240 5856 26292 5908
rect 29644 5856 29696 5908
rect 29736 5856 29788 5908
rect 30012 5899 30064 5908
rect 30012 5865 30021 5899
rect 30021 5865 30055 5899
rect 30055 5865 30064 5899
rect 30012 5856 30064 5865
rect 15660 5763 15712 5772
rect 15660 5729 15669 5763
rect 15669 5729 15703 5763
rect 15703 5729 15712 5763
rect 15660 5720 15712 5729
rect 15844 5720 15896 5772
rect 15476 5652 15528 5704
rect 16396 5652 16448 5704
rect 17040 5695 17092 5704
rect 17040 5661 17049 5695
rect 17049 5661 17083 5695
rect 17083 5661 17092 5695
rect 17040 5652 17092 5661
rect 17408 5720 17460 5772
rect 17776 5652 17828 5704
rect 18144 5720 18196 5772
rect 18972 5652 19024 5704
rect 19432 5652 19484 5704
rect 19616 5695 19668 5704
rect 19616 5661 19625 5695
rect 19625 5661 19659 5695
rect 19659 5661 19668 5695
rect 19616 5652 19668 5661
rect 20260 5652 20312 5704
rect 23112 5720 23164 5772
rect 21456 5695 21508 5704
rect 21456 5661 21465 5695
rect 21465 5661 21499 5695
rect 21499 5661 21508 5695
rect 21456 5652 21508 5661
rect 23204 5652 23256 5704
rect 26608 5788 26660 5840
rect 28908 5788 28960 5840
rect 14280 5627 14332 5636
rect 14280 5593 14289 5627
rect 14289 5593 14323 5627
rect 14323 5593 14332 5627
rect 14280 5584 14332 5593
rect 13912 5516 13964 5568
rect 15568 5584 15620 5636
rect 16856 5584 16908 5636
rect 23296 5584 23348 5636
rect 18512 5516 18564 5568
rect 18604 5516 18656 5568
rect 21088 5516 21140 5568
rect 24860 5652 24912 5704
rect 26608 5652 26660 5704
rect 28540 5695 28592 5704
rect 28540 5661 28549 5695
rect 28549 5661 28583 5695
rect 28583 5661 28592 5695
rect 28540 5652 28592 5661
rect 28816 5652 28868 5704
rect 23664 5584 23716 5636
rect 28724 5584 28776 5636
rect 30104 5763 30156 5772
rect 30104 5729 30113 5763
rect 30113 5729 30147 5763
rect 30147 5729 30156 5763
rect 30104 5720 30156 5729
rect 30196 5720 30248 5772
rect 32956 5652 33008 5704
rect 33784 5652 33836 5704
rect 35808 5788 35860 5840
rect 37648 5788 37700 5840
rect 35348 5720 35400 5772
rect 48320 5856 48372 5908
rect 38384 5831 38436 5840
rect 38384 5797 38393 5831
rect 38393 5797 38427 5831
rect 38427 5797 38436 5831
rect 38384 5788 38436 5797
rect 40500 5788 40552 5840
rect 41420 5788 41472 5840
rect 34796 5652 34848 5704
rect 35440 5652 35492 5704
rect 37372 5652 37424 5704
rect 37740 5652 37792 5704
rect 38568 5720 38620 5772
rect 26516 5516 26568 5568
rect 27620 5516 27672 5568
rect 31944 5584 31996 5636
rect 34060 5584 34112 5636
rect 38016 5584 38068 5636
rect 38844 5584 38896 5636
rect 55864 5652 55916 5704
rect 57980 5720 58032 5772
rect 58164 5763 58216 5772
rect 58164 5729 58173 5763
rect 58173 5729 58207 5763
rect 58207 5729 58216 5763
rect 58164 5720 58216 5729
rect 57796 5652 57848 5704
rect 31576 5516 31628 5568
rect 31852 5516 31904 5568
rect 34244 5559 34296 5568
rect 34244 5525 34253 5559
rect 34253 5525 34287 5559
rect 34287 5525 34296 5559
rect 34244 5516 34296 5525
rect 36360 5559 36412 5568
rect 36360 5525 36369 5559
rect 36369 5525 36403 5559
rect 36403 5525 36412 5559
rect 36360 5516 36412 5525
rect 37556 5516 37608 5568
rect 38936 5516 38988 5568
rect 40040 5584 40092 5636
rect 41420 5627 41472 5636
rect 41420 5593 41429 5627
rect 41429 5593 41463 5627
rect 41463 5593 41472 5627
rect 57244 5627 57296 5636
rect 41420 5584 41472 5593
rect 57244 5593 57253 5627
rect 57253 5593 57287 5627
rect 57287 5593 57296 5627
rect 57244 5584 57296 5593
rect 39948 5516 40000 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 9588 5312 9640 5364
rect 10140 5355 10192 5364
rect 10140 5321 10149 5355
rect 10149 5321 10183 5355
rect 10183 5321 10192 5355
rect 10140 5312 10192 5321
rect 8944 5287 8996 5296
rect 8944 5253 8953 5287
rect 8953 5253 8987 5287
rect 8987 5253 8996 5287
rect 8944 5244 8996 5253
rect 14280 5312 14332 5364
rect 18604 5312 18656 5364
rect 19340 5312 19392 5364
rect 26056 5312 26108 5364
rect 31116 5355 31168 5364
rect 1584 5219 1636 5228
rect 1584 5185 1593 5219
rect 1593 5185 1627 5219
rect 1627 5185 1636 5219
rect 1584 5176 1636 5185
rect 8116 5176 8168 5228
rect 9588 5176 9640 5228
rect 10048 5176 10100 5228
rect 10508 5219 10560 5228
rect 10508 5185 10517 5219
rect 10517 5185 10551 5219
rect 10551 5185 10560 5219
rect 10508 5176 10560 5185
rect 11980 5176 12032 5228
rect 14740 5244 14792 5296
rect 20904 5244 20956 5296
rect 26424 5244 26476 5296
rect 27988 5244 28040 5296
rect 28448 5287 28500 5296
rect 28448 5253 28457 5287
rect 28457 5253 28491 5287
rect 28491 5253 28500 5287
rect 30840 5287 30892 5296
rect 28448 5244 28500 5253
rect 1768 5151 1820 5160
rect 1768 5117 1777 5151
rect 1777 5117 1811 5151
rect 1811 5117 1820 5151
rect 1768 5108 1820 5117
rect 8760 5040 8812 5092
rect 10600 5151 10652 5160
rect 10600 5117 10609 5151
rect 10609 5117 10643 5151
rect 10643 5117 10652 5151
rect 10600 5108 10652 5117
rect 13728 5176 13780 5228
rect 13820 5108 13872 5160
rect 17408 5176 17460 5228
rect 18052 5219 18104 5228
rect 18052 5185 18061 5219
rect 18061 5185 18095 5219
rect 18095 5185 18104 5219
rect 18052 5176 18104 5185
rect 19340 5176 19392 5228
rect 20260 5176 20312 5228
rect 20628 5176 20680 5228
rect 23388 5176 23440 5228
rect 17132 5108 17184 5160
rect 19892 5151 19944 5160
rect 19892 5117 19901 5151
rect 19901 5117 19935 5151
rect 19935 5117 19944 5151
rect 19892 5108 19944 5117
rect 21364 5108 21416 5160
rect 22468 5108 22520 5160
rect 24952 5176 25004 5228
rect 25136 5219 25188 5228
rect 25136 5185 25145 5219
rect 25145 5185 25179 5219
rect 25179 5185 25188 5219
rect 25136 5176 25188 5185
rect 24216 5108 24268 5160
rect 27160 5219 27212 5228
rect 27160 5185 27169 5219
rect 27169 5185 27203 5219
rect 27203 5185 27212 5219
rect 27160 5176 27212 5185
rect 27252 5219 27304 5228
rect 27252 5185 27261 5219
rect 27261 5185 27295 5219
rect 27295 5185 27304 5219
rect 28540 5219 28592 5228
rect 27252 5176 27304 5185
rect 28540 5185 28549 5219
rect 28549 5185 28583 5219
rect 28583 5185 28592 5219
rect 28540 5176 28592 5185
rect 29736 5219 29788 5228
rect 26332 5151 26384 5160
rect 26332 5117 26341 5151
rect 26341 5117 26375 5151
rect 26375 5117 26384 5151
rect 26332 5108 26384 5117
rect 26516 5151 26568 5160
rect 26516 5117 26525 5151
rect 26525 5117 26559 5151
rect 26559 5117 26568 5151
rect 26516 5108 26568 5117
rect 26884 5108 26936 5160
rect 28080 5108 28132 5160
rect 29736 5185 29745 5219
rect 29745 5185 29779 5219
rect 29779 5185 29788 5219
rect 29736 5176 29788 5185
rect 30564 5176 30616 5228
rect 30840 5253 30849 5287
rect 30849 5253 30883 5287
rect 30883 5253 30892 5287
rect 30840 5244 30892 5253
rect 31116 5321 31125 5355
rect 31125 5321 31159 5355
rect 31159 5321 31168 5355
rect 31116 5312 31168 5321
rect 31392 5312 31444 5364
rect 35624 5312 35676 5364
rect 32588 5244 32640 5296
rect 33784 5244 33836 5296
rect 34796 5244 34848 5296
rect 31024 5219 31076 5228
rect 31024 5185 31033 5219
rect 31033 5185 31067 5219
rect 31067 5185 31076 5219
rect 31024 5176 31076 5185
rect 31300 5176 31352 5228
rect 35348 5176 35400 5228
rect 35900 5219 35952 5228
rect 35900 5185 35909 5219
rect 35909 5185 35943 5219
rect 35943 5185 35952 5219
rect 35900 5176 35952 5185
rect 36452 5244 36504 5296
rect 40224 5244 40276 5296
rect 40684 5312 40736 5364
rect 42800 5355 42852 5364
rect 42800 5321 42809 5355
rect 42809 5321 42843 5355
rect 42843 5321 42852 5355
rect 42800 5312 42852 5321
rect 43168 5312 43220 5364
rect 37188 5176 37240 5228
rect 37372 5176 37424 5228
rect 37648 5219 37700 5228
rect 7104 4972 7156 5024
rect 9680 4972 9732 5024
rect 16672 4972 16724 5024
rect 20628 4972 20680 5024
rect 24676 5015 24728 5024
rect 24676 4981 24685 5015
rect 24685 4981 24719 5015
rect 24719 4981 24728 5015
rect 24676 4972 24728 4981
rect 24952 4972 25004 5024
rect 28632 5040 28684 5092
rect 28816 5040 28868 5092
rect 30196 5040 30248 5092
rect 25780 4972 25832 5024
rect 25872 4972 25924 5024
rect 27528 5015 27580 5024
rect 27528 4981 27537 5015
rect 27537 4981 27571 5015
rect 27571 4981 27580 5015
rect 27528 4972 27580 4981
rect 28080 5015 28132 5024
rect 28080 4981 28089 5015
rect 28089 4981 28123 5015
rect 28123 4981 28132 5015
rect 28080 4972 28132 4981
rect 30012 4972 30064 5024
rect 33232 5108 33284 5160
rect 34796 5108 34848 5160
rect 35440 5108 35492 5160
rect 37648 5185 37657 5219
rect 37657 5185 37691 5219
rect 37691 5185 37700 5219
rect 37648 5176 37700 5185
rect 38936 5219 38988 5228
rect 38936 5185 38945 5219
rect 38945 5185 38979 5219
rect 38979 5185 38988 5219
rect 38936 5176 38988 5185
rect 39672 5219 39724 5228
rect 39672 5185 39681 5219
rect 39681 5185 39715 5219
rect 39715 5185 39724 5219
rect 39672 5176 39724 5185
rect 33048 5083 33100 5092
rect 33048 5049 33057 5083
rect 33057 5049 33091 5083
rect 33091 5049 33100 5083
rect 33048 5040 33100 5049
rect 34152 4972 34204 5024
rect 34428 5015 34480 5024
rect 34428 4981 34437 5015
rect 34437 4981 34471 5015
rect 34471 4981 34480 5015
rect 34428 4972 34480 4981
rect 38476 5040 38528 5092
rect 40500 5176 40552 5228
rect 41604 5176 41656 5228
rect 41880 5176 41932 5228
rect 42892 5176 42944 5228
rect 44180 5219 44232 5228
rect 44180 5185 44189 5219
rect 44189 5185 44223 5219
rect 44223 5185 44232 5219
rect 44180 5176 44232 5185
rect 44548 5176 44600 5228
rect 45652 5176 45704 5228
rect 48780 5219 48832 5228
rect 48780 5185 48789 5219
rect 48789 5185 48823 5219
rect 48823 5185 48832 5219
rect 48780 5176 48832 5185
rect 40224 5040 40276 5092
rect 46756 5108 46808 5160
rect 58072 5219 58124 5228
rect 58072 5185 58081 5219
rect 58081 5185 58115 5219
rect 58115 5185 58124 5219
rect 58072 5176 58124 5185
rect 44456 5040 44508 5092
rect 44640 5040 44692 5092
rect 45192 5040 45244 5092
rect 34704 4972 34756 5024
rect 37832 5015 37884 5024
rect 37832 4981 37841 5015
rect 37841 4981 37875 5015
rect 37875 4981 37884 5015
rect 37832 4972 37884 4981
rect 38844 4972 38896 5024
rect 39212 4972 39264 5024
rect 40684 4972 40736 5024
rect 41144 4972 41196 5024
rect 41696 4972 41748 5024
rect 44272 4972 44324 5024
rect 45008 5015 45060 5024
rect 45008 4981 45017 5015
rect 45017 4981 45051 5015
rect 45051 4981 45060 5015
rect 45008 4972 45060 4981
rect 51448 4972 51500 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 1584 4700 1636 4752
rect 9864 4768 9916 4820
rect 11244 4768 11296 4820
rect 13728 4768 13780 4820
rect 17500 4768 17552 4820
rect 24676 4768 24728 4820
rect 25596 4768 25648 4820
rect 10048 4700 10100 4752
rect 12072 4700 12124 4752
rect 9680 4632 9732 4684
rect 9772 4675 9824 4684
rect 9772 4641 9781 4675
rect 9781 4641 9815 4675
rect 9815 4641 9824 4675
rect 9772 4632 9824 4641
rect 9956 4675 10008 4684
rect 9956 4641 9965 4675
rect 9965 4641 9999 4675
rect 9999 4641 10008 4675
rect 9956 4632 10008 4641
rect 10416 4632 10468 4684
rect 14740 4743 14792 4752
rect 14740 4709 14749 4743
rect 14749 4709 14783 4743
rect 14783 4709 14792 4743
rect 14740 4700 14792 4709
rect 15200 4700 15252 4752
rect 15660 4700 15712 4752
rect 17316 4700 17368 4752
rect 19892 4700 19944 4752
rect 23756 4700 23808 4752
rect 18880 4632 18932 4684
rect 18972 4632 19024 4684
rect 21180 4675 21232 4684
rect 4620 4564 4672 4616
rect 9864 4607 9916 4616
rect 9864 4573 9873 4607
rect 9873 4573 9907 4607
rect 9907 4573 9916 4607
rect 9864 4564 9916 4573
rect 6920 4539 6972 4548
rect 6920 4505 6929 4539
rect 6929 4505 6963 4539
rect 6963 4505 6972 4539
rect 6920 4496 6972 4505
rect 8300 4496 8352 4548
rect 7012 4471 7064 4480
rect 7012 4437 7021 4471
rect 7021 4437 7055 4471
rect 7055 4437 7064 4471
rect 7012 4428 7064 4437
rect 7564 4428 7616 4480
rect 8852 4496 8904 4548
rect 9772 4428 9824 4480
rect 12992 4564 13044 4616
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 14740 4564 14792 4616
rect 16396 4564 16448 4616
rect 16580 4607 16632 4616
rect 16580 4573 16589 4607
rect 16589 4573 16623 4607
rect 16623 4573 16632 4607
rect 16580 4564 16632 4573
rect 17868 4564 17920 4616
rect 18328 4564 18380 4616
rect 11796 4496 11848 4548
rect 13084 4496 13136 4548
rect 18052 4496 18104 4548
rect 19432 4564 19484 4616
rect 20076 4564 20128 4616
rect 21180 4641 21189 4675
rect 21189 4641 21223 4675
rect 21223 4641 21232 4675
rect 21180 4632 21232 4641
rect 25228 4700 25280 4752
rect 25872 4700 25924 4752
rect 25964 4700 26016 4752
rect 27712 4811 27764 4820
rect 27712 4777 27721 4811
rect 27721 4777 27755 4811
rect 27755 4777 27764 4811
rect 27712 4768 27764 4777
rect 31760 4768 31812 4820
rect 35348 4768 35400 4820
rect 26332 4700 26384 4752
rect 31852 4700 31904 4752
rect 24952 4632 25004 4684
rect 21364 4564 21416 4616
rect 22008 4564 22060 4616
rect 22376 4607 22428 4616
rect 22376 4573 22385 4607
rect 22385 4573 22419 4607
rect 22419 4573 22428 4607
rect 22376 4564 22428 4573
rect 19892 4539 19944 4548
rect 19892 4505 19901 4539
rect 19901 4505 19935 4539
rect 19935 4505 19944 4539
rect 19892 4496 19944 4505
rect 17224 4428 17276 4480
rect 17316 4428 17368 4480
rect 20536 4471 20588 4480
rect 20536 4437 20545 4471
rect 20545 4437 20579 4471
rect 20579 4437 20588 4471
rect 20536 4428 20588 4437
rect 24492 4564 24544 4616
rect 24676 4607 24728 4616
rect 24676 4573 24685 4607
rect 24685 4573 24719 4607
rect 24719 4573 24728 4607
rect 24676 4564 24728 4573
rect 25412 4564 25464 4616
rect 25964 4564 26016 4616
rect 26424 4607 26476 4616
rect 26424 4573 26433 4607
rect 26433 4573 26467 4607
rect 26467 4573 26476 4607
rect 26424 4564 26476 4573
rect 28356 4632 28408 4684
rect 31944 4632 31996 4684
rect 32036 4632 32088 4684
rect 32864 4632 32916 4684
rect 22744 4496 22796 4548
rect 25504 4496 25556 4548
rect 25596 4496 25648 4548
rect 26240 4496 26292 4548
rect 28724 4564 28776 4616
rect 30564 4564 30616 4616
rect 27068 4496 27120 4548
rect 27620 4496 27672 4548
rect 28632 4496 28684 4548
rect 21456 4428 21508 4480
rect 23572 4428 23624 4480
rect 23756 4471 23808 4480
rect 23756 4437 23765 4471
rect 23765 4437 23799 4471
rect 23799 4437 23808 4471
rect 23756 4428 23808 4437
rect 23940 4428 23992 4480
rect 28816 4428 28868 4480
rect 30012 4428 30064 4480
rect 32220 4564 32272 4616
rect 33140 4564 33192 4616
rect 36544 4700 36596 4752
rect 36820 4700 36872 4752
rect 40776 4768 40828 4820
rect 37372 4632 37424 4684
rect 37924 4632 37976 4684
rect 35624 4564 35676 4616
rect 37832 4564 37884 4616
rect 40316 4700 40368 4752
rect 39028 4632 39080 4684
rect 39488 4632 39540 4684
rect 31116 4496 31168 4548
rect 31576 4428 31628 4480
rect 32220 4428 32272 4480
rect 32496 4539 32548 4548
rect 32496 4505 32505 4539
rect 32505 4505 32539 4539
rect 32539 4505 32548 4539
rect 32496 4496 32548 4505
rect 34520 4496 34572 4548
rect 37188 4496 37240 4548
rect 38200 4496 38252 4548
rect 40960 4564 41012 4616
rect 43352 4700 43404 4752
rect 43628 4768 43680 4820
rect 44272 4768 44324 4820
rect 56508 4768 56560 4820
rect 50712 4700 50764 4752
rect 38752 4496 38804 4548
rect 40132 4539 40184 4548
rect 33416 4428 33468 4480
rect 33508 4428 33560 4480
rect 36360 4428 36412 4480
rect 37464 4428 37516 4480
rect 39212 4428 39264 4480
rect 40132 4505 40141 4539
rect 40141 4505 40175 4539
rect 40175 4505 40184 4539
rect 40132 4496 40184 4505
rect 40776 4496 40828 4548
rect 42524 4496 42576 4548
rect 42984 4632 43036 4684
rect 43628 4607 43680 4616
rect 40316 4428 40368 4480
rect 43628 4573 43637 4607
rect 43637 4573 43671 4607
rect 43671 4573 43680 4607
rect 43628 4564 43680 4573
rect 43904 4632 43956 4684
rect 53104 4632 53156 4684
rect 43996 4607 44048 4616
rect 43996 4573 44010 4607
rect 44010 4573 44044 4607
rect 44044 4573 44048 4607
rect 43996 4564 44048 4573
rect 51264 4607 51316 4616
rect 51264 4573 51273 4607
rect 51273 4573 51307 4607
rect 51307 4573 51316 4607
rect 51264 4564 51316 4573
rect 51448 4607 51500 4616
rect 51448 4573 51457 4607
rect 51457 4573 51491 4607
rect 51491 4573 51500 4607
rect 51448 4564 51500 4573
rect 57796 4564 57848 4616
rect 45100 4496 45152 4548
rect 46020 4539 46072 4548
rect 46020 4505 46029 4539
rect 46029 4505 46063 4539
rect 46063 4505 46072 4539
rect 46020 4496 46072 4505
rect 44364 4428 44416 4480
rect 53564 4428 53616 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 7012 4224 7064 4276
rect 6460 4156 6512 4208
rect 7288 4156 7340 4208
rect 8484 4156 8536 4208
rect 5908 4088 5960 4140
rect 6828 4131 6880 4140
rect 6828 4097 6837 4131
rect 6837 4097 6871 4131
rect 6871 4097 6880 4131
rect 6828 4088 6880 4097
rect 8208 4088 8260 4140
rect 9588 4156 9640 4208
rect 11704 4156 11756 4208
rect 12440 4156 12492 4208
rect 9496 4088 9548 4140
rect 11152 4131 11204 4140
rect 1768 4063 1820 4072
rect 1768 4029 1777 4063
rect 1777 4029 1811 4063
rect 1811 4029 1820 4063
rect 1768 4020 1820 4029
rect 6644 3952 6696 4004
rect 8668 3952 8720 4004
rect 8944 4020 8996 4072
rect 9220 4063 9272 4072
rect 9220 4029 9229 4063
rect 9229 4029 9263 4063
rect 9263 4029 9272 4063
rect 9220 4020 9272 4029
rect 9404 4063 9456 4072
rect 9404 4029 9413 4063
rect 9413 4029 9447 4063
rect 9447 4029 9456 4063
rect 9404 4020 9456 4029
rect 9588 4020 9640 4072
rect 10324 4020 10376 4072
rect 11152 4097 11161 4131
rect 11161 4097 11195 4131
rect 11195 4097 11204 4131
rect 11152 4088 11204 4097
rect 12072 4088 12124 4140
rect 14280 4199 14332 4208
rect 14280 4165 14289 4199
rect 14289 4165 14323 4199
rect 14323 4165 14332 4199
rect 14280 4156 14332 4165
rect 16580 4224 16632 4276
rect 19340 4224 19392 4276
rect 22376 4224 22428 4276
rect 24124 4224 24176 4276
rect 24676 4267 24728 4276
rect 24676 4233 24685 4267
rect 24685 4233 24719 4267
rect 24719 4233 24728 4267
rect 24676 4224 24728 4233
rect 27804 4224 27856 4276
rect 27988 4224 28040 4276
rect 31576 4224 31628 4276
rect 33324 4224 33376 4276
rect 33692 4224 33744 4276
rect 34152 4224 34204 4276
rect 52460 4224 52512 4276
rect 53104 4267 53156 4276
rect 53104 4233 53113 4267
rect 53113 4233 53147 4267
rect 53147 4233 53156 4267
rect 53104 4224 53156 4233
rect 19524 4156 19576 4208
rect 20536 4156 20588 4208
rect 12348 4020 12400 4072
rect 10048 3952 10100 4004
rect 7472 3927 7524 3936
rect 7472 3893 7481 3927
rect 7481 3893 7515 3927
rect 7515 3893 7524 3927
rect 7472 3884 7524 3893
rect 8576 3884 8628 3936
rect 9036 3884 9088 3936
rect 11244 3952 11296 4004
rect 12900 4063 12952 4072
rect 12900 4029 12909 4063
rect 12909 4029 12943 4063
rect 12943 4029 12952 4063
rect 12900 4020 12952 4029
rect 12992 3952 13044 4004
rect 16948 4131 17000 4140
rect 14832 4020 14884 4072
rect 11152 3884 11204 3936
rect 16948 4097 16957 4131
rect 16957 4097 16991 4131
rect 16991 4097 17000 4131
rect 16948 4088 17000 4097
rect 17592 4088 17644 4140
rect 16120 4063 16172 4072
rect 16120 4029 16129 4063
rect 16129 4029 16163 4063
rect 16163 4029 16172 4063
rect 16120 4020 16172 4029
rect 18604 4088 18656 4140
rect 19064 4088 19116 4140
rect 18512 4020 18564 4072
rect 19616 4088 19668 4140
rect 19800 4088 19852 4140
rect 20996 4088 21048 4140
rect 16764 3884 16816 3936
rect 18144 3884 18196 3936
rect 18420 3884 18472 3936
rect 18788 3927 18840 3936
rect 18788 3893 18797 3927
rect 18797 3893 18831 3927
rect 18831 3893 18840 3927
rect 18788 3884 18840 3893
rect 18972 3952 19024 4004
rect 19432 4020 19484 4072
rect 19984 4063 20036 4072
rect 19984 4029 19993 4063
rect 19993 4029 20027 4063
rect 20027 4029 20036 4063
rect 19984 4020 20036 4029
rect 19432 3884 19484 3936
rect 19616 3884 19668 3936
rect 24860 4156 24912 4208
rect 28080 4156 28132 4208
rect 28172 4156 28224 4208
rect 22376 4131 22428 4140
rect 22376 4097 22385 4131
rect 22385 4097 22419 4131
rect 22419 4097 22428 4131
rect 22376 4088 22428 4097
rect 23572 4131 23624 4140
rect 23572 4097 23606 4131
rect 23606 4097 23624 4131
rect 23572 4088 23624 4097
rect 28448 4088 28500 4140
rect 29736 4131 29788 4140
rect 29736 4097 29745 4131
rect 29745 4097 29779 4131
rect 29779 4097 29788 4131
rect 29736 4088 29788 4097
rect 30472 4156 30524 4208
rect 30932 4156 30984 4208
rect 33416 4156 33468 4208
rect 37372 4156 37424 4208
rect 37648 4156 37700 4208
rect 42064 4156 42116 4208
rect 45376 4156 45428 4208
rect 46112 4156 46164 4208
rect 52000 4156 52052 4208
rect 52828 4156 52880 4208
rect 53380 4156 53432 4208
rect 57888 4156 57940 4208
rect 31208 4088 31260 4140
rect 31484 4088 31536 4140
rect 34428 4131 34480 4140
rect 34428 4097 34437 4131
rect 34437 4097 34471 4131
rect 34471 4097 34480 4131
rect 34428 4088 34480 4097
rect 23020 4020 23072 4072
rect 23296 4063 23348 4072
rect 23296 4029 23305 4063
rect 23305 4029 23339 4063
rect 23339 4029 23348 4063
rect 23296 4020 23348 4029
rect 24676 4020 24728 4072
rect 24492 3952 24544 4004
rect 27252 3952 27304 4004
rect 21364 3927 21416 3936
rect 21364 3893 21373 3927
rect 21373 3893 21407 3927
rect 21407 3893 21416 3927
rect 21364 3884 21416 3893
rect 23204 3884 23256 3936
rect 25964 3884 26016 3936
rect 29644 4020 29696 4072
rect 32772 4063 32824 4072
rect 32772 4029 32781 4063
rect 32781 4029 32815 4063
rect 32815 4029 32824 4063
rect 32772 4020 32824 4029
rect 32864 4063 32916 4072
rect 32864 4029 32873 4063
rect 32873 4029 32907 4063
rect 32907 4029 32916 4063
rect 32864 4020 32916 4029
rect 29000 3952 29052 4004
rect 30104 3952 30156 4004
rect 28724 3927 28776 3936
rect 28724 3893 28733 3927
rect 28733 3893 28767 3927
rect 28767 3893 28776 3927
rect 28724 3884 28776 3893
rect 30840 3927 30892 3936
rect 30840 3893 30849 3927
rect 30849 3893 30883 3927
rect 30883 3893 30892 3927
rect 30840 3884 30892 3893
rect 32036 3884 32088 3936
rect 32680 3952 32732 4004
rect 34060 4020 34112 4072
rect 36268 4131 36320 4140
rect 36268 4097 36277 4131
rect 36277 4097 36311 4131
rect 36311 4097 36320 4131
rect 36268 4088 36320 4097
rect 37188 4088 37240 4140
rect 38844 4131 38896 4140
rect 38844 4097 38878 4131
rect 38878 4097 38896 4131
rect 38844 4088 38896 4097
rect 33416 3884 33468 3936
rect 33600 3884 33652 3936
rect 35440 3884 35492 3936
rect 35716 4020 35768 4072
rect 36728 4020 36780 4072
rect 35624 3952 35676 4004
rect 37832 3884 37884 3936
rect 40132 4088 40184 4140
rect 40592 4131 40644 4140
rect 40592 4097 40601 4131
rect 40601 4097 40635 4131
rect 40635 4097 40644 4131
rect 40592 4088 40644 4097
rect 41512 4131 41564 4140
rect 41512 4097 41521 4131
rect 41521 4097 41555 4131
rect 41555 4097 41564 4131
rect 41512 4088 41564 4097
rect 43352 4131 43404 4140
rect 43352 4097 43361 4131
rect 43361 4097 43395 4131
rect 43395 4097 43404 4131
rect 43352 4088 43404 4097
rect 39856 4020 39908 4072
rect 43444 4063 43496 4072
rect 43444 4029 43453 4063
rect 43453 4029 43487 4063
rect 43487 4029 43496 4063
rect 43444 4020 43496 4029
rect 39948 3995 40000 4004
rect 39948 3961 39957 3995
rect 39957 3961 39991 3995
rect 39991 3961 40000 3995
rect 39948 3952 40000 3961
rect 43536 3952 43588 4004
rect 44364 4088 44416 4140
rect 45928 4131 45980 4140
rect 45928 4097 45937 4131
rect 45937 4097 45971 4131
rect 45971 4097 45980 4131
rect 45928 4088 45980 4097
rect 44732 4020 44784 4072
rect 45468 4020 45520 4072
rect 44364 3952 44416 4004
rect 44824 3952 44876 4004
rect 48136 4088 48188 4140
rect 51724 4088 51776 4140
rect 54484 4088 54536 4140
rect 58348 4131 58400 4140
rect 58348 4097 58357 4131
rect 58357 4097 58391 4131
rect 58391 4097 58400 4131
rect 58348 4088 58400 4097
rect 46848 4020 46900 4072
rect 53472 4020 53524 4072
rect 48412 3995 48464 4004
rect 48412 3961 48421 3995
rect 48421 3961 48455 3995
rect 48455 3961 48464 3995
rect 48412 3952 48464 3961
rect 53656 3952 53708 4004
rect 42524 3884 42576 3936
rect 43628 3884 43680 3936
rect 43996 3884 44048 3936
rect 45928 3884 45980 3936
rect 47032 3884 47084 3936
rect 47308 3884 47360 3936
rect 47492 3884 47544 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 7012 3680 7064 3732
rect 7472 3680 7524 3732
rect 6000 3655 6052 3664
rect 6000 3621 6009 3655
rect 6009 3621 6043 3655
rect 6043 3621 6052 3655
rect 6000 3612 6052 3621
rect 7564 3655 7616 3664
rect 7564 3621 7573 3655
rect 7573 3621 7607 3655
rect 7607 3621 7616 3655
rect 7564 3612 7616 3621
rect 7656 3655 7708 3664
rect 7656 3621 7665 3655
rect 7665 3621 7699 3655
rect 7699 3621 7708 3655
rect 7656 3612 7708 3621
rect 6184 3476 6236 3528
rect 8852 3612 8904 3664
rect 10600 3680 10652 3732
rect 11888 3655 11940 3664
rect 11888 3621 11897 3655
rect 11897 3621 11931 3655
rect 11931 3621 11940 3655
rect 11888 3612 11940 3621
rect 12624 3655 12676 3664
rect 12624 3621 12633 3655
rect 12633 3621 12667 3655
rect 12667 3621 12676 3655
rect 12624 3612 12676 3621
rect 12900 3680 12952 3732
rect 14648 3680 14700 3732
rect 17960 3680 18012 3732
rect 18512 3680 18564 3732
rect 19248 3680 19300 3732
rect 13544 3612 13596 3664
rect 13820 3612 13872 3664
rect 15936 3655 15988 3664
rect 15936 3621 15945 3655
rect 15945 3621 15979 3655
rect 15979 3621 15988 3655
rect 15936 3612 15988 3621
rect 20352 3680 20404 3732
rect 20720 3680 20772 3732
rect 20996 3655 21048 3664
rect 12532 3544 12584 3596
rect 20996 3621 21005 3655
rect 21005 3621 21039 3655
rect 21039 3621 21048 3655
rect 20996 3612 21048 3621
rect 9588 3519 9640 3528
rect 9588 3485 9597 3519
rect 9597 3485 9631 3519
rect 9631 3485 9640 3519
rect 9588 3476 9640 3485
rect 1860 3451 1912 3460
rect 1860 3417 1869 3451
rect 1869 3417 1903 3451
rect 1903 3417 1912 3451
rect 1860 3408 1912 3417
rect 7012 3340 7064 3392
rect 8208 3408 8260 3460
rect 8392 3408 8444 3460
rect 8484 3408 8536 3460
rect 8852 3408 8904 3460
rect 9864 3519 9916 3528
rect 9864 3485 9873 3519
rect 9873 3485 9907 3519
rect 9907 3485 9916 3519
rect 9864 3476 9916 3485
rect 10324 3476 10376 3528
rect 13360 3476 13412 3528
rect 15108 3476 15160 3528
rect 15660 3519 15712 3528
rect 15660 3485 15669 3519
rect 15669 3485 15703 3519
rect 15703 3485 15712 3519
rect 15660 3476 15712 3485
rect 17224 3476 17276 3528
rect 17500 3519 17552 3528
rect 17500 3485 17509 3519
rect 17509 3485 17543 3519
rect 17543 3485 17552 3519
rect 17500 3476 17552 3485
rect 18972 3544 19024 3596
rect 18420 3519 18472 3528
rect 18420 3485 18429 3519
rect 18429 3485 18463 3519
rect 18463 3485 18472 3519
rect 19524 3544 19576 3596
rect 21180 3544 21232 3596
rect 22376 3544 22428 3596
rect 18420 3476 18472 3485
rect 9956 3408 10008 3460
rect 12348 3451 12400 3460
rect 12348 3417 12357 3451
rect 12357 3417 12391 3451
rect 12391 3417 12400 3451
rect 12348 3408 12400 3417
rect 8576 3340 8628 3392
rect 9220 3340 9272 3392
rect 12532 3340 12584 3392
rect 12808 3340 12860 3392
rect 14188 3408 14240 3460
rect 15568 3408 15620 3460
rect 16580 3408 16632 3460
rect 17776 3408 17828 3460
rect 13544 3340 13596 3392
rect 23296 3476 23348 3528
rect 23756 3680 23808 3732
rect 27712 3723 27764 3732
rect 27712 3689 27721 3723
rect 27721 3689 27755 3723
rect 27755 3689 27764 3723
rect 27712 3680 27764 3689
rect 33692 3723 33744 3732
rect 28264 3612 28316 3664
rect 29736 3612 29788 3664
rect 33692 3689 33701 3723
rect 33701 3689 33735 3723
rect 33735 3689 33744 3723
rect 33692 3680 33744 3689
rect 37188 3680 37240 3732
rect 39672 3680 39724 3732
rect 42432 3680 42484 3732
rect 43720 3680 43772 3732
rect 44180 3680 44232 3732
rect 44364 3680 44416 3732
rect 47032 3723 47084 3732
rect 47032 3689 47041 3723
rect 47041 3689 47075 3723
rect 47075 3689 47084 3723
rect 47032 3680 47084 3689
rect 47860 3680 47912 3732
rect 48596 3680 48648 3732
rect 49424 3723 49476 3732
rect 49424 3689 49433 3723
rect 49433 3689 49467 3723
rect 49467 3689 49476 3723
rect 49424 3680 49476 3689
rect 52460 3680 52512 3732
rect 54208 3723 54260 3732
rect 54208 3689 54217 3723
rect 54217 3689 54251 3723
rect 54251 3689 54260 3723
rect 54208 3680 54260 3689
rect 55036 3680 55088 3732
rect 26516 3476 26568 3528
rect 18788 3408 18840 3460
rect 19524 3340 19576 3392
rect 19984 3408 20036 3460
rect 20076 3408 20128 3460
rect 20904 3408 20956 3460
rect 21824 3451 21876 3460
rect 21088 3340 21140 3392
rect 21456 3383 21508 3392
rect 21456 3349 21465 3383
rect 21465 3349 21499 3383
rect 21499 3349 21508 3383
rect 21456 3340 21508 3349
rect 21824 3417 21833 3451
rect 21833 3417 21867 3451
rect 21867 3417 21876 3451
rect 21824 3408 21876 3417
rect 23204 3408 23256 3460
rect 24124 3408 24176 3460
rect 26700 3451 26752 3460
rect 26700 3417 26709 3451
rect 26709 3417 26743 3451
rect 26743 3417 26752 3451
rect 26700 3408 26752 3417
rect 27436 3544 27488 3596
rect 29368 3544 29420 3596
rect 30104 3544 30156 3596
rect 32220 3544 32272 3596
rect 28724 3476 28776 3528
rect 27252 3451 27304 3460
rect 27252 3417 27261 3451
rect 27261 3417 27295 3451
rect 27295 3417 27304 3451
rect 27252 3408 27304 3417
rect 27344 3408 27396 3460
rect 29092 3476 29144 3528
rect 31576 3519 31628 3528
rect 31576 3485 31585 3519
rect 31585 3485 31619 3519
rect 31619 3485 31628 3519
rect 31576 3476 31628 3485
rect 32036 3476 32088 3528
rect 29276 3408 29328 3460
rect 30196 3408 30248 3460
rect 33232 3544 33284 3596
rect 36084 3544 36136 3596
rect 36820 3544 36872 3596
rect 32864 3476 32916 3528
rect 33324 3476 33376 3528
rect 33416 3476 33468 3528
rect 33968 3476 34020 3528
rect 34704 3476 34756 3528
rect 36176 3519 36228 3528
rect 36176 3485 36185 3519
rect 36185 3485 36219 3519
rect 36219 3485 36228 3519
rect 36176 3476 36228 3485
rect 38292 3612 38344 3664
rect 40776 3612 40828 3664
rect 41972 3655 42024 3664
rect 39120 3544 39172 3596
rect 40132 3587 40184 3596
rect 40132 3553 40141 3587
rect 40141 3553 40175 3587
rect 40175 3553 40184 3587
rect 40132 3544 40184 3553
rect 40868 3587 40920 3596
rect 40868 3553 40877 3587
rect 40877 3553 40911 3587
rect 40911 3553 40920 3587
rect 40868 3544 40920 3553
rect 41972 3621 41981 3655
rect 41981 3621 42015 3655
rect 42015 3621 42024 3655
rect 41972 3612 42024 3621
rect 42708 3612 42760 3664
rect 43352 3544 43404 3596
rect 43812 3544 43864 3596
rect 37372 3476 37424 3528
rect 37556 3519 37608 3528
rect 37556 3485 37565 3519
rect 37565 3485 37599 3519
rect 37599 3485 37608 3519
rect 37556 3476 37608 3485
rect 23664 3340 23716 3392
rect 26884 3340 26936 3392
rect 28080 3383 28132 3392
rect 28080 3349 28089 3383
rect 28089 3349 28123 3383
rect 28123 3349 28132 3383
rect 28080 3340 28132 3349
rect 28448 3340 28500 3392
rect 32864 3340 32916 3392
rect 32956 3340 33008 3392
rect 34336 3408 34388 3460
rect 34612 3408 34664 3460
rect 35716 3408 35768 3460
rect 33324 3340 33376 3392
rect 33876 3340 33928 3392
rect 34060 3340 34112 3392
rect 35440 3340 35492 3392
rect 36544 3340 36596 3392
rect 40960 3476 41012 3528
rect 41144 3519 41196 3528
rect 41144 3485 41153 3519
rect 41153 3485 41187 3519
rect 41187 3485 41196 3519
rect 41144 3476 41196 3485
rect 38292 3408 38344 3460
rect 42524 3476 42576 3528
rect 44088 3544 44140 3596
rect 45100 3612 45152 3664
rect 46020 3612 46072 3664
rect 47400 3612 47452 3664
rect 44180 3519 44232 3528
rect 44180 3485 44189 3519
rect 44189 3485 44223 3519
rect 44223 3485 44232 3519
rect 44180 3476 44232 3485
rect 46848 3544 46900 3596
rect 47584 3476 47636 3528
rect 48780 3476 48832 3528
rect 49332 3476 49384 3528
rect 56876 3587 56928 3596
rect 56876 3553 56885 3587
rect 56885 3553 56919 3587
rect 56919 3553 56928 3587
rect 56876 3544 56928 3553
rect 51724 3476 51776 3528
rect 53196 3476 53248 3528
rect 54760 3476 54812 3528
rect 38568 3340 38620 3392
rect 40592 3340 40644 3392
rect 43260 3340 43312 3392
rect 46756 3408 46808 3460
rect 43628 3340 43680 3392
rect 45468 3340 45520 3392
rect 49884 3408 49936 3460
rect 50620 3408 50672 3460
rect 51264 3408 51316 3460
rect 52276 3408 52328 3460
rect 53564 3408 53616 3460
rect 50804 3340 50856 3392
rect 57244 3340 57296 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 8024 3136 8076 3188
rect 9864 3136 9916 3188
rect 12900 3136 12952 3188
rect 15936 3136 15988 3188
rect 23204 3179 23256 3188
rect 5908 3068 5960 3120
rect 4620 3000 4672 3052
rect 9128 3068 9180 3120
rect 1768 2975 1820 2984
rect 1768 2941 1777 2975
rect 1777 2941 1811 2975
rect 1811 2941 1820 2975
rect 1768 2932 1820 2941
rect 7564 2932 7616 2984
rect 9220 3000 9272 3052
rect 9588 3043 9640 3052
rect 9588 3009 9597 3043
rect 9597 3009 9631 3043
rect 9631 3009 9640 3043
rect 9588 3000 9640 3009
rect 10048 3000 10100 3052
rect 10324 3068 10376 3120
rect 12808 3000 12860 3052
rect 8208 2932 8260 2984
rect 8392 2932 8444 2984
rect 8760 2907 8812 2916
rect 8760 2873 8769 2907
rect 8769 2873 8803 2907
rect 8803 2873 8812 2907
rect 8760 2864 8812 2873
rect 7104 2796 7156 2848
rect 7380 2796 7432 2848
rect 7932 2839 7984 2848
rect 7932 2805 7941 2839
rect 7941 2805 7975 2839
rect 7975 2805 7984 2839
rect 7932 2796 7984 2805
rect 8024 2796 8076 2848
rect 9956 2932 10008 2984
rect 11796 2932 11848 2984
rect 12256 2932 12308 2984
rect 13636 3000 13688 3052
rect 14372 3000 14424 3052
rect 14464 3043 14516 3052
rect 14464 3009 14473 3043
rect 14473 3009 14507 3043
rect 14507 3009 14516 3043
rect 14464 3000 14516 3009
rect 15292 3000 15344 3052
rect 15660 3000 15712 3052
rect 18144 3068 18196 3120
rect 18236 3068 18288 3120
rect 17776 3043 17828 3052
rect 17776 3009 17785 3043
rect 17785 3009 17819 3043
rect 17819 3009 17828 3043
rect 17776 3000 17828 3009
rect 9588 2864 9640 2916
rect 10600 2864 10652 2916
rect 11796 2796 11848 2848
rect 13912 2796 13964 2848
rect 14004 2796 14056 2848
rect 16948 2864 17000 2916
rect 19708 3000 19760 3052
rect 21456 3068 21508 3120
rect 23204 3145 23213 3179
rect 23213 3145 23247 3179
rect 23247 3145 23256 3179
rect 23204 3136 23256 3145
rect 27436 3136 27488 3188
rect 23664 3111 23716 3120
rect 23664 3077 23673 3111
rect 23673 3077 23707 3111
rect 23707 3077 23716 3111
rect 23664 3068 23716 3077
rect 26516 3068 26568 3120
rect 29552 3136 29604 3188
rect 33048 3136 33100 3188
rect 30748 3068 30800 3120
rect 21916 3000 21968 3052
rect 22284 3043 22336 3052
rect 22284 3009 22293 3043
rect 22293 3009 22327 3043
rect 22327 3009 22336 3043
rect 22284 3000 22336 3009
rect 22376 3000 22428 3052
rect 23572 3043 23624 3052
rect 17960 2864 18012 2916
rect 19524 2864 19576 2916
rect 16580 2796 16632 2848
rect 16856 2796 16908 2848
rect 19156 2796 19208 2848
rect 23572 3009 23581 3043
rect 23581 3009 23615 3043
rect 23615 3009 23624 3043
rect 23572 3000 23624 3009
rect 20628 2864 20680 2916
rect 22192 2864 22244 2916
rect 23940 2932 23992 2984
rect 23848 2864 23900 2916
rect 25228 2864 25280 2916
rect 27344 3000 27396 3052
rect 27528 3043 27580 3052
rect 27528 3009 27537 3043
rect 27537 3009 27571 3043
rect 27571 3009 27580 3043
rect 27528 3000 27580 3009
rect 29000 3000 29052 3052
rect 30840 3043 30892 3052
rect 30840 3009 30849 3043
rect 30849 3009 30883 3043
rect 30883 3009 30892 3043
rect 30840 3000 30892 3009
rect 32220 3068 32272 3120
rect 35624 3068 35676 3120
rect 34520 3000 34572 3052
rect 37096 3136 37148 3188
rect 37740 3136 37792 3188
rect 38384 3136 38436 3188
rect 38844 3136 38896 3188
rect 36544 3111 36596 3120
rect 36544 3077 36553 3111
rect 36553 3077 36587 3111
rect 36587 3077 36596 3111
rect 36544 3068 36596 3077
rect 40224 3068 40276 3120
rect 40408 3111 40460 3120
rect 40408 3077 40417 3111
rect 40417 3077 40451 3111
rect 40451 3077 40460 3111
rect 40408 3068 40460 3077
rect 40684 3136 40736 3188
rect 44916 3136 44968 3188
rect 45192 3179 45244 3188
rect 45192 3145 45201 3179
rect 45201 3145 45235 3179
rect 45235 3145 45244 3179
rect 45192 3136 45244 3145
rect 46480 3179 46532 3188
rect 46480 3145 46489 3179
rect 46489 3145 46523 3179
rect 46523 3145 46532 3179
rect 46480 3136 46532 3145
rect 47952 3179 48004 3188
rect 47952 3145 47961 3179
rect 47961 3145 47995 3179
rect 47995 3145 48004 3179
rect 47952 3136 48004 3145
rect 48872 3179 48924 3188
rect 48872 3145 48881 3179
rect 48881 3145 48915 3179
rect 48915 3145 48924 3179
rect 48872 3136 48924 3145
rect 49792 3179 49844 3188
rect 49792 3145 49801 3179
rect 49801 3145 49835 3179
rect 49835 3145 49844 3179
rect 49792 3136 49844 3145
rect 50712 3179 50764 3188
rect 50712 3145 50721 3179
rect 50721 3145 50755 3179
rect 50755 3145 50764 3179
rect 50712 3136 50764 3145
rect 52184 3179 52236 3188
rect 52184 3145 52193 3179
rect 52193 3145 52227 3179
rect 52227 3145 52236 3179
rect 52184 3136 52236 3145
rect 55220 3136 55272 3188
rect 36268 3043 36320 3052
rect 36268 3009 36277 3043
rect 36277 3009 36311 3043
rect 36311 3009 36320 3043
rect 36268 3000 36320 3009
rect 36452 3043 36504 3052
rect 36452 3009 36459 3043
rect 36459 3009 36504 3043
rect 36452 3000 36504 3009
rect 26424 2975 26476 2984
rect 26424 2941 26433 2975
rect 26433 2941 26467 2975
rect 26467 2941 26476 2975
rect 26424 2932 26476 2941
rect 28172 2864 28224 2916
rect 20260 2796 20312 2848
rect 20904 2796 20956 2848
rect 22008 2796 22060 2848
rect 23296 2796 23348 2848
rect 23388 2796 23440 2848
rect 27160 2796 27212 2848
rect 28356 2932 28408 2984
rect 29092 2932 29144 2984
rect 30748 2932 30800 2984
rect 31576 2932 31628 2984
rect 33508 2975 33560 2984
rect 33508 2941 33517 2975
rect 33517 2941 33551 2975
rect 33551 2941 33560 2975
rect 33508 2932 33560 2941
rect 33876 2932 33928 2984
rect 34336 2932 34388 2984
rect 36084 2932 36136 2984
rect 38108 2932 38160 2984
rect 38936 3000 38988 3052
rect 39304 3000 39356 3052
rect 39580 3000 39632 3052
rect 41144 3043 41196 3052
rect 38568 2932 38620 2984
rect 41144 3009 41153 3043
rect 41153 3009 41187 3043
rect 41187 3009 41196 3043
rect 41144 3000 41196 3009
rect 41512 3000 41564 3052
rect 42156 3000 42208 3052
rect 42616 3043 42668 3052
rect 42616 3009 42625 3043
rect 42625 3009 42659 3043
rect 42659 3009 42668 3043
rect 42616 3000 42668 3009
rect 42984 3000 43036 3052
rect 43168 3000 43220 3052
rect 43628 3043 43680 3052
rect 43628 3009 43637 3043
rect 43637 3009 43671 3043
rect 43671 3009 43680 3043
rect 43628 3000 43680 3009
rect 45560 3068 45612 3120
rect 49332 3068 49384 3120
rect 49516 3068 49568 3120
rect 50896 3068 50948 3120
rect 54944 3068 54996 3120
rect 58164 3111 58216 3120
rect 58164 3077 58173 3111
rect 58173 3077 58207 3111
rect 58207 3077 58216 3111
rect 58164 3068 58216 3077
rect 44364 3000 44416 3052
rect 45008 3000 45060 3052
rect 46204 3000 46256 3052
rect 47032 3000 47084 3052
rect 48412 3000 48464 3052
rect 48964 3000 49016 3052
rect 50160 3000 50212 3052
rect 51448 3000 51500 3052
rect 53932 3000 53984 3052
rect 54208 3000 54260 3052
rect 55312 3000 55364 3052
rect 58256 3000 58308 3052
rect 43352 2975 43404 2984
rect 36820 2864 36872 2916
rect 37464 2864 37516 2916
rect 43352 2941 43361 2975
rect 43361 2941 43395 2975
rect 43395 2941 43404 2975
rect 43352 2932 43404 2941
rect 43536 2975 43588 2984
rect 43536 2941 43545 2975
rect 43545 2941 43579 2975
rect 43579 2941 43588 2975
rect 43536 2932 43588 2941
rect 45284 2932 45336 2984
rect 29092 2796 29144 2848
rect 32496 2796 32548 2848
rect 34520 2796 34572 2848
rect 40960 2864 41012 2916
rect 43444 2864 43496 2916
rect 45376 2864 45428 2916
rect 47676 2932 47728 2984
rect 53288 2932 53340 2984
rect 49608 2864 49660 2916
rect 49700 2864 49752 2916
rect 50804 2864 50856 2916
rect 41604 2796 41656 2848
rect 42340 2796 42392 2848
rect 44180 2796 44232 2848
rect 47860 2796 47912 2848
rect 50436 2796 50488 2848
rect 50528 2796 50580 2848
rect 53472 2864 53524 2916
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 7196 2592 7248 2644
rect 7380 2592 7432 2644
rect 9036 2592 9088 2644
rect 7656 2524 7708 2576
rect 11244 2592 11296 2644
rect 14004 2592 14056 2644
rect 17408 2592 17460 2644
rect 11060 2524 11112 2576
rect 12624 2524 12676 2576
rect 19432 2592 19484 2644
rect 19524 2592 19576 2644
rect 21364 2592 21416 2644
rect 26792 2592 26844 2644
rect 1584 2431 1636 2440
rect 1584 2397 1593 2431
rect 1593 2397 1627 2431
rect 1627 2397 1636 2431
rect 1584 2388 1636 2397
rect 4528 2388 4580 2440
rect 1860 2363 1912 2372
rect 1860 2329 1869 2363
rect 1869 2329 1903 2363
rect 1903 2329 1912 2363
rect 1860 2320 1912 2329
rect 7840 2456 7892 2508
rect 5724 2320 5776 2372
rect 9312 2456 9364 2508
rect 13636 2456 13688 2508
rect 4436 2295 4488 2304
rect 4436 2261 4445 2295
rect 4445 2261 4479 2295
rect 4479 2261 4488 2295
rect 4436 2252 4488 2261
rect 7380 2320 7432 2372
rect 7656 2363 7708 2372
rect 7656 2329 7665 2363
rect 7665 2329 7699 2363
rect 7699 2329 7708 2363
rect 7656 2320 7708 2329
rect 9496 2363 9548 2372
rect 9496 2329 9505 2363
rect 9505 2329 9539 2363
rect 9539 2329 9548 2363
rect 9496 2320 9548 2329
rect 11796 2388 11848 2440
rect 12348 2431 12400 2440
rect 12348 2397 12357 2431
rect 12357 2397 12391 2431
rect 12391 2397 12400 2431
rect 12348 2388 12400 2397
rect 12992 2388 13044 2440
rect 16856 2456 16908 2508
rect 17776 2456 17828 2508
rect 20628 2524 20680 2576
rect 17316 2388 17368 2440
rect 17500 2431 17552 2440
rect 17500 2397 17509 2431
rect 17509 2397 17543 2431
rect 17543 2397 17552 2431
rect 17500 2388 17552 2397
rect 18420 2431 18472 2440
rect 18420 2397 18429 2431
rect 18429 2397 18463 2431
rect 18463 2397 18472 2431
rect 18420 2388 18472 2397
rect 11428 2320 11480 2372
rect 6920 2252 6972 2304
rect 7472 2252 7524 2304
rect 7748 2295 7800 2304
rect 7748 2261 7757 2295
rect 7757 2261 7791 2295
rect 7791 2261 7800 2295
rect 7748 2252 7800 2261
rect 8484 2295 8536 2304
rect 8484 2261 8493 2295
rect 8493 2261 8527 2295
rect 8527 2261 8536 2295
rect 8484 2252 8536 2261
rect 9220 2252 9272 2304
rect 10876 2252 10928 2304
rect 15752 2320 15804 2372
rect 15016 2252 15068 2304
rect 19892 2431 19944 2440
rect 19892 2397 19901 2431
rect 19901 2397 19935 2431
rect 19935 2397 19944 2431
rect 19892 2388 19944 2397
rect 22008 2456 22060 2508
rect 24400 2456 24452 2508
rect 20076 2320 20128 2372
rect 19432 2295 19484 2304
rect 19432 2261 19441 2295
rect 19441 2261 19475 2295
rect 19475 2261 19484 2295
rect 19432 2252 19484 2261
rect 19524 2252 19576 2304
rect 20444 2252 20496 2304
rect 20996 2431 21048 2440
rect 20996 2397 21005 2431
rect 21005 2397 21039 2431
rect 21039 2397 21048 2431
rect 20996 2388 21048 2397
rect 22652 2431 22704 2440
rect 22652 2397 22661 2431
rect 22661 2397 22695 2431
rect 22695 2397 22704 2431
rect 22652 2388 22704 2397
rect 23480 2320 23532 2372
rect 23664 2388 23716 2440
rect 28816 2524 28868 2576
rect 29368 2456 29420 2508
rect 27896 2388 27948 2440
rect 28908 2388 28960 2440
rect 29184 2388 29236 2440
rect 30932 2388 30984 2440
rect 34336 2592 34388 2644
rect 34244 2524 34296 2576
rect 31300 2456 31352 2508
rect 34520 2456 34572 2508
rect 32404 2388 32456 2440
rect 34888 2431 34940 2440
rect 34888 2397 34897 2431
rect 34897 2397 34931 2431
rect 34931 2397 34940 2431
rect 34888 2388 34940 2397
rect 23756 2320 23808 2372
rect 24952 2320 25004 2372
rect 25504 2363 25556 2372
rect 25504 2329 25513 2363
rect 25513 2329 25547 2363
rect 25547 2329 25556 2363
rect 25504 2320 25556 2329
rect 28816 2320 28868 2372
rect 29920 2320 29972 2372
rect 30472 2363 30524 2372
rect 30472 2329 30481 2363
rect 30481 2329 30515 2363
rect 30515 2329 30524 2363
rect 30472 2320 30524 2329
rect 31024 2320 31076 2372
rect 31852 2320 31904 2372
rect 33876 2320 33928 2372
rect 36912 2456 36964 2508
rect 40868 2592 40920 2644
rect 42800 2592 42852 2644
rect 45008 2592 45060 2644
rect 45376 2635 45428 2644
rect 45376 2601 45385 2635
rect 45385 2601 45419 2635
rect 45419 2601 45428 2635
rect 45376 2592 45428 2601
rect 46112 2592 46164 2644
rect 47124 2635 47176 2644
rect 47124 2601 47133 2635
rect 47133 2601 47167 2635
rect 47167 2601 47176 2635
rect 47124 2592 47176 2601
rect 47768 2592 47820 2644
rect 48688 2592 48740 2644
rect 49056 2592 49108 2644
rect 58256 2635 58308 2644
rect 50712 2524 50764 2576
rect 37924 2388 37976 2440
rect 21640 2252 21692 2304
rect 23388 2252 23440 2304
rect 26148 2252 26200 2304
rect 26884 2252 26936 2304
rect 32128 2252 32180 2304
rect 36636 2320 36688 2372
rect 42984 2456 43036 2508
rect 45008 2456 45060 2508
rect 40224 2388 40276 2440
rect 42616 2431 42668 2440
rect 42616 2397 42625 2431
rect 42625 2397 42659 2431
rect 42659 2397 42668 2431
rect 42616 2388 42668 2397
rect 42800 2431 42852 2440
rect 42800 2397 42807 2431
rect 42807 2397 42852 2431
rect 42800 2388 42852 2397
rect 43536 2388 43588 2440
rect 39304 2320 39356 2372
rect 44456 2388 44508 2440
rect 45192 2431 45244 2440
rect 45192 2397 45201 2431
rect 45201 2397 45235 2431
rect 45235 2397 45244 2431
rect 45192 2388 45244 2397
rect 46480 2388 46532 2440
rect 49240 2456 49292 2508
rect 49700 2388 49752 2440
rect 50436 2431 50488 2440
rect 50436 2397 50445 2431
rect 50445 2397 50479 2431
rect 50479 2397 50488 2431
rect 50436 2388 50488 2397
rect 50988 2456 51040 2508
rect 58256 2601 58265 2635
rect 58265 2601 58299 2635
rect 58299 2601 58308 2635
rect 58256 2592 58308 2601
rect 53656 2388 53708 2440
rect 55036 2388 55088 2440
rect 57244 2388 57296 2440
rect 58164 2431 58216 2440
rect 58164 2397 58173 2431
rect 58173 2397 58207 2431
rect 58207 2397 58216 2431
rect 58164 2388 58216 2397
rect 43904 2363 43956 2372
rect 43904 2329 43913 2363
rect 43913 2329 43947 2363
rect 43947 2329 43956 2363
rect 43904 2320 43956 2329
rect 45928 2320 45980 2372
rect 35532 2252 35584 2304
rect 42248 2252 42300 2304
rect 43352 2252 43404 2304
rect 44180 2252 44232 2304
rect 47308 2320 47360 2372
rect 50068 2252 50120 2304
rect 52552 2320 52604 2372
rect 57336 2363 57388 2372
rect 57336 2329 57345 2363
rect 57345 2329 57379 2363
rect 57379 2329 57388 2363
rect 57336 2320 57388 2329
rect 51264 2295 51316 2304
rect 51264 2261 51273 2295
rect 51273 2261 51307 2295
rect 51307 2261 51316 2295
rect 51264 2252 51316 2261
rect 53104 2295 53156 2304
rect 53104 2261 53113 2295
rect 53113 2261 53147 2295
rect 53147 2261 53156 2295
rect 53104 2252 53156 2261
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 1584 2048 1636 2100
rect 4436 1980 4488 2032
rect 8668 1980 8720 2032
rect 9496 1980 9548 2032
rect 12808 1980 12860 2032
rect 8484 1912 8536 1964
rect 11336 1912 11388 1964
rect 19432 2048 19484 2100
rect 27988 2048 28040 2100
rect 41052 2048 41104 2100
rect 43352 2048 43404 2100
rect 43628 2048 43680 2100
rect 50712 2048 50764 2100
rect 18420 1980 18472 2032
rect 22836 1980 22888 2032
rect 23756 1980 23808 2032
rect 26700 1912 26752 1964
rect 26976 1912 27028 1964
rect 34888 1912 34940 1964
rect 7656 1844 7708 1896
rect 11152 1844 11204 1896
rect 7748 1776 7800 1828
rect 12716 1776 12768 1828
rect 13176 1776 13228 1828
rect 23664 1776 23716 1828
rect 37004 1980 37056 2032
rect 42248 1980 42300 2032
rect 39764 1912 39816 1964
rect 51264 1912 51316 1964
rect 36912 1844 36964 1896
rect 53104 1844 53156 1896
rect 7472 1708 7524 1760
rect 13268 1708 13320 1760
rect 17316 1708 17368 1760
rect 20168 1708 20220 1760
rect 26056 1708 26108 1760
rect 43076 1708 43128 1760
rect 36912 1640 36964 1692
rect 37924 1640 37976 1692
rect 43904 1640 43956 1692
rect 26424 1504 26476 1556
rect 28540 1504 28592 1556
rect 35716 1504 35768 1556
rect 36728 1504 36780 1556
rect 6920 1436 6972 1488
rect 10048 1436 10100 1488
rect 5724 1368 5776 1420
rect 9496 1368 9548 1420
rect 26148 1368 26200 1420
rect 28264 1368 28316 1420
rect 35992 1368 36044 1420
rect 37464 1368 37516 1420
rect 36820 1300 36872 1352
rect 37832 1300 37884 1352
rect 46940 1300 46992 1352
rect 55956 1300 56008 1352
rect 35440 1164 35492 1216
rect 38568 1164 38620 1216
rect 39028 1028 39080 1080
rect 45192 1028 45244 1080
<< metal2 >>
rect 846 63200 902 64000
rect 1582 63200 1638 64000
rect 2318 63322 2374 64000
rect 3054 63322 3110 64000
rect 3790 63322 3846 64000
rect 4526 63322 4582 64000
rect 5262 63322 5318 64000
rect 5998 63322 6054 64000
rect 6734 63322 6790 64000
rect 2318 63294 2636 63322
rect 2318 63200 2374 63294
rect 860 59022 888 63200
rect 1596 61962 1624 63200
rect 1596 61934 1808 61962
rect 1674 61840 1730 61849
rect 1674 61775 1730 61784
rect 1688 61198 1716 61775
rect 1676 61192 1728 61198
rect 1676 61134 1728 61140
rect 1584 60716 1636 60722
rect 1584 60658 1636 60664
rect 1596 60489 1624 60658
rect 1582 60480 1638 60489
rect 1582 60415 1638 60424
rect 1676 60036 1728 60042
rect 1676 59978 1728 59984
rect 1688 59809 1716 59978
rect 1674 59800 1730 59809
rect 1674 59735 1730 59744
rect 1780 59702 1808 61934
rect 2608 60110 2636 63294
rect 3054 63294 3280 63322
rect 3054 63200 3110 63294
rect 2780 61192 2832 61198
rect 2778 61160 2780 61169
rect 2832 61160 2834 61169
rect 2778 61095 2834 61104
rect 3252 60790 3280 63294
rect 3790 63294 4016 63322
rect 3790 63200 3846 63294
rect 3988 60790 4016 63294
rect 4526 63294 4660 63322
rect 4526 63200 4582 63294
rect 4214 61500 4522 61509
rect 4214 61498 4220 61500
rect 4276 61498 4300 61500
rect 4356 61498 4380 61500
rect 4436 61498 4460 61500
rect 4516 61498 4522 61500
rect 4276 61446 4278 61498
rect 4458 61446 4460 61498
rect 4214 61444 4220 61446
rect 4276 61444 4300 61446
rect 4356 61444 4380 61446
rect 4436 61444 4460 61446
rect 4516 61444 4522 61446
rect 4214 61435 4522 61444
rect 4632 61198 4660 63294
rect 5092 63294 5318 63322
rect 5092 61198 5120 63294
rect 5262 63200 5318 63294
rect 5736 63294 6054 63322
rect 5736 61198 5764 63294
rect 5998 63200 6054 63294
rect 6656 63294 6790 63322
rect 6656 61198 6684 63294
rect 6734 63200 6790 63294
rect 7470 63322 7526 64000
rect 7470 63294 7604 63322
rect 7470 63200 7526 63294
rect 7576 61198 7604 63294
rect 8206 63200 8262 64000
rect 8942 63322 8998 64000
rect 8942 63294 9076 63322
rect 8942 63200 8998 63294
rect 7656 61396 7708 61402
rect 7656 61338 7708 61344
rect 4620 61192 4672 61198
rect 4620 61134 4672 61140
rect 5080 61192 5132 61198
rect 5080 61134 5132 61140
rect 5724 61192 5776 61198
rect 5724 61134 5776 61140
rect 6644 61192 6696 61198
rect 6644 61134 6696 61140
rect 7564 61192 7616 61198
rect 7564 61134 7616 61140
rect 5632 61124 5684 61130
rect 5632 61066 5684 61072
rect 6920 61124 6972 61130
rect 6920 61066 6972 61072
rect 4712 61056 4764 61062
rect 4712 60998 4764 61004
rect 5172 61056 5224 61062
rect 5172 60998 5224 61004
rect 3240 60784 3292 60790
rect 3240 60726 3292 60732
rect 3976 60784 4028 60790
rect 3976 60726 4028 60732
rect 4620 60580 4672 60586
rect 4620 60522 4672 60528
rect 3332 60512 3384 60518
rect 3332 60454 3384 60460
rect 3344 60314 3372 60454
rect 4214 60412 4522 60421
rect 4214 60410 4220 60412
rect 4276 60410 4300 60412
rect 4356 60410 4380 60412
rect 4436 60410 4460 60412
rect 4516 60410 4522 60412
rect 4276 60358 4278 60410
rect 4458 60358 4460 60410
rect 4214 60356 4220 60358
rect 4276 60356 4300 60358
rect 4356 60356 4380 60358
rect 4436 60356 4460 60358
rect 4516 60356 4522 60358
rect 4214 60347 4522 60356
rect 3332 60308 3384 60314
rect 3332 60250 3384 60256
rect 2596 60104 2648 60110
rect 2596 60046 2648 60052
rect 2044 60036 2096 60042
rect 2044 59978 2096 59984
rect 1768 59696 1820 59702
rect 1768 59638 1820 59644
rect 1676 59628 1728 59634
rect 1676 59570 1728 59576
rect 1688 59129 1716 59570
rect 1952 59424 2004 59430
rect 1952 59366 2004 59372
rect 1674 59120 1730 59129
rect 1964 59090 1992 59366
rect 1674 59055 1730 59064
rect 1952 59084 2004 59090
rect 1952 59026 2004 59032
rect 848 59016 900 59022
rect 848 58958 900 58964
rect 2056 58682 2084 59978
rect 2504 59968 2556 59974
rect 2504 59910 2556 59916
rect 2320 59424 2372 59430
rect 2320 59366 2372 59372
rect 2044 58676 2096 58682
rect 2044 58618 2096 58624
rect 1584 58540 1636 58546
rect 1584 58482 1636 58488
rect 1596 58449 1624 58482
rect 1582 58440 1638 58449
rect 1582 58375 1638 58384
rect 1584 57928 1636 57934
rect 1584 57870 1636 57876
rect 1596 57769 1624 57870
rect 1582 57760 1638 57769
rect 1582 57695 1638 57704
rect 1584 57452 1636 57458
rect 1584 57394 1636 57400
rect 1596 57089 1624 57394
rect 1768 57248 1820 57254
rect 1768 57190 1820 57196
rect 1582 57080 1638 57089
rect 1582 57015 1638 57024
rect 1676 56772 1728 56778
rect 1676 56714 1728 56720
rect 1688 56409 1716 56714
rect 1780 56506 1808 57190
rect 2044 56772 2096 56778
rect 2044 56714 2096 56720
rect 1768 56500 1820 56506
rect 1768 56442 1820 56448
rect 2056 56438 2084 56714
rect 2044 56432 2096 56438
rect 1674 56400 1730 56409
rect 2044 56374 2096 56380
rect 1674 56335 1730 56344
rect 1768 55888 1820 55894
rect 1768 55830 1820 55836
rect 1674 55720 1730 55729
rect 1674 55655 1676 55664
rect 1728 55655 1730 55664
rect 1676 55626 1728 55632
rect 1780 55418 1808 55830
rect 1768 55412 1820 55418
rect 1768 55354 1820 55360
rect 1584 55276 1636 55282
rect 1584 55218 1636 55224
rect 1596 55049 1624 55218
rect 1582 55040 1638 55049
rect 1582 54975 1638 54984
rect 1676 54596 1728 54602
rect 1676 54538 1728 54544
rect 1688 54369 1716 54538
rect 1674 54360 1730 54369
rect 1674 54295 1730 54304
rect 1584 54188 1636 54194
rect 1584 54130 1636 54136
rect 1596 53689 1624 54130
rect 1768 53984 1820 53990
rect 1768 53926 1820 53932
rect 1582 53680 1638 53689
rect 1582 53615 1638 53624
rect 1780 53582 1808 53926
rect 1768 53576 1820 53582
rect 1768 53518 1820 53524
rect 1676 53100 1728 53106
rect 1676 53042 1728 53048
rect 1688 53009 1716 53042
rect 1674 53000 1730 53009
rect 1674 52935 1730 52944
rect 1584 52488 1636 52494
rect 1584 52430 1636 52436
rect 1596 52329 1624 52430
rect 1582 52320 1638 52329
rect 1582 52255 1638 52264
rect 1676 52012 1728 52018
rect 1676 51954 1728 51960
rect 1688 51649 1716 51954
rect 1674 51640 1730 51649
rect 1674 51575 1730 51584
rect 1676 51332 1728 51338
rect 1676 51274 1728 51280
rect 1688 50969 1716 51274
rect 1674 50960 1730 50969
rect 1674 50895 1730 50904
rect 1674 50280 1730 50289
rect 1674 50215 1676 50224
rect 1728 50215 1730 50224
rect 2044 50244 2096 50250
rect 1676 50186 1728 50192
rect 2044 50186 2096 50192
rect 1584 49836 1636 49842
rect 1584 49778 1636 49784
rect 1596 49609 1624 49778
rect 1582 49600 1638 49609
rect 1582 49535 1638 49544
rect 1584 49224 1636 49230
rect 1584 49166 1636 49172
rect 1596 48929 1624 49166
rect 1582 48920 1638 48929
rect 1582 48855 1638 48864
rect 1676 48748 1728 48754
rect 1676 48690 1728 48696
rect 1688 48249 1716 48690
rect 1952 48612 2004 48618
rect 1952 48554 2004 48560
rect 1674 48240 1730 48249
rect 1674 48175 1730 48184
rect 1860 48000 1912 48006
rect 1860 47942 1912 47948
rect 1676 47660 1728 47666
rect 1676 47602 1728 47608
rect 1688 47569 1716 47602
rect 1674 47560 1730 47569
rect 1674 47495 1730 47504
rect 1584 47048 1636 47054
rect 1584 46990 1636 46996
rect 1596 46889 1624 46990
rect 1582 46880 1638 46889
rect 1582 46815 1638 46824
rect 1584 46572 1636 46578
rect 1584 46514 1636 46520
rect 1596 46209 1624 46514
rect 1582 46200 1638 46209
rect 1582 46135 1638 46144
rect 1676 45892 1728 45898
rect 1676 45834 1728 45840
rect 1688 45529 1716 45834
rect 1674 45520 1730 45529
rect 1674 45455 1730 45464
rect 1584 44872 1636 44878
rect 1582 44840 1584 44849
rect 1636 44840 1638 44849
rect 1582 44775 1638 44784
rect 1676 44396 1728 44402
rect 1676 44338 1728 44344
rect 1688 44169 1716 44338
rect 1674 44160 1730 44169
rect 1674 44095 1730 44104
rect 1676 43716 1728 43722
rect 1676 43658 1728 43664
rect 1688 43489 1716 43658
rect 1674 43480 1730 43489
rect 1674 43415 1730 43424
rect 1584 43308 1636 43314
rect 1584 43250 1636 43256
rect 1596 42809 1624 43250
rect 1768 43104 1820 43110
rect 1768 43046 1820 43052
rect 1582 42800 1638 42809
rect 1582 42735 1638 42744
rect 1780 42362 1808 43046
rect 1768 42356 1820 42362
rect 1768 42298 1820 42304
rect 1584 42220 1636 42226
rect 1584 42162 1636 42168
rect 1596 42129 1624 42162
rect 1582 42120 1638 42129
rect 1582 42055 1638 42064
rect 1676 41540 1728 41546
rect 1676 41482 1728 41488
rect 1688 41449 1716 41482
rect 1674 41440 1730 41449
rect 1674 41375 1730 41384
rect 1676 41132 1728 41138
rect 1676 41074 1728 41080
rect 1688 40769 1716 41074
rect 1674 40760 1730 40769
rect 1872 40746 1900 47942
rect 1674 40695 1730 40704
rect 1780 40718 1900 40746
rect 1676 40452 1728 40458
rect 1676 40394 1728 40400
rect 1688 40089 1716 40394
rect 1674 40080 1730 40089
rect 1674 40015 1730 40024
rect 1674 39400 1730 39409
rect 1674 39335 1676 39344
rect 1728 39335 1730 39344
rect 1676 39306 1728 39312
rect 1676 38956 1728 38962
rect 1676 38898 1728 38904
rect 1688 38729 1716 38898
rect 1674 38720 1730 38729
rect 1674 38655 1730 38664
rect 1676 38276 1728 38282
rect 1676 38218 1728 38224
rect 1688 38049 1716 38218
rect 1674 38040 1730 38049
rect 1674 37975 1730 37984
rect 1674 37360 1730 37369
rect 1674 37295 1730 37304
rect 1688 37262 1716 37295
rect 1676 37256 1728 37262
rect 1676 37198 1728 37204
rect 1584 36780 1636 36786
rect 1584 36722 1636 36728
rect 1596 36689 1624 36722
rect 1582 36680 1638 36689
rect 1582 36615 1638 36624
rect 1676 36100 1728 36106
rect 1676 36042 1728 36048
rect 1688 36009 1716 36042
rect 1674 36000 1730 36009
rect 1674 35935 1730 35944
rect 1780 35834 1808 40718
rect 1860 38820 1912 38826
rect 1860 38762 1912 38768
rect 1872 38418 1900 38762
rect 1860 38412 1912 38418
rect 1860 38354 1912 38360
rect 1964 37874 1992 48554
rect 2056 48142 2084 50186
rect 2044 48136 2096 48142
rect 2044 48078 2096 48084
rect 2136 42016 2188 42022
rect 2136 41958 2188 41964
rect 1952 37868 2004 37874
rect 1952 37810 2004 37816
rect 1768 35828 1820 35834
rect 1768 35770 1820 35776
rect 1676 35692 1728 35698
rect 1676 35634 1728 35640
rect 1688 35329 1716 35634
rect 1674 35320 1730 35329
rect 1674 35255 1730 35264
rect 1676 35012 1728 35018
rect 1676 34954 1728 34960
rect 1688 34649 1716 34954
rect 1674 34640 1730 34649
rect 1674 34575 1730 34584
rect 1674 33960 1730 33969
rect 1674 33895 1676 33904
rect 1728 33895 1730 33904
rect 1676 33866 1728 33872
rect 1768 33856 1820 33862
rect 1768 33798 1820 33804
rect 1780 33658 1808 33798
rect 1768 33652 1820 33658
rect 1768 33594 1820 33600
rect 1676 33516 1728 33522
rect 1676 33458 1728 33464
rect 1688 33289 1716 33458
rect 1674 33280 1730 33289
rect 1674 33215 1730 33224
rect 1676 32836 1728 32842
rect 1676 32778 1728 32784
rect 1688 32609 1716 32778
rect 1674 32600 1730 32609
rect 1674 32535 1730 32544
rect 1676 32428 1728 32434
rect 1676 32370 1728 32376
rect 1688 31929 1716 32370
rect 1674 31920 1730 31929
rect 1674 31855 1730 31864
rect 1676 31340 1728 31346
rect 1676 31282 1728 31288
rect 1688 31249 1716 31282
rect 1674 31240 1730 31249
rect 1674 31175 1730 31184
rect 1676 30660 1728 30666
rect 1676 30602 1728 30608
rect 1688 30569 1716 30602
rect 1674 30560 1730 30569
rect 1674 30495 1730 30504
rect 1584 30252 1636 30258
rect 1584 30194 1636 30200
rect 1596 29306 1624 30194
rect 1768 30184 1820 30190
rect 1768 30126 1820 30132
rect 1780 29889 1808 30126
rect 1766 29880 1822 29889
rect 1766 29815 1822 29824
rect 1952 29640 2004 29646
rect 1952 29582 2004 29588
rect 1860 29572 1912 29578
rect 1860 29514 1912 29520
rect 1584 29300 1636 29306
rect 1584 29242 1636 29248
rect 1872 29209 1900 29514
rect 1858 29200 1914 29209
rect 1858 29135 1914 29144
rect 1858 28520 1914 28529
rect 1858 28455 1860 28464
rect 1912 28455 1914 28464
rect 1860 28426 1912 28432
rect 1768 28008 1820 28014
rect 1768 27950 1820 27956
rect 1780 27849 1808 27950
rect 1766 27840 1822 27849
rect 1766 27775 1822 27784
rect 1584 27464 1636 27470
rect 1584 27406 1636 27412
rect 1596 27130 1624 27406
rect 1860 27396 1912 27402
rect 1860 27338 1912 27344
rect 1872 27169 1900 27338
rect 1858 27160 1914 27169
rect 1584 27124 1636 27130
rect 1858 27095 1914 27104
rect 1584 27066 1636 27072
rect 1584 26988 1636 26994
rect 1584 26930 1636 26936
rect 1596 21434 1624 26930
rect 1768 26920 1820 26926
rect 1768 26862 1820 26868
rect 1780 26489 1808 26862
rect 1766 26480 1822 26489
rect 1766 26415 1822 26424
rect 1768 25832 1820 25838
rect 1766 25800 1768 25809
rect 1820 25800 1822 25809
rect 1766 25735 1822 25744
rect 1860 25220 1912 25226
rect 1860 25162 1912 25168
rect 1872 25129 1900 25162
rect 1858 25120 1914 25129
rect 1858 25055 1914 25064
rect 1768 24744 1820 24750
rect 1768 24686 1820 24692
rect 1780 24449 1808 24686
rect 1766 24440 1822 24449
rect 1766 24375 1822 24384
rect 1860 24132 1912 24138
rect 1860 24074 1912 24080
rect 1872 23769 1900 24074
rect 1858 23760 1914 23769
rect 1858 23695 1914 23704
rect 1858 23080 1914 23089
rect 1858 23015 1860 23024
rect 1912 23015 1914 23024
rect 1860 22986 1912 22992
rect 1768 22568 1820 22574
rect 1768 22510 1820 22516
rect 1780 22409 1808 22510
rect 1766 22400 1822 22409
rect 1766 22335 1822 22344
rect 1860 21956 1912 21962
rect 1860 21898 1912 21904
rect 1872 21729 1900 21898
rect 1858 21720 1914 21729
rect 1858 21655 1914 21664
rect 1596 21406 1716 21434
rect 1584 17672 1636 17678
rect 1584 17614 1636 17620
rect 1596 16726 1624 17614
rect 1584 16720 1636 16726
rect 1584 16662 1636 16668
rect 1584 14884 1636 14890
rect 1584 14826 1636 14832
rect 1596 13938 1624 14826
rect 1584 13932 1636 13938
rect 1584 13874 1636 13880
rect 1584 13728 1636 13734
rect 1584 13670 1636 13676
rect 1596 13326 1624 13670
rect 1584 13320 1636 13326
rect 1584 13262 1636 13268
rect 1584 11008 1636 11014
rect 1584 10950 1636 10956
rect 1596 10674 1624 10950
rect 1688 10810 1716 21406
rect 1768 21344 1820 21350
rect 1768 21286 1820 21292
rect 1780 21049 1808 21286
rect 1766 21040 1822 21049
rect 1766 20975 1822 20984
rect 1768 20392 1820 20398
rect 1766 20360 1768 20369
rect 1820 20360 1822 20369
rect 1766 20295 1822 20304
rect 1860 19780 1912 19786
rect 1860 19722 1912 19728
rect 1872 19689 1900 19722
rect 1858 19680 1914 19689
rect 1858 19615 1914 19624
rect 1860 19372 1912 19378
rect 1860 19314 1912 19320
rect 1872 19009 1900 19314
rect 1858 19000 1914 19009
rect 1858 18935 1914 18944
rect 1860 18692 1912 18698
rect 1860 18634 1912 18640
rect 1872 18329 1900 18634
rect 1858 18320 1914 18329
rect 1858 18255 1914 18264
rect 1858 17640 1914 17649
rect 1858 17575 1860 17584
rect 1912 17575 1914 17584
rect 1860 17546 1912 17552
rect 1768 17128 1820 17134
rect 1768 17070 1820 17076
rect 1780 16969 1808 17070
rect 1766 16960 1822 16969
rect 1766 16895 1822 16904
rect 1860 16516 1912 16522
rect 1860 16458 1912 16464
rect 1872 16289 1900 16458
rect 1858 16280 1914 16289
rect 1858 16215 1914 16224
rect 1768 16040 1820 16046
rect 1768 15982 1820 15988
rect 1780 15609 1808 15982
rect 1766 15600 1822 15609
rect 1766 15535 1822 15544
rect 1768 14952 1820 14958
rect 1766 14920 1768 14929
rect 1820 14920 1822 14929
rect 1766 14855 1822 14864
rect 1860 14340 1912 14346
rect 1860 14282 1912 14288
rect 1872 14249 1900 14282
rect 1858 14240 1914 14249
rect 1858 14175 1914 14184
rect 1768 13864 1820 13870
rect 1768 13806 1820 13812
rect 1780 13569 1808 13806
rect 1766 13560 1822 13569
rect 1766 13495 1822 13504
rect 1860 13252 1912 13258
rect 1860 13194 1912 13200
rect 1872 12889 1900 13194
rect 1858 12880 1914 12889
rect 1858 12815 1914 12824
rect 1858 12200 1914 12209
rect 1858 12135 1914 12144
rect 1872 11830 1900 12135
rect 1860 11824 1912 11830
rect 1860 11766 1912 11772
rect 1766 11520 1822 11529
rect 1766 11455 1822 11464
rect 1780 11218 1808 11455
rect 1768 11212 1820 11218
rect 1768 11154 1820 11160
rect 1858 10840 1914 10849
rect 1676 10804 1728 10810
rect 1858 10775 1914 10784
rect 1676 10746 1728 10752
rect 1872 10742 1900 10775
rect 1860 10736 1912 10742
rect 1860 10678 1912 10684
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 1766 10160 1822 10169
rect 1766 10095 1768 10104
rect 1820 10095 1822 10104
rect 1768 10066 1820 10072
rect 1582 10024 1638 10033
rect 1582 9959 1638 9968
rect 1596 9586 1624 9959
rect 1964 9926 1992 29582
rect 2148 27538 2176 41958
rect 2228 39568 2280 39574
rect 2228 39510 2280 39516
rect 2240 37806 2268 39510
rect 2332 39438 2360 59366
rect 2412 48136 2464 48142
rect 2412 48078 2464 48084
rect 2424 39574 2452 48078
rect 2412 39568 2464 39574
rect 2412 39510 2464 39516
rect 2320 39432 2372 39438
rect 2320 39374 2372 39380
rect 2412 39296 2464 39302
rect 2412 39238 2464 39244
rect 2228 37800 2280 37806
rect 2228 37742 2280 37748
rect 2320 37732 2372 37738
rect 2320 37674 2372 37680
rect 2332 33590 2360 37674
rect 2424 36106 2452 39238
rect 2516 36174 2544 59910
rect 4214 59324 4522 59333
rect 4214 59322 4220 59324
rect 4276 59322 4300 59324
rect 4356 59322 4380 59324
rect 4436 59322 4460 59324
rect 4516 59322 4522 59324
rect 4276 59270 4278 59322
rect 4458 59270 4460 59322
rect 4214 59268 4220 59270
rect 4276 59268 4300 59270
rect 4356 59268 4380 59270
rect 4436 59268 4460 59270
rect 4516 59268 4522 59270
rect 4214 59259 4522 59268
rect 4214 58236 4522 58245
rect 4214 58234 4220 58236
rect 4276 58234 4300 58236
rect 4356 58234 4380 58236
rect 4436 58234 4460 58236
rect 4516 58234 4522 58236
rect 4276 58182 4278 58234
rect 4458 58182 4460 58234
rect 4214 58180 4220 58182
rect 4276 58180 4300 58182
rect 4356 58180 4380 58182
rect 4436 58180 4460 58182
rect 4516 58180 4522 58182
rect 4214 58171 4522 58180
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 4068 51944 4120 51950
rect 4068 51886 4120 51892
rect 3976 51332 4028 51338
rect 3976 51274 4028 51280
rect 3988 50998 4016 51274
rect 3976 50992 4028 50998
rect 3976 50934 4028 50940
rect 4080 50930 4108 51886
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 4632 51066 4660 60522
rect 4724 57322 4752 60998
rect 5184 60858 5212 60998
rect 5172 60852 5224 60858
rect 5172 60794 5224 60800
rect 5540 60648 5592 60654
rect 5540 60590 5592 60596
rect 4804 58472 4856 58478
rect 4804 58414 4856 58420
rect 4712 57316 4764 57322
rect 4712 57258 4764 57264
rect 4620 51060 4672 51066
rect 4620 51002 4672 51008
rect 4068 50924 4120 50930
rect 4068 50866 4120 50872
rect 2596 50856 2648 50862
rect 2596 50798 2648 50804
rect 2608 39302 2636 50798
rect 4080 48210 4108 50866
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 2872 48204 2924 48210
rect 2872 48146 2924 48152
rect 4068 48204 4120 48210
rect 4068 48146 4120 48152
rect 2780 39976 2832 39982
rect 2780 39918 2832 39924
rect 2792 39438 2820 39918
rect 2780 39432 2832 39438
rect 2780 39374 2832 39380
rect 2596 39296 2648 39302
rect 2596 39238 2648 39244
rect 2792 38350 2820 39374
rect 2780 38344 2832 38350
rect 2780 38286 2832 38292
rect 2596 37664 2648 37670
rect 2596 37606 2648 37612
rect 2608 37466 2636 37606
rect 2596 37460 2648 37466
rect 2596 37402 2648 37408
rect 2792 37346 2820 38286
rect 2884 37942 2912 48146
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 2872 37936 2924 37942
rect 2872 37878 2924 37884
rect 3056 37868 3108 37874
rect 3056 37810 3108 37816
rect 2688 37324 2740 37330
rect 2792 37318 3004 37346
rect 3068 37330 3096 37810
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 2688 37266 2740 37272
rect 2596 36576 2648 36582
rect 2596 36518 2648 36524
rect 2504 36168 2556 36174
rect 2504 36110 2556 36116
rect 2412 36100 2464 36106
rect 2412 36042 2464 36048
rect 2320 33584 2372 33590
rect 2320 33526 2372 33532
rect 2608 29646 2636 36518
rect 2700 35290 2728 37266
rect 2872 36168 2924 36174
rect 2872 36110 2924 36116
rect 2780 36100 2832 36106
rect 2780 36042 2832 36048
rect 2688 35284 2740 35290
rect 2688 35226 2740 35232
rect 2792 35222 2820 36042
rect 2780 35216 2832 35222
rect 2780 35158 2832 35164
rect 2596 29640 2648 29646
rect 2596 29582 2648 29588
rect 2884 28994 2912 36110
rect 2516 28966 2912 28994
rect 2228 28076 2280 28082
rect 2228 28018 2280 28024
rect 2136 27532 2188 27538
rect 2136 27474 2188 27480
rect 2240 12442 2268 28018
rect 2516 27282 2544 28966
rect 2976 28558 3004 37318
rect 3056 37324 3108 37330
rect 3056 37266 3108 37272
rect 3068 36174 3096 37266
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 3056 36168 3108 36174
rect 3056 36110 3108 36116
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 2964 28552 3016 28558
rect 2964 28494 3016 28500
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 2516 27254 2636 27282
rect 2608 26994 2636 27254
rect 2504 26988 2556 26994
rect 2504 26930 2556 26936
rect 2596 26988 2648 26994
rect 2596 26930 2648 26936
rect 2516 25294 2544 26930
rect 2608 26234 2636 26930
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 2608 26206 2728 26234
rect 2504 25288 2556 25294
rect 2504 25230 2556 25236
rect 2596 25288 2648 25294
rect 2596 25230 2648 25236
rect 2412 19168 2464 19174
rect 2412 19110 2464 19116
rect 2424 18873 2452 19110
rect 2410 18864 2466 18873
rect 2410 18799 2466 18808
rect 2410 18728 2466 18737
rect 2410 18663 2412 18672
rect 2464 18663 2466 18672
rect 2412 18634 2464 18640
rect 2410 17232 2466 17241
rect 2410 17167 2412 17176
rect 2464 17167 2466 17176
rect 2412 17138 2464 17144
rect 2412 16040 2464 16046
rect 2410 16008 2412 16017
rect 2464 16008 2466 16017
rect 2410 15943 2466 15952
rect 2410 14512 2466 14521
rect 2410 14447 2412 14456
rect 2464 14447 2466 14456
rect 2412 14418 2464 14424
rect 2228 12436 2280 12442
rect 2228 12378 2280 12384
rect 2608 10130 2636 25230
rect 2596 10124 2648 10130
rect 2596 10066 2648 10072
rect 1952 9920 2004 9926
rect 1952 9862 2004 9868
rect 1584 9580 1636 9586
rect 1584 9522 1636 9528
rect 1768 9512 1820 9518
rect 1766 9480 1768 9489
rect 1820 9480 1822 9489
rect 1766 9415 1822 9424
rect 1860 8900 1912 8906
rect 1860 8842 1912 8848
rect 1872 8809 1900 8842
rect 1858 8800 1914 8809
rect 1858 8735 1914 8744
rect 1768 8424 1820 8430
rect 1768 8366 1820 8372
rect 1780 8129 1808 8366
rect 1766 8120 1822 8129
rect 2700 8090 2728 26206
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 2872 25220 2924 25226
rect 2872 25162 2924 25168
rect 2884 24206 2912 25162
rect 3056 24812 3108 24818
rect 3056 24754 3108 24760
rect 3068 24410 3096 24754
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 3056 24404 3108 24410
rect 3056 24346 3108 24352
rect 4816 24274 4844 58414
rect 5552 57254 5580 60590
rect 5644 60110 5672 61066
rect 5908 61056 5960 61062
rect 5908 60998 5960 61004
rect 5632 60104 5684 60110
rect 5632 60046 5684 60052
rect 5540 57248 5592 57254
rect 5540 57190 5592 57196
rect 5920 38010 5948 60998
rect 6276 50720 6328 50726
rect 6276 50662 6328 50668
rect 6184 47524 6236 47530
rect 6184 47466 6236 47472
rect 5908 38004 5960 38010
rect 5908 37946 5960 37952
rect 6196 37942 6224 47466
rect 6184 37936 6236 37942
rect 6184 37878 6236 37884
rect 6288 37262 6316 50662
rect 6000 37256 6052 37262
rect 6000 37198 6052 37204
rect 6276 37256 6328 37262
rect 6276 37198 6328 37204
rect 6736 37256 6788 37262
rect 6736 37198 6788 37204
rect 5540 37120 5592 37126
rect 5540 37062 5592 37068
rect 5552 28626 5580 37062
rect 6012 36922 6040 37198
rect 6000 36916 6052 36922
rect 6000 36858 6052 36864
rect 6748 36310 6776 37198
rect 6736 36304 6788 36310
rect 6736 36246 6788 36252
rect 5540 28620 5592 28626
rect 5540 28562 5592 28568
rect 4804 24268 4856 24274
rect 4804 24210 4856 24216
rect 2872 24200 2924 24206
rect 2872 24142 2924 24148
rect 2884 11082 2912 24142
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 6828 21548 6880 21554
rect 6828 21490 6880 21496
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 6840 19378 6868 21490
rect 6828 19372 6880 19378
rect 6828 19314 6880 19320
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 6840 18766 6868 19314
rect 6828 18760 6880 18766
rect 6828 18702 6880 18708
rect 6840 18426 6868 18702
rect 6828 18420 6880 18426
rect 6828 18362 6880 18368
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 6932 13297 6960 61066
rect 7668 60110 7696 61338
rect 8220 60874 8248 63200
rect 8944 61124 8996 61130
rect 8944 61066 8996 61072
rect 8220 60846 8340 60874
rect 8312 60790 8340 60846
rect 8300 60784 8352 60790
rect 8300 60726 8352 60732
rect 7656 60104 7708 60110
rect 7656 60046 7708 60052
rect 8024 59968 8076 59974
rect 8024 59910 8076 59916
rect 8036 52018 8064 59910
rect 8024 52012 8076 52018
rect 8024 51954 8076 51960
rect 7840 51808 7892 51814
rect 7840 51750 7892 51756
rect 7852 26994 7880 51750
rect 8956 28558 8984 61066
rect 9048 60722 9076 63294
rect 9678 63200 9734 64000
rect 10414 63322 10470 64000
rect 10244 63294 10470 63322
rect 9692 61198 9720 63200
rect 10244 61198 10272 63294
rect 10414 63200 10470 63294
rect 11150 63200 11206 64000
rect 11886 63322 11942 64000
rect 12622 63322 12678 64000
rect 13358 63322 13414 64000
rect 14094 63322 14150 64000
rect 14830 63322 14886 64000
rect 15566 63322 15622 64000
rect 16302 63322 16358 64000
rect 11886 63294 12020 63322
rect 11886 63200 11942 63294
rect 11060 61668 11112 61674
rect 11060 61610 11112 61616
rect 9680 61192 9732 61198
rect 9680 61134 9732 61140
rect 10232 61192 10284 61198
rect 10232 61134 10284 61140
rect 11072 61062 11100 61610
rect 11164 61198 11192 63200
rect 11992 61198 12020 63294
rect 12622 63294 12756 63322
rect 12622 63200 12678 63294
rect 12728 61198 12756 63294
rect 13358 63294 13584 63322
rect 13358 63200 13414 63294
rect 11152 61192 11204 61198
rect 11152 61134 11204 61140
rect 11980 61192 12032 61198
rect 11980 61134 12032 61140
rect 12716 61192 12768 61198
rect 12992 61192 13044 61198
rect 12716 61134 12768 61140
rect 12990 61160 12992 61169
rect 13044 61160 13046 61169
rect 12990 61095 13046 61104
rect 11060 61056 11112 61062
rect 11060 60998 11112 61004
rect 12164 61056 12216 61062
rect 12164 60998 12216 61004
rect 9036 60716 9088 60722
rect 9036 60658 9088 60664
rect 9220 60512 9272 60518
rect 9220 60454 9272 60460
rect 9232 44470 9260 60454
rect 10140 57860 10192 57866
rect 10140 57802 10192 57808
rect 10152 50386 10180 57802
rect 10784 52556 10836 52562
rect 10784 52498 10836 52504
rect 10140 50380 10192 50386
rect 10140 50322 10192 50328
rect 10796 47598 10824 52498
rect 10784 47592 10836 47598
rect 10784 47534 10836 47540
rect 10324 46980 10376 46986
rect 10324 46922 10376 46928
rect 9220 44464 9272 44470
rect 9220 44406 9272 44412
rect 9588 44260 9640 44266
rect 9588 44202 9640 44208
rect 9600 43858 9628 44202
rect 9588 43852 9640 43858
rect 9588 43794 9640 43800
rect 9036 37324 9088 37330
rect 9036 37266 9088 37272
rect 9048 37126 9076 37266
rect 9036 37120 9088 37126
rect 9036 37062 9088 37068
rect 10336 31210 10364 46922
rect 12176 33590 12204 60998
rect 13556 60790 13584 63294
rect 14094 63294 14320 63322
rect 14094 63200 14150 63294
rect 14292 60790 14320 63294
rect 14830 63294 14964 63322
rect 14830 63200 14886 63294
rect 14936 61198 14964 63294
rect 15566 63294 15792 63322
rect 15566 63200 15622 63294
rect 14924 61192 14976 61198
rect 14924 61134 14976 61140
rect 14648 61124 14700 61130
rect 14648 61066 14700 61072
rect 15200 61124 15252 61130
rect 15200 61066 15252 61072
rect 13544 60784 13596 60790
rect 13544 60726 13596 60732
rect 14280 60784 14332 60790
rect 14280 60726 14332 60732
rect 13636 60512 13688 60518
rect 13636 60454 13688 60460
rect 14372 60512 14424 60518
rect 14372 60454 14424 60460
rect 13648 60246 13676 60454
rect 13636 60240 13688 60246
rect 13636 60182 13688 60188
rect 14384 59770 14412 60454
rect 14372 59764 14424 59770
rect 14372 59706 14424 59712
rect 13084 49768 13136 49774
rect 13084 49710 13136 49716
rect 13096 39370 13124 49710
rect 13084 39364 13136 39370
rect 13084 39306 13136 39312
rect 13820 35284 13872 35290
rect 13820 35226 13872 35232
rect 12164 33584 12216 33590
rect 12164 33526 12216 33532
rect 10324 31204 10376 31210
rect 10324 31146 10376 31152
rect 13832 29714 13860 35226
rect 14660 31754 14688 61066
rect 15212 55214 15240 61066
rect 15764 60790 15792 63294
rect 16132 63294 16358 63322
rect 15844 61328 15896 61334
rect 15844 61270 15896 61276
rect 15856 60790 15884 61270
rect 16132 61198 16160 63294
rect 16302 63200 16358 63294
rect 17038 63322 17094 64000
rect 17774 63322 17830 64000
rect 18510 63322 18566 64000
rect 17038 63294 17264 63322
rect 17038 63200 17094 63294
rect 17236 61198 17264 63294
rect 17774 63294 17908 63322
rect 17774 63200 17830 63294
rect 16120 61192 16172 61198
rect 16120 61134 16172 61140
rect 17224 61192 17276 61198
rect 17880 61180 17908 63294
rect 18510 63294 18736 63322
rect 18510 63200 18566 63294
rect 18236 61328 18288 61334
rect 18236 61270 18288 61276
rect 17960 61192 18012 61198
rect 17880 61152 17960 61180
rect 17224 61134 17276 61140
rect 17960 61134 18012 61140
rect 17408 61124 17460 61130
rect 17408 61066 17460 61072
rect 17316 61056 17368 61062
rect 17316 60998 17368 61004
rect 15752 60784 15804 60790
rect 15752 60726 15804 60732
rect 15844 60784 15896 60790
rect 15844 60726 15896 60732
rect 15936 57316 15988 57322
rect 15936 57258 15988 57264
rect 15212 55186 15332 55214
rect 15200 45824 15252 45830
rect 15200 45766 15252 45772
rect 15212 45558 15240 45766
rect 15200 45552 15252 45558
rect 15200 45494 15252 45500
rect 15304 42129 15332 55186
rect 15290 42120 15346 42129
rect 15290 42055 15346 42064
rect 15752 36032 15804 36038
rect 15752 35974 15804 35980
rect 14660 31726 14780 31754
rect 13820 29708 13872 29714
rect 13820 29650 13872 29656
rect 9956 29640 10008 29646
rect 9956 29582 10008 29588
rect 9680 29096 9732 29102
rect 9680 29038 9732 29044
rect 8944 28552 8996 28558
rect 8944 28494 8996 28500
rect 9692 28490 9720 29038
rect 9680 28484 9732 28490
rect 9680 28426 9732 28432
rect 7840 26988 7892 26994
rect 7840 26930 7892 26936
rect 9692 25906 9720 28426
rect 9680 25900 9732 25906
rect 9680 25842 9732 25848
rect 9680 22636 9732 22642
rect 9680 22578 9732 22584
rect 9692 22234 9720 22578
rect 9680 22228 9732 22234
rect 9680 22170 9732 22176
rect 7288 22024 7340 22030
rect 7288 21966 7340 21972
rect 7300 21690 7328 21966
rect 7288 21684 7340 21690
rect 7288 21626 7340 21632
rect 7380 20460 7432 20466
rect 7380 20402 7432 20408
rect 8024 20460 8076 20466
rect 8024 20402 8076 20408
rect 7012 18692 7064 18698
rect 7012 18634 7064 18640
rect 7024 17134 7052 18634
rect 7104 18624 7156 18630
rect 7104 18566 7156 18572
rect 7116 18290 7144 18566
rect 7104 18284 7156 18290
rect 7104 18226 7156 18232
rect 7012 17128 7064 17134
rect 7012 17070 7064 17076
rect 6918 13288 6974 13297
rect 6918 13223 6974 13232
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 2872 11076 2924 11082
rect 2872 11018 2924 11024
rect 7392 10810 7420 20402
rect 7472 19712 7524 19718
rect 7472 19654 7524 19660
rect 7484 19446 7512 19654
rect 7472 19440 7524 19446
rect 7472 19382 7524 19388
rect 8036 17882 8064 20402
rect 9404 20256 9456 20262
rect 9404 20198 9456 20204
rect 9416 19990 9444 20198
rect 9404 19984 9456 19990
rect 9404 19926 9456 19932
rect 9312 19848 9364 19854
rect 9312 19790 9364 19796
rect 9220 19712 9272 19718
rect 9220 19654 9272 19660
rect 8208 18760 8260 18766
rect 8208 18702 8260 18708
rect 8116 18284 8168 18290
rect 8116 18226 8168 18232
rect 8024 17876 8076 17882
rect 8024 17818 8076 17824
rect 8128 17814 8156 18226
rect 8116 17808 8168 17814
rect 8116 17750 8168 17756
rect 8220 17202 8248 18702
rect 9128 17876 9180 17882
rect 9128 17818 9180 17824
rect 8208 17196 8260 17202
rect 8208 17138 8260 17144
rect 7564 16584 7616 16590
rect 7564 16526 7616 16532
rect 7576 16182 7604 16526
rect 7564 16176 7616 16182
rect 7564 16118 7616 16124
rect 8220 15178 8248 17138
rect 9140 16590 9168 17818
rect 9232 17678 9260 19654
rect 9220 17672 9272 17678
rect 9220 17614 9272 17620
rect 9128 16584 9180 16590
rect 9128 16526 9180 16532
rect 9324 16454 9352 19790
rect 9588 19780 9640 19786
rect 9588 19722 9640 19728
rect 9496 17808 9548 17814
rect 9496 17750 9548 17756
rect 9508 17678 9536 17750
rect 9496 17672 9548 17678
rect 9496 17614 9548 17620
rect 9404 17604 9456 17610
rect 9404 17546 9456 17552
rect 9416 16658 9444 17546
rect 9600 17542 9628 19722
rect 9680 18692 9732 18698
rect 9680 18634 9732 18640
rect 9692 17882 9720 18634
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9588 17536 9640 17542
rect 9588 17478 9640 17484
rect 9600 16998 9628 17478
rect 9784 17134 9812 18022
rect 9772 17128 9824 17134
rect 9772 17070 9824 17076
rect 9588 16992 9640 16998
rect 9588 16934 9640 16940
rect 9404 16652 9456 16658
rect 9404 16594 9456 16600
rect 9312 16448 9364 16454
rect 9312 16390 9364 16396
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 9876 15502 9904 15846
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 8220 15150 8340 15178
rect 8312 14482 8340 15150
rect 9772 15020 9824 15026
rect 9772 14962 9824 14968
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 9312 14476 9364 14482
rect 9312 14418 9364 14424
rect 9324 13938 9352 14418
rect 8852 13932 8904 13938
rect 8852 13874 8904 13880
rect 9312 13932 9364 13938
rect 9312 13874 9364 13880
rect 8864 12782 8892 13874
rect 9324 13394 9352 13874
rect 9692 13394 9720 14758
rect 9312 13388 9364 13394
rect 9312 13330 9364 13336
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 9784 12986 9812 14962
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 8852 12776 8904 12782
rect 8852 12718 8904 12724
rect 9496 12776 9548 12782
rect 9496 12718 9548 12724
rect 9508 11898 9536 12718
rect 9496 11892 9548 11898
rect 9496 11834 9548 11840
rect 8576 11076 8628 11082
rect 8576 11018 8628 11024
rect 7380 10804 7432 10810
rect 7380 10746 7432 10752
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 6826 10296 6882 10305
rect 6826 10231 6882 10240
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 1766 8055 1822 8064
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 6000 7880 6052 7886
rect 6000 7822 6052 7828
rect 1596 7478 1624 7822
rect 1860 7812 1912 7818
rect 1860 7754 1912 7760
rect 1584 7472 1636 7478
rect 1872 7449 1900 7754
rect 1584 7414 1636 7420
rect 1858 7440 1914 7449
rect 1858 7375 1914 7384
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 1858 6760 1914 6769
rect 1858 6695 1860 6704
rect 1912 6695 1914 6704
rect 1860 6666 1912 6672
rect 1768 6248 1820 6254
rect 1768 6190 1820 6196
rect 1780 6089 1808 6190
rect 1766 6080 1822 6089
rect 1766 6015 1822 6024
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 1860 5636 1912 5642
rect 1860 5578 1912 5584
rect 1872 5409 1900 5578
rect 1858 5400 1914 5409
rect 1858 5335 1914 5344
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 1596 4758 1624 5170
rect 1768 5160 1820 5166
rect 1768 5102 1820 5108
rect 1584 4752 1636 4758
rect 1780 4729 1808 5102
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 1584 4694 1636 4700
rect 1766 4720 1822 4729
rect 1766 4655 1822 4664
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 1768 4072 1820 4078
rect 1766 4040 1768 4049
rect 1820 4040 1822 4049
rect 1766 3975 1822 3984
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 1860 3460 1912 3466
rect 1860 3402 1912 3408
rect 1872 3369 1900 3402
rect 1858 3360 1914 3369
rect 1858 3295 1914 3304
rect 4632 3058 4660 4558
rect 5908 4140 5960 4146
rect 5908 4082 5960 4088
rect 5920 4049 5948 4082
rect 5906 4040 5962 4049
rect 5906 3975 5962 3984
rect 6012 3670 6040 7822
rect 6460 4208 6512 4214
rect 6460 4150 6512 4156
rect 6000 3664 6052 3670
rect 6000 3606 6052 3612
rect 6184 3528 6236 3534
rect 6184 3470 6236 3476
rect 5908 3120 5960 3126
rect 5908 3062 5960 3068
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 1768 2984 1820 2990
rect 1768 2926 1820 2932
rect 1780 2689 1808 2926
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 1766 2680 1822 2689
rect 4214 2683 4522 2692
rect 1766 2615 1822 2624
rect 1584 2440 1636 2446
rect 1584 2382 1636 2388
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 1596 2106 1624 2382
rect 1860 2372 1912 2378
rect 1860 2314 1912 2320
rect 1584 2100 1636 2106
rect 1584 2042 1636 2048
rect 1872 2009 1900 2314
rect 4436 2304 4488 2310
rect 4436 2246 4488 2252
rect 4448 2038 4476 2246
rect 4436 2032 4488 2038
rect 1858 2000 1914 2009
rect 4436 1974 4488 1980
rect 1858 1935 1914 1944
rect 4540 800 4568 2382
rect 5724 2372 5776 2378
rect 5724 2314 5776 2320
rect 5736 1426 5764 2314
rect 5724 1420 5776 1426
rect 5724 1362 5776 1368
rect 5920 800 5948 3062
rect 6196 800 6224 3470
rect 6472 800 6500 4150
rect 6840 4146 6868 10231
rect 7196 9444 7248 9450
rect 7196 9386 7248 9392
rect 7104 5024 7156 5030
rect 7104 4966 7156 4972
rect 6920 4548 6972 4554
rect 6920 4490 6972 4496
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6644 4004 6696 4010
rect 6644 3946 6696 3952
rect 6656 2825 6684 3946
rect 6642 2816 6698 2825
rect 6932 2774 6960 4490
rect 7012 4480 7064 4486
rect 7012 4422 7064 4428
rect 7024 4282 7052 4422
rect 7012 4276 7064 4282
rect 7012 4218 7064 4224
rect 7010 3768 7066 3777
rect 7010 3703 7012 3712
rect 7064 3703 7066 3712
rect 7012 3674 7064 3680
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 6642 2751 6698 2760
rect 6748 2746 6960 2774
rect 6748 800 6776 2746
rect 6920 2304 6972 2310
rect 6920 2246 6972 2252
rect 6932 1494 6960 2246
rect 6920 1488 6972 1494
rect 6920 1430 6972 1436
rect 7024 800 7052 3334
rect 7116 2854 7144 4966
rect 7104 2848 7156 2854
rect 7104 2790 7156 2796
rect 7208 2650 7236 9386
rect 8300 8968 8352 8974
rect 8298 8936 8300 8945
rect 8352 8936 8354 8945
rect 8298 8871 8354 8880
rect 7930 7984 7986 7993
rect 7930 7919 7986 7928
rect 7944 7886 7972 7919
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 8588 7818 8616 11018
rect 9496 10600 9548 10606
rect 9494 10568 9496 10577
rect 9680 10600 9732 10606
rect 9548 10568 9550 10577
rect 9680 10542 9732 10548
rect 9494 10503 9550 10512
rect 9692 9518 9720 10542
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 8772 7886 8800 9454
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 8576 7812 8628 7818
rect 8576 7754 8628 7760
rect 7380 7268 7432 7274
rect 7380 7210 7432 7216
rect 7288 4208 7340 4214
rect 7288 4150 7340 4156
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 7300 800 7328 4150
rect 7392 2854 7420 7210
rect 8772 6866 8800 7822
rect 9772 7812 9824 7818
rect 9772 7754 9824 7760
rect 9496 7404 9548 7410
rect 9496 7346 9548 7352
rect 9588 7404 9640 7410
rect 9588 7346 9640 7352
rect 9404 7200 9456 7206
rect 9404 7142 9456 7148
rect 8760 6860 8812 6866
rect 8760 6802 8812 6808
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 9140 6458 9168 6734
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 9312 6316 9364 6322
rect 9312 6258 9364 6264
rect 8944 6248 8996 6254
rect 8944 6190 8996 6196
rect 7932 5840 7984 5846
rect 7932 5782 7984 5788
rect 7748 5568 7800 5574
rect 7748 5510 7800 5516
rect 7564 4480 7616 4486
rect 7564 4422 7616 4428
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 7484 3738 7512 3878
rect 7472 3732 7524 3738
rect 7472 3674 7524 3680
rect 7576 3670 7604 4422
rect 7654 3904 7710 3913
rect 7654 3839 7710 3848
rect 7668 3670 7696 3839
rect 7564 3664 7616 3670
rect 7564 3606 7616 3612
rect 7656 3664 7708 3670
rect 7656 3606 7708 3612
rect 7564 2984 7616 2990
rect 7564 2926 7616 2932
rect 7380 2848 7432 2854
rect 7380 2790 7432 2796
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 7392 2378 7420 2586
rect 7380 2372 7432 2378
rect 7380 2314 7432 2320
rect 7472 2304 7524 2310
rect 7472 2246 7524 2252
rect 7484 1766 7512 2246
rect 7472 1760 7524 1766
rect 7472 1702 7524 1708
rect 7576 800 7604 2926
rect 7760 2774 7788 5510
rect 7944 2854 7972 5782
rect 8956 5302 8984 6190
rect 9140 5914 9168 6258
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 9324 5710 9352 6258
rect 9416 6236 9444 7142
rect 9508 6662 9536 7346
rect 9600 6798 9628 7346
rect 9784 7177 9812 7754
rect 9968 7750 9996 29582
rect 12808 28552 12860 28558
rect 12808 28494 12860 28500
rect 10692 25900 10744 25906
rect 10692 25842 10744 25848
rect 10704 23118 10732 25842
rect 12164 24132 12216 24138
rect 12164 24074 12216 24080
rect 12176 23322 12204 24074
rect 12820 23798 12848 28494
rect 13728 24132 13780 24138
rect 13728 24074 13780 24080
rect 12808 23792 12860 23798
rect 12808 23734 12860 23740
rect 12164 23316 12216 23322
rect 12164 23258 12216 23264
rect 12820 23118 12848 23734
rect 13740 23730 13768 24074
rect 13728 23724 13780 23730
rect 13728 23666 13780 23672
rect 10140 23112 10192 23118
rect 10140 23054 10192 23060
rect 10692 23112 10744 23118
rect 10692 23054 10744 23060
rect 10876 23112 10928 23118
rect 10876 23054 10928 23060
rect 12808 23112 12860 23118
rect 12808 23054 12860 23060
rect 10152 22098 10180 23054
rect 10888 22982 10916 23054
rect 10876 22976 10928 22982
rect 10876 22918 10928 22924
rect 10140 22094 10192 22098
rect 10140 22092 10364 22094
rect 10192 22066 10364 22092
rect 10140 22034 10192 22040
rect 10336 21554 10364 22066
rect 11060 22024 11112 22030
rect 11060 21966 11112 21972
rect 10324 21548 10376 21554
rect 10324 21490 10376 21496
rect 10048 19168 10100 19174
rect 10048 19110 10100 19116
rect 10060 17678 10088 19110
rect 10048 17672 10100 17678
rect 10048 17614 10100 17620
rect 10140 16108 10192 16114
rect 10140 16050 10192 16056
rect 10048 16040 10100 16046
rect 10048 15982 10100 15988
rect 10060 14074 10088 15982
rect 10048 14068 10100 14074
rect 10048 14010 10100 14016
rect 10152 12442 10180 16050
rect 10232 15360 10284 15366
rect 10232 15302 10284 15308
rect 10244 14482 10272 15302
rect 10232 14476 10284 14482
rect 10232 14418 10284 14424
rect 10140 12436 10192 12442
rect 10140 12378 10192 12384
rect 10336 12306 10364 21490
rect 11072 21321 11100 21966
rect 12716 21548 12768 21554
rect 12716 21490 12768 21496
rect 13268 21548 13320 21554
rect 13268 21490 13320 21496
rect 11058 21312 11114 21321
rect 11058 21247 11114 21256
rect 12728 21078 12756 21490
rect 12900 21480 12952 21486
rect 12900 21422 12952 21428
rect 13176 21480 13228 21486
rect 13176 21422 13228 21428
rect 12808 21344 12860 21350
rect 12808 21286 12860 21292
rect 12716 21072 12768 21078
rect 12716 21014 12768 21020
rect 11704 21004 11756 21010
rect 11704 20946 11756 20952
rect 12256 21004 12308 21010
rect 12256 20946 12308 20952
rect 11152 20800 11204 20806
rect 11152 20742 11204 20748
rect 11164 20466 11192 20742
rect 11716 20534 11744 20946
rect 11704 20528 11756 20534
rect 11704 20470 11756 20476
rect 11152 20460 11204 20466
rect 11152 20402 11204 20408
rect 11888 20392 11940 20398
rect 11888 20334 11940 20340
rect 11060 20256 11112 20262
rect 11060 20198 11112 20204
rect 10692 19712 10744 19718
rect 10692 19654 10744 19660
rect 10704 19378 10732 19654
rect 10692 19372 10744 19378
rect 10692 19314 10744 19320
rect 11072 18222 11100 20198
rect 11900 19378 11928 20334
rect 11888 19372 11940 19378
rect 11888 19314 11940 19320
rect 12164 19304 12216 19310
rect 12164 19246 12216 19252
rect 12176 18970 12204 19246
rect 12164 18964 12216 18970
rect 12164 18906 12216 18912
rect 12268 18290 12296 20946
rect 12716 20936 12768 20942
rect 12716 20878 12768 20884
rect 12348 18692 12400 18698
rect 12348 18634 12400 18640
rect 12256 18284 12308 18290
rect 12256 18226 12308 18232
rect 11060 18216 11112 18222
rect 11060 18158 11112 18164
rect 11888 16108 11940 16114
rect 11888 16050 11940 16056
rect 11612 15496 11664 15502
rect 11612 15438 11664 15444
rect 11152 14408 11204 14414
rect 11152 14350 11204 14356
rect 11164 12986 11192 14350
rect 11428 13320 11480 13326
rect 11428 13262 11480 13268
rect 11244 13184 11296 13190
rect 11244 13126 11296 13132
rect 11152 12980 11204 12986
rect 11152 12922 11204 12928
rect 11256 12714 11284 13126
rect 11244 12708 11296 12714
rect 11244 12650 11296 12656
rect 11440 12442 11468 13262
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 10324 12300 10376 12306
rect 10324 12242 10376 12248
rect 10336 11558 10364 12242
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 10520 11762 10548 12174
rect 11060 12164 11112 12170
rect 11060 12106 11112 12112
rect 11072 11830 11100 12106
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 11060 11824 11112 11830
rect 11060 11766 11112 11772
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 11152 10532 11204 10538
rect 11152 10474 11204 10480
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10600 8492 10652 8498
rect 10600 8434 10652 8440
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 10060 7886 10088 8026
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 9956 7744 10008 7750
rect 9956 7686 10008 7692
rect 9770 7168 9826 7177
rect 9770 7103 9826 7112
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9496 6248 9548 6254
rect 9416 6208 9496 6236
rect 9496 6190 9548 6196
rect 9588 6248 9640 6254
rect 9588 6190 9640 6196
rect 9404 6112 9456 6118
rect 9404 6054 9456 6060
rect 9416 5778 9444 6054
rect 9600 5794 9628 6190
rect 9404 5772 9456 5778
rect 9404 5714 9456 5720
rect 9508 5766 9628 5794
rect 9692 5778 9720 6598
rect 9680 5772 9732 5778
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 8944 5296 8996 5302
rect 8944 5238 8996 5244
rect 8116 5228 8168 5234
rect 8116 5170 8168 5176
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 8036 2854 8064 3130
rect 7932 2848 7984 2854
rect 7932 2790 7984 2796
rect 8024 2848 8076 2854
rect 8024 2790 8076 2796
rect 7668 2746 7788 2774
rect 7668 2582 7696 2746
rect 7656 2576 7708 2582
rect 7656 2518 7708 2524
rect 7840 2508 7892 2514
rect 7840 2450 7892 2456
rect 7656 2372 7708 2378
rect 7656 2314 7708 2320
rect 7668 1902 7696 2314
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 7656 1896 7708 1902
rect 7656 1838 7708 1844
rect 7760 1834 7788 2246
rect 7748 1828 7800 1834
rect 7748 1770 7800 1776
rect 7852 800 7880 2450
rect 8128 800 8156 5170
rect 8760 5092 8812 5098
rect 8760 5034 8812 5040
rect 8300 4548 8352 4554
rect 8300 4490 8352 4496
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 8220 3466 8248 4082
rect 8208 3460 8260 3466
rect 8208 3402 8260 3408
rect 8208 2984 8260 2990
rect 8206 2952 8208 2961
rect 8260 2952 8262 2961
rect 8206 2887 8262 2896
rect 8312 2774 8340 4490
rect 8484 4208 8536 4214
rect 8484 4150 8536 4156
rect 8496 3466 8524 4150
rect 8574 4040 8630 4049
rect 8574 3975 8630 3984
rect 8668 4004 8720 4010
rect 8588 3942 8616 3975
rect 8668 3946 8720 3952
rect 8576 3936 8628 3942
rect 8576 3878 8628 3884
rect 8392 3460 8444 3466
rect 8392 3402 8444 3408
rect 8484 3460 8536 3466
rect 8484 3402 8536 3408
rect 8404 2990 8432 3402
rect 8576 3392 8628 3398
rect 8576 3334 8628 3340
rect 8392 2984 8444 2990
rect 8392 2926 8444 2932
rect 8312 2746 8432 2774
rect 8404 800 8432 2746
rect 8484 2304 8536 2310
rect 8484 2246 8536 2252
rect 8496 1970 8524 2246
rect 8484 1964 8536 1970
rect 8484 1906 8536 1912
rect 8588 1442 8616 3334
rect 8680 2038 8708 3946
rect 8772 2922 8800 5034
rect 8852 4548 8904 4554
rect 8852 4490 8904 4496
rect 8864 3670 8892 4490
rect 9508 4146 9536 5766
rect 9680 5714 9732 5720
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 9600 5370 9628 5646
rect 9588 5364 9640 5370
rect 9588 5306 9640 5312
rect 9588 5228 9640 5234
rect 9588 5170 9640 5176
rect 9600 4214 9628 5170
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9692 4690 9720 4966
rect 9784 4690 9812 7103
rect 10060 5234 10088 7822
rect 10612 7546 10640 8434
rect 10600 7540 10652 7546
rect 10600 7482 10652 7488
rect 10704 7342 10732 8978
rect 10784 7472 10836 7478
rect 10784 7414 10836 7420
rect 10692 7336 10744 7342
rect 10692 7278 10744 7284
rect 10704 6798 10732 7278
rect 10796 6866 10824 7414
rect 10876 7336 10928 7342
rect 10876 7278 10928 7284
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 10888 7002 10916 7278
rect 10876 6996 10928 7002
rect 10876 6938 10928 6944
rect 10784 6860 10836 6866
rect 10784 6802 10836 6808
rect 10876 6860 10928 6866
rect 10876 6802 10928 6808
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10888 6390 10916 6802
rect 10876 6384 10928 6390
rect 10876 6326 10928 6332
rect 11072 5914 11100 7278
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 10140 5636 10192 5642
rect 10140 5578 10192 5584
rect 10416 5636 10468 5642
rect 10416 5578 10468 5584
rect 10152 5370 10180 5578
rect 10140 5364 10192 5370
rect 10140 5306 10192 5312
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 10428 5216 10456 5578
rect 10508 5228 10560 5234
rect 10428 5188 10508 5216
rect 9876 4826 10088 4842
rect 9864 4820 10088 4826
rect 9916 4814 10088 4820
rect 9864 4762 9916 4768
rect 10060 4758 10088 4814
rect 10048 4752 10100 4758
rect 9862 4720 9918 4729
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9772 4684 9824 4690
rect 10048 4694 10100 4700
rect 10428 4690 10456 5188
rect 10508 5170 10560 5176
rect 10600 5160 10652 5166
rect 10600 5102 10652 5108
rect 9862 4655 9918 4664
rect 9956 4684 10008 4690
rect 9772 4626 9824 4632
rect 9876 4622 9904 4655
rect 9956 4626 10008 4632
rect 10416 4684 10468 4690
rect 10416 4626 10468 4632
rect 9864 4616 9916 4622
rect 9864 4558 9916 4564
rect 9772 4480 9824 4486
rect 9772 4422 9824 4428
rect 9588 4208 9640 4214
rect 9588 4150 9640 4156
rect 9496 4140 9548 4146
rect 9496 4082 9548 4088
rect 9600 4078 9628 4150
rect 8944 4072 8996 4078
rect 8944 4014 8996 4020
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 9404 4072 9456 4078
rect 9404 4014 9456 4020
rect 9588 4072 9640 4078
rect 9588 4014 9640 4020
rect 8852 3664 8904 3670
rect 8852 3606 8904 3612
rect 8852 3460 8904 3466
rect 8852 3402 8904 3408
rect 8760 2916 8812 2922
rect 8760 2858 8812 2864
rect 8668 2032 8720 2038
rect 8668 1974 8720 1980
rect 8864 1442 8892 3402
rect 8956 2553 8984 4014
rect 9036 3936 9088 3942
rect 9036 3878 9088 3884
rect 9048 2650 9076 3878
rect 9232 3398 9260 4014
rect 9416 3913 9444 4014
rect 9402 3904 9458 3913
rect 9402 3839 9458 3848
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9220 3392 9272 3398
rect 9220 3334 9272 3340
rect 9128 3120 9180 3126
rect 9600 3097 9628 3470
rect 9128 3062 9180 3068
rect 9586 3088 9642 3097
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 8942 2544 8998 2553
rect 8942 2479 8998 2488
rect 9140 1442 9168 3062
rect 9220 3052 9272 3058
rect 9586 3023 9588 3032
rect 9220 2994 9272 3000
rect 9640 3023 9642 3032
rect 9588 2994 9640 3000
rect 9232 2310 9260 2994
rect 9588 2916 9640 2922
rect 9588 2858 9640 2864
rect 9600 2774 9628 2858
rect 9324 2746 9628 2774
rect 9324 2514 9352 2746
rect 9312 2508 9364 2514
rect 9312 2450 9364 2456
rect 9496 2372 9548 2378
rect 9496 2314 9548 2320
rect 9220 2304 9272 2310
rect 9220 2246 9272 2252
rect 9508 2038 9536 2314
rect 9496 2032 9548 2038
rect 9496 1974 9548 1980
rect 8588 1414 8708 1442
rect 8864 1414 8984 1442
rect 9140 1414 9260 1442
rect 8680 800 8708 1414
rect 8956 800 8984 1414
rect 9232 800 9260 1414
rect 9496 1420 9548 1426
rect 9496 1362 9548 1368
rect 9508 800 9536 1362
rect 9784 800 9812 4422
rect 9864 3528 9916 3534
rect 9864 3470 9916 3476
rect 9876 3194 9904 3470
rect 9968 3466 9996 4626
rect 10324 4072 10376 4078
rect 10324 4014 10376 4020
rect 10048 4004 10100 4010
rect 10048 3946 10100 3952
rect 9956 3460 10008 3466
rect 9956 3402 10008 3408
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9968 2990 9996 3402
rect 10060 3058 10088 3946
rect 10336 3534 10364 4014
rect 10612 3738 10640 5102
rect 11164 4146 11192 10474
rect 11256 9654 11284 12038
rect 11624 11506 11652 15438
rect 11900 15366 11928 16050
rect 12256 15904 12308 15910
rect 12256 15846 12308 15852
rect 11888 15360 11940 15366
rect 11888 15302 11940 15308
rect 12268 15026 12296 15846
rect 12256 15020 12308 15026
rect 12256 14962 12308 14968
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 11992 13938 12020 14214
rect 11980 13932 12032 13938
rect 11980 13874 12032 13880
rect 11886 13016 11942 13025
rect 11886 12951 11942 12960
rect 11900 12918 11928 12951
rect 11888 12912 11940 12918
rect 11888 12854 11940 12860
rect 11980 12912 12032 12918
rect 11980 12854 12032 12860
rect 11900 12170 11928 12854
rect 11992 12442 12020 12854
rect 12072 12844 12124 12850
rect 12072 12786 12124 12792
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 12084 12238 12112 12786
rect 12256 12436 12308 12442
rect 12256 12378 12308 12384
rect 12072 12232 12124 12238
rect 12070 12200 12072 12209
rect 12124 12200 12126 12209
rect 11888 12164 11940 12170
rect 12070 12135 12126 12144
rect 11888 12106 11940 12112
rect 12084 12109 12112 12135
rect 12268 11830 12296 12378
rect 12256 11824 12308 11830
rect 11886 11792 11942 11801
rect 12256 11766 12308 11772
rect 11886 11727 11888 11736
rect 11940 11727 11942 11736
rect 11888 11698 11940 11704
rect 11796 11620 11848 11626
rect 11796 11562 11848 11568
rect 11808 11506 11836 11562
rect 11624 11478 11836 11506
rect 11716 11218 11744 11478
rect 11900 11354 11928 11698
rect 12164 11688 12216 11694
rect 12164 11630 12216 11636
rect 11888 11348 11940 11354
rect 11888 11290 11940 11296
rect 11704 11212 11756 11218
rect 11704 11154 11756 11160
rect 11428 11144 11480 11150
rect 11428 11086 11480 11092
rect 11440 10266 11468 11086
rect 11716 10606 11744 11154
rect 12176 10810 12204 11630
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 12268 10606 12296 11766
rect 12360 11762 12388 18634
rect 12728 18358 12756 20878
rect 12820 19854 12848 21286
rect 12912 20806 12940 21422
rect 13188 21010 13216 21422
rect 13176 21004 13228 21010
rect 13176 20946 13228 20952
rect 13280 20874 13308 21490
rect 13636 21004 13688 21010
rect 13636 20946 13688 20952
rect 13268 20868 13320 20874
rect 13268 20810 13320 20816
rect 12900 20800 12952 20806
rect 12900 20742 12952 20748
rect 13084 20800 13136 20806
rect 13084 20742 13136 20748
rect 12912 20602 12940 20742
rect 12900 20596 12952 20602
rect 12900 20538 12952 20544
rect 12808 19848 12860 19854
rect 12808 19790 12860 19796
rect 12716 18352 12768 18358
rect 12716 18294 12768 18300
rect 12532 18148 12584 18154
rect 12532 18090 12584 18096
rect 12544 17202 12572 18090
rect 12992 17808 13044 17814
rect 13096 17796 13124 20742
rect 13360 20460 13412 20466
rect 13360 20402 13412 20408
rect 13176 19916 13228 19922
rect 13176 19858 13228 19864
rect 13188 17814 13216 19858
rect 13372 17882 13400 20402
rect 13648 20330 13676 20946
rect 13636 20324 13688 20330
rect 13636 20266 13688 20272
rect 13636 20052 13688 20058
rect 13636 19994 13688 20000
rect 13452 18080 13504 18086
rect 13452 18022 13504 18028
rect 13360 17876 13412 17882
rect 13360 17818 13412 17824
rect 13044 17768 13124 17796
rect 12992 17750 13044 17756
rect 13096 17678 13124 17768
rect 13176 17808 13228 17814
rect 13176 17750 13228 17756
rect 13084 17672 13136 17678
rect 13084 17614 13136 17620
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 12808 16584 12860 16590
rect 12808 16526 12860 16532
rect 13360 16584 13412 16590
rect 13360 16526 13412 16532
rect 12624 16040 12676 16046
rect 12624 15982 12676 15988
rect 12636 15026 12664 15982
rect 12716 15428 12768 15434
rect 12716 15370 12768 15376
rect 12624 15020 12676 15026
rect 12624 14962 12676 14968
rect 12440 14340 12492 14346
rect 12440 14282 12492 14288
rect 12452 12434 12480 14282
rect 12636 12850 12664 14962
rect 12624 12844 12676 12850
rect 12624 12786 12676 12792
rect 12728 12434 12756 15370
rect 12452 12406 12572 12434
rect 12544 12238 12572 12406
rect 12636 12406 12756 12434
rect 12532 12232 12584 12238
rect 12532 12174 12584 12180
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 11704 10600 11756 10606
rect 11704 10542 11756 10548
rect 12256 10600 12308 10606
rect 12256 10542 12308 10548
rect 11428 10260 11480 10266
rect 11428 10202 11480 10208
rect 11336 10192 11388 10198
rect 11336 10134 11388 10140
rect 11244 9648 11296 9654
rect 11244 9590 11296 9596
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 11256 4826 11284 6734
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 11244 4004 11296 4010
rect 11244 3946 11296 3952
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 10600 3732 10652 3738
rect 10600 3674 10652 3680
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 10336 3126 10364 3470
rect 10324 3120 10376 3126
rect 10324 3062 10376 3068
rect 10048 3052 10100 3058
rect 10048 2994 10100 3000
rect 9956 2984 10008 2990
rect 9956 2926 10008 2932
rect 10322 2952 10378 2961
rect 10322 2887 10378 2896
rect 10600 2916 10652 2922
rect 10048 1488 10100 1494
rect 10048 1430 10100 1436
rect 10060 800 10088 1430
rect 10336 800 10364 2887
rect 10600 2858 10652 2864
rect 10612 800 10640 2858
rect 11060 2576 11112 2582
rect 11164 2564 11192 3878
rect 11256 2650 11284 3946
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 11112 2536 11192 2564
rect 11060 2518 11112 2524
rect 10876 2304 10928 2310
rect 10876 2246 10928 2252
rect 10888 800 10916 2246
rect 11348 1970 11376 10134
rect 11716 9994 11744 10542
rect 12164 10464 12216 10470
rect 12164 10406 12216 10412
rect 11704 9988 11756 9994
rect 11704 9930 11756 9936
rect 11428 7404 11480 7410
rect 11428 7346 11480 7352
rect 11440 6730 11468 7346
rect 11428 6724 11480 6730
rect 11428 6666 11480 6672
rect 11716 6390 11744 9930
rect 11704 6384 11756 6390
rect 11704 6326 11756 6332
rect 11888 5840 11940 5846
rect 11888 5782 11940 5788
rect 11796 4548 11848 4554
rect 11796 4490 11848 4496
rect 11704 4208 11756 4214
rect 11704 4150 11756 4156
rect 11428 2372 11480 2378
rect 11428 2314 11480 2320
rect 11336 1964 11388 1970
rect 11336 1906 11388 1912
rect 11152 1896 11204 1902
rect 11152 1838 11204 1844
rect 11164 800 11192 1838
rect 11440 800 11468 2314
rect 11716 800 11744 4150
rect 11808 2990 11836 4490
rect 11900 3670 11928 5782
rect 11980 5228 12032 5234
rect 11980 5170 12032 5176
rect 11888 3664 11940 3670
rect 11888 3606 11940 3612
rect 11796 2984 11848 2990
rect 11796 2926 11848 2932
rect 11796 2848 11848 2854
rect 11796 2790 11848 2796
rect 11808 2446 11836 2790
rect 11796 2440 11848 2446
rect 11796 2382 11848 2388
rect 11992 800 12020 5170
rect 12072 4752 12124 4758
rect 12072 4694 12124 4700
rect 12084 4146 12112 4694
rect 12072 4140 12124 4146
rect 12072 4082 12124 4088
rect 12176 3210 12204 10406
rect 12440 8900 12492 8906
rect 12440 8842 12492 8848
rect 12452 7818 12480 8842
rect 12440 7812 12492 7818
rect 12440 7754 12492 7760
rect 12452 7342 12480 7754
rect 12544 7585 12572 12174
rect 12530 7576 12586 7585
rect 12530 7511 12586 7520
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 12452 6186 12480 7278
rect 12440 6180 12492 6186
rect 12440 6122 12492 6128
rect 12440 4208 12492 4214
rect 12440 4150 12492 4156
rect 12348 4072 12400 4078
rect 12348 4014 12400 4020
rect 12360 3466 12388 4014
rect 12348 3460 12400 3466
rect 12348 3402 12400 3408
rect 12176 3182 12388 3210
rect 12256 2984 12308 2990
rect 12256 2926 12308 2932
rect 12268 800 12296 2926
rect 12360 2446 12388 3182
rect 12348 2440 12400 2446
rect 12348 2382 12400 2388
rect 12452 2122 12480 4150
rect 12544 3913 12572 7511
rect 12636 5914 12664 12406
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 12728 9382 12756 10610
rect 12716 9376 12768 9382
rect 12716 9318 12768 9324
rect 12716 8016 12768 8022
rect 12716 7958 12768 7964
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 12530 3904 12586 3913
rect 12530 3839 12586 3848
rect 12624 3664 12676 3670
rect 12624 3606 12676 3612
rect 12532 3596 12584 3602
rect 12532 3538 12584 3544
rect 12544 3398 12572 3538
rect 12532 3392 12584 3398
rect 12532 3334 12584 3340
rect 12636 2582 12664 3606
rect 12624 2576 12676 2582
rect 12624 2518 12676 2524
rect 12452 2094 12572 2122
rect 12544 800 12572 2094
rect 12728 1834 12756 7958
rect 12820 3754 12848 16526
rect 12900 16516 12952 16522
rect 12900 16458 12952 16464
rect 12912 15162 12940 16458
rect 13084 16176 13136 16182
rect 13084 16118 13136 16124
rect 13096 15706 13124 16118
rect 13372 15910 13400 16526
rect 13464 16114 13492 18022
rect 13648 16250 13676 19994
rect 14648 19848 14700 19854
rect 14648 19790 14700 19796
rect 14660 19310 14688 19790
rect 14648 19304 14700 19310
rect 14568 19264 14648 19292
rect 14568 18766 14596 19264
rect 14648 19246 14700 19252
rect 13728 18760 13780 18766
rect 13728 18702 13780 18708
rect 14556 18760 14608 18766
rect 14556 18702 14608 18708
rect 13740 17338 13768 18702
rect 13728 17332 13780 17338
rect 13728 17274 13780 17280
rect 14280 16788 14332 16794
rect 14280 16730 14332 16736
rect 14292 16590 14320 16730
rect 13728 16584 13780 16590
rect 13728 16526 13780 16532
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 13636 16244 13688 16250
rect 13636 16186 13688 16192
rect 13740 16114 13768 16526
rect 14292 16182 14320 16526
rect 14280 16176 14332 16182
rect 14280 16118 14332 16124
rect 13452 16108 13504 16114
rect 13452 16050 13504 16056
rect 13728 16108 13780 16114
rect 13728 16050 13780 16056
rect 13360 15904 13412 15910
rect 13360 15846 13412 15852
rect 13084 15700 13136 15706
rect 13084 15642 13136 15648
rect 13372 15570 13400 15846
rect 13740 15570 13768 16050
rect 14292 15570 14320 16118
rect 13360 15564 13412 15570
rect 13360 15506 13412 15512
rect 13728 15564 13780 15570
rect 13728 15506 13780 15512
rect 14280 15564 14332 15570
rect 14280 15506 14332 15512
rect 14648 15564 14700 15570
rect 14648 15506 14700 15512
rect 12900 15156 12952 15162
rect 12900 15098 12952 15104
rect 14292 14482 14320 15506
rect 14556 15088 14608 15094
rect 14556 15030 14608 15036
rect 14568 14618 14596 15030
rect 14556 14612 14608 14618
rect 14556 14554 14608 14560
rect 14280 14476 14332 14482
rect 14280 14418 14332 14424
rect 14292 14006 14320 14418
rect 14280 14000 14332 14006
rect 14280 13942 14332 13948
rect 13728 13932 13780 13938
rect 13728 13874 13780 13880
rect 13544 13320 13596 13326
rect 13544 13262 13596 13268
rect 13556 12986 13584 13262
rect 13544 12980 13596 12986
rect 13544 12922 13596 12928
rect 13084 12776 13136 12782
rect 13084 12718 13136 12724
rect 13096 12442 13124 12718
rect 13084 12436 13136 12442
rect 13084 12378 13136 12384
rect 13740 12374 13768 13874
rect 14292 13394 14320 13942
rect 14280 13388 14332 13394
rect 14280 13330 14332 13336
rect 14004 12844 14056 12850
rect 14004 12786 14056 12792
rect 13728 12368 13780 12374
rect 13728 12310 13780 12316
rect 14016 11898 14044 12786
rect 14004 11892 14056 11898
rect 14004 11834 14056 11840
rect 13268 11824 13320 11830
rect 13268 11766 13320 11772
rect 13636 11824 13688 11830
rect 13636 11766 13688 11772
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 13188 11218 13216 11494
rect 13176 11212 13228 11218
rect 13176 11154 13228 11160
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 12912 9994 12940 10610
rect 13188 10538 13216 11154
rect 13176 10532 13228 10538
rect 13176 10474 13228 10480
rect 13188 10198 13216 10474
rect 13176 10192 13228 10198
rect 13176 10134 13228 10140
rect 12900 9988 12952 9994
rect 12900 9930 12952 9936
rect 13280 9518 13308 11766
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 13372 10674 13400 11494
rect 13360 10668 13412 10674
rect 13360 10610 13412 10616
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13360 9988 13412 9994
rect 13360 9930 13412 9936
rect 13372 9586 13400 9930
rect 13464 9586 13492 9998
rect 13544 9648 13596 9654
rect 13544 9590 13596 9596
rect 13360 9580 13412 9586
rect 13360 9522 13412 9528
rect 13452 9580 13504 9586
rect 13452 9522 13504 9528
rect 13268 9512 13320 9518
rect 13268 9454 13320 9460
rect 13176 9376 13228 9382
rect 13176 9318 13228 9324
rect 12898 8800 12954 8809
rect 12898 8735 12954 8744
rect 12912 4078 12940 8735
rect 12992 4616 13044 4622
rect 12992 4558 13044 4564
rect 12900 4072 12952 4078
rect 12900 4014 12952 4020
rect 13004 4010 13032 4558
rect 13084 4548 13136 4554
rect 13084 4490 13136 4496
rect 12992 4004 13044 4010
rect 12992 3946 13044 3952
rect 12990 3904 13046 3913
rect 12990 3839 13046 3848
rect 12820 3738 12940 3754
rect 12820 3732 12952 3738
rect 12820 3726 12900 3732
rect 12900 3674 12952 3680
rect 12898 3496 12954 3505
rect 12898 3431 12954 3440
rect 12808 3392 12860 3398
rect 12808 3334 12860 3340
rect 12820 3058 12848 3334
rect 12912 3194 12940 3431
rect 12900 3188 12952 3194
rect 12900 3130 12952 3136
rect 12808 3052 12860 3058
rect 12808 2994 12860 3000
rect 13004 2446 13032 3839
rect 12992 2440 13044 2446
rect 12992 2382 13044 2388
rect 12808 2032 12860 2038
rect 12808 1974 12860 1980
rect 12716 1828 12768 1834
rect 12716 1770 12768 1776
rect 12820 800 12848 1974
rect 13096 800 13124 4490
rect 13188 1834 13216 9318
rect 13268 9104 13320 9110
rect 13268 9046 13320 9052
rect 13176 1828 13228 1834
rect 13176 1770 13228 1776
rect 13280 1766 13308 9046
rect 13372 8362 13400 9522
rect 13464 8838 13492 9522
rect 13556 9042 13584 9590
rect 13648 9382 13676 11766
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 13648 8906 13676 9318
rect 13832 9178 13860 10202
rect 14188 9920 14240 9926
rect 14188 9862 14240 9868
rect 14200 9586 14228 9862
rect 14188 9580 14240 9586
rect 14188 9522 14240 9528
rect 14280 9512 14332 9518
rect 14280 9454 14332 9460
rect 13820 9172 13872 9178
rect 13820 9114 13872 9120
rect 14292 8974 14320 9454
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 13636 8900 13688 8906
rect 13636 8842 13688 8848
rect 13452 8832 13504 8838
rect 13452 8774 13504 8780
rect 13464 8634 13492 8774
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 14004 8492 14056 8498
rect 14004 8434 14056 8440
rect 13360 8356 13412 8362
rect 13360 8298 13412 8304
rect 14016 8022 14044 8434
rect 14004 8016 14056 8022
rect 14004 7958 14056 7964
rect 13728 6180 13780 6186
rect 13728 6122 13780 6128
rect 13740 5234 13768 6122
rect 14462 5944 14518 5953
rect 13820 5908 13872 5914
rect 14462 5879 14518 5888
rect 13820 5850 13872 5856
rect 13728 5228 13780 5234
rect 13728 5170 13780 5176
rect 13832 5166 13860 5850
rect 14280 5636 14332 5642
rect 14280 5578 14332 5584
rect 13912 5568 13964 5574
rect 13912 5510 13964 5516
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 13544 3664 13596 3670
rect 13544 3606 13596 3612
rect 13740 3618 13768 4762
rect 13820 3664 13872 3670
rect 13740 3612 13820 3618
rect 13740 3606 13872 3612
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 13268 1760 13320 1766
rect 13268 1702 13320 1708
rect 13372 800 13400 3470
rect 13556 3398 13584 3606
rect 13740 3590 13860 3606
rect 13544 3392 13596 3398
rect 13544 3334 13596 3340
rect 13636 3052 13688 3058
rect 13924 3040 13952 5510
rect 14292 5370 14320 5578
rect 14280 5364 14332 5370
rect 14280 5306 14332 5312
rect 14292 4622 14320 5306
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14292 4214 14320 4558
rect 14280 4208 14332 4214
rect 14280 4150 14332 4156
rect 14188 3460 14240 3466
rect 14188 3402 14240 3408
rect 13688 3012 13952 3040
rect 13636 2994 13688 3000
rect 13912 2848 13964 2854
rect 13912 2790 13964 2796
rect 14004 2848 14056 2854
rect 14004 2790 14056 2796
rect 13636 2508 13688 2514
rect 13636 2450 13688 2456
rect 13648 800 13676 2450
rect 13924 800 13952 2790
rect 14016 2650 14044 2790
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 14200 800 14228 3402
rect 14476 3058 14504 5879
rect 14660 3738 14688 15506
rect 14752 15094 14780 31726
rect 15108 30320 15160 30326
rect 15108 30262 15160 30268
rect 15120 29170 15148 30262
rect 15108 29164 15160 29170
rect 15108 29106 15160 29112
rect 14924 20052 14976 20058
rect 14924 19994 14976 20000
rect 14832 17876 14884 17882
rect 14832 17818 14884 17824
rect 14844 17678 14872 17818
rect 14832 17672 14884 17678
rect 14832 17614 14884 17620
rect 14936 15910 14964 19994
rect 15016 16992 15068 16998
rect 15016 16934 15068 16940
rect 15028 16522 15056 16934
rect 15016 16516 15068 16522
rect 15016 16458 15068 16464
rect 14924 15904 14976 15910
rect 14924 15846 14976 15852
rect 14740 15088 14792 15094
rect 14740 15030 14792 15036
rect 15120 13433 15148 29106
rect 15384 21888 15436 21894
rect 15384 21830 15436 21836
rect 15292 21344 15344 21350
rect 15292 21286 15344 21292
rect 15200 20256 15252 20262
rect 15200 20198 15252 20204
rect 15212 19854 15240 20198
rect 15200 19848 15252 19854
rect 15200 19790 15252 19796
rect 15304 19378 15332 21286
rect 15396 20942 15424 21830
rect 15384 20936 15436 20942
rect 15384 20878 15436 20884
rect 15568 20936 15620 20942
rect 15568 20878 15620 20884
rect 15384 20800 15436 20806
rect 15384 20742 15436 20748
rect 15396 20466 15424 20742
rect 15384 20460 15436 20466
rect 15384 20402 15436 20408
rect 15292 19372 15344 19378
rect 15292 19314 15344 19320
rect 15200 19168 15252 19174
rect 15200 19110 15252 19116
rect 15212 18766 15240 19110
rect 15200 18760 15252 18766
rect 15200 18702 15252 18708
rect 15580 17882 15608 20878
rect 15568 17876 15620 17882
rect 15568 17818 15620 17824
rect 15384 17536 15436 17542
rect 15384 17478 15436 17484
rect 15396 17338 15424 17478
rect 15384 17332 15436 17338
rect 15384 17274 15436 17280
rect 15382 16144 15438 16153
rect 15382 16079 15384 16088
rect 15436 16079 15438 16088
rect 15384 16050 15436 16056
rect 15568 16040 15620 16046
rect 15568 15982 15620 15988
rect 15580 15570 15608 15982
rect 15568 15564 15620 15570
rect 15568 15506 15620 15512
rect 15200 15496 15252 15502
rect 15200 15438 15252 15444
rect 15212 13870 15240 15438
rect 15660 14884 15712 14890
rect 15660 14826 15712 14832
rect 15672 14482 15700 14826
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 15384 14408 15436 14414
rect 15384 14350 15436 14356
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 15106 13424 15162 13433
rect 15106 13359 15162 13368
rect 15016 12640 15068 12646
rect 15016 12582 15068 12588
rect 14924 12300 14976 12306
rect 14924 12242 14976 12248
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14752 11665 14780 12038
rect 14936 11762 14964 12242
rect 14924 11756 14976 11762
rect 14924 11698 14976 11704
rect 14832 11688 14884 11694
rect 14738 11656 14794 11665
rect 14832 11630 14884 11636
rect 14738 11591 14794 11600
rect 14844 11529 14872 11630
rect 14830 11520 14886 11529
rect 14830 11455 14886 11464
rect 14830 11248 14886 11257
rect 14830 11183 14832 11192
rect 14884 11183 14886 11192
rect 14832 11154 14884 11160
rect 15028 11150 15056 12582
rect 15016 11144 15068 11150
rect 15016 11086 15068 11092
rect 15120 10130 15148 13359
rect 15396 12986 15424 14350
rect 15660 14272 15712 14278
rect 15660 14214 15712 14220
rect 15568 13184 15620 13190
rect 15568 13126 15620 13132
rect 15384 12980 15436 12986
rect 15384 12922 15436 12928
rect 15200 12912 15252 12918
rect 15200 12854 15252 12860
rect 15212 10538 15240 12854
rect 15384 12232 15436 12238
rect 15384 12174 15436 12180
rect 15292 11688 15344 11694
rect 15290 11656 15292 11665
rect 15344 11656 15346 11665
rect 15290 11591 15346 11600
rect 15292 10668 15344 10674
rect 15292 10610 15344 10616
rect 15200 10532 15252 10538
rect 15200 10474 15252 10480
rect 15304 10130 15332 10610
rect 15108 10124 15160 10130
rect 15108 10066 15160 10072
rect 15292 10124 15344 10130
rect 15292 10066 15344 10072
rect 15120 9654 15148 10066
rect 15292 9988 15344 9994
rect 15292 9930 15344 9936
rect 15108 9648 15160 9654
rect 15108 9590 15160 9596
rect 15304 9489 15332 9930
rect 15290 9480 15346 9489
rect 15200 9444 15252 9450
rect 15290 9415 15346 9424
rect 15200 9386 15252 9392
rect 15212 9178 15240 9386
rect 15200 9172 15252 9178
rect 15200 9114 15252 9120
rect 15396 9092 15424 12174
rect 15580 10146 15608 13126
rect 15672 12238 15700 14214
rect 15660 12232 15712 12238
rect 15660 12174 15712 12180
rect 15660 12096 15712 12102
rect 15660 12038 15712 12044
rect 15672 11694 15700 12038
rect 15660 11688 15712 11694
rect 15660 11630 15712 11636
rect 15660 11552 15712 11558
rect 15660 11494 15712 11500
rect 15672 10674 15700 11494
rect 15764 11014 15792 35974
rect 15948 31754 15976 57258
rect 17040 56908 17092 56914
rect 17040 56850 17092 56856
rect 16304 38548 16356 38554
rect 16304 38490 16356 38496
rect 16316 37466 16344 38490
rect 16304 37460 16356 37466
rect 16304 37402 16356 37408
rect 16488 37460 16540 37466
rect 16488 37402 16540 37408
rect 16500 36038 16528 37402
rect 16488 36032 16540 36038
rect 16488 35974 16540 35980
rect 16580 35692 16632 35698
rect 16580 35634 16632 35640
rect 16592 32774 16620 35634
rect 16948 33312 17000 33318
rect 16948 33254 17000 33260
rect 16580 32768 16632 32774
rect 16580 32710 16632 32716
rect 16488 32496 16540 32502
rect 16488 32438 16540 32444
rect 15948 31726 16252 31754
rect 15936 22024 15988 22030
rect 15936 21966 15988 21972
rect 15844 21684 15896 21690
rect 15844 21626 15896 21632
rect 15856 20942 15884 21626
rect 15948 21146 15976 21966
rect 16028 21548 16080 21554
rect 16028 21490 16080 21496
rect 16040 21146 16068 21490
rect 16120 21344 16172 21350
rect 16120 21286 16172 21292
rect 15936 21140 15988 21146
rect 15936 21082 15988 21088
rect 16028 21140 16080 21146
rect 16028 21082 16080 21088
rect 15844 20936 15896 20942
rect 16028 20936 16080 20942
rect 15844 20878 15896 20884
rect 15948 20884 16028 20890
rect 15948 20878 16080 20884
rect 15948 20862 16068 20878
rect 15844 20392 15896 20398
rect 15844 20334 15896 20340
rect 15856 17542 15884 20334
rect 15948 17610 15976 20862
rect 16028 19168 16080 19174
rect 16028 19110 16080 19116
rect 16040 18290 16068 19110
rect 16028 18284 16080 18290
rect 16028 18226 16080 18232
rect 16028 18080 16080 18086
rect 16028 18022 16080 18028
rect 15936 17604 15988 17610
rect 15936 17546 15988 17552
rect 15844 17536 15896 17542
rect 15844 17478 15896 17484
rect 16040 17354 16068 18022
rect 16132 17626 16160 21286
rect 16224 18086 16252 31726
rect 16396 21956 16448 21962
rect 16396 21898 16448 21904
rect 16304 21548 16356 21554
rect 16304 21490 16356 21496
rect 16316 21078 16344 21490
rect 16304 21072 16356 21078
rect 16304 21014 16356 21020
rect 16408 20942 16436 21898
rect 16396 20936 16448 20942
rect 16396 20878 16448 20884
rect 16396 18828 16448 18834
rect 16396 18770 16448 18776
rect 16408 18290 16436 18770
rect 16396 18284 16448 18290
rect 16396 18226 16448 18232
rect 16212 18080 16264 18086
rect 16212 18022 16264 18028
rect 16396 18080 16448 18086
rect 16396 18022 16448 18028
rect 16132 17610 16344 17626
rect 16132 17604 16356 17610
rect 16132 17598 16304 17604
rect 16304 17546 16356 17552
rect 16040 17326 16252 17354
rect 16120 17196 16172 17202
rect 16120 17138 16172 17144
rect 16132 16114 16160 17138
rect 16120 16108 16172 16114
rect 16120 16050 16172 16056
rect 15844 15088 15896 15094
rect 15844 15030 15896 15036
rect 15752 11008 15804 11014
rect 15752 10950 15804 10956
rect 15856 10742 15884 15030
rect 16028 15020 16080 15026
rect 16028 14962 16080 14968
rect 15936 14952 15988 14958
rect 15936 14894 15988 14900
rect 15948 14822 15976 14894
rect 15936 14816 15988 14822
rect 15936 14758 15988 14764
rect 16040 13530 16068 14962
rect 16028 13524 16080 13530
rect 16028 13466 16080 13472
rect 15936 13184 15988 13190
rect 15936 13126 15988 13132
rect 15948 12918 15976 13126
rect 15936 12912 15988 12918
rect 15936 12854 15988 12860
rect 16132 12442 16160 16050
rect 16120 12436 16172 12442
rect 16120 12378 16172 12384
rect 15936 12232 15988 12238
rect 15936 12174 15988 12180
rect 15948 11898 15976 12174
rect 16120 12164 16172 12170
rect 16120 12106 16172 12112
rect 15936 11892 15988 11898
rect 15936 11834 15988 11840
rect 16132 11801 16160 12106
rect 16118 11792 16174 11801
rect 16118 11727 16174 11736
rect 16224 10826 16252 17326
rect 16408 17134 16436 18022
rect 16396 17128 16448 17134
rect 16396 17070 16448 17076
rect 16396 16448 16448 16454
rect 16396 16390 16448 16396
rect 16304 16108 16356 16114
rect 16304 16050 16356 16056
rect 16316 15638 16344 16050
rect 16304 15632 16356 15638
rect 16304 15574 16356 15580
rect 16408 15094 16436 16390
rect 16396 15088 16448 15094
rect 16396 15030 16448 15036
rect 16304 13388 16356 13394
rect 16304 13330 16356 13336
rect 16040 10798 16252 10826
rect 15844 10736 15896 10742
rect 15844 10678 15896 10684
rect 15660 10668 15712 10674
rect 15660 10610 15712 10616
rect 15580 10118 15792 10146
rect 15660 10056 15712 10062
rect 15660 9998 15712 10004
rect 15568 9580 15620 9586
rect 15568 9522 15620 9528
rect 15580 9194 15608 9522
rect 15672 9382 15700 9998
rect 15660 9376 15712 9382
rect 15660 9318 15712 9324
rect 15580 9166 15700 9194
rect 15396 9064 15608 9092
rect 14924 8900 14976 8906
rect 14924 8842 14976 8848
rect 14936 8634 14964 8842
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 14924 8628 14976 8634
rect 14924 8570 14976 8576
rect 15120 8566 15148 8774
rect 15108 8560 15160 8566
rect 15108 8502 15160 8508
rect 15292 8492 15344 8498
rect 15476 8492 15528 8498
rect 15344 8452 15476 8480
rect 15292 8434 15344 8440
rect 15476 8434 15528 8440
rect 15106 8256 15162 8265
rect 15106 8191 15162 8200
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 15028 7546 15056 7822
rect 15016 7540 15068 7546
rect 15016 7482 15068 7488
rect 14830 6080 14886 6089
rect 14830 6015 14886 6024
rect 14740 5296 14792 5302
rect 14740 5238 14792 5244
rect 14752 4758 14780 5238
rect 14740 4752 14792 4758
rect 14740 4694 14792 4700
rect 14740 4616 14792 4622
rect 14740 4558 14792 4564
rect 14648 3732 14700 3738
rect 14648 3674 14700 3680
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 14464 3052 14516 3058
rect 14464 2994 14516 3000
rect 14384 1578 14412 2994
rect 14384 1550 14504 1578
rect 14476 800 14504 1550
rect 14752 800 14780 4558
rect 14844 4078 14872 6015
rect 14832 4072 14884 4078
rect 14832 4014 14884 4020
rect 15120 3534 15148 8191
rect 15290 8120 15346 8129
rect 15290 8055 15346 8064
rect 15200 8016 15252 8022
rect 15200 7958 15252 7964
rect 15212 7886 15240 7958
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 15304 7750 15332 8055
rect 15488 7886 15516 8434
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15292 7744 15344 7750
rect 15292 7686 15344 7692
rect 15488 7478 15516 7822
rect 15476 7472 15528 7478
rect 15476 7414 15528 7420
rect 15198 7304 15254 7313
rect 15198 7239 15200 7248
rect 15252 7239 15254 7248
rect 15200 7210 15252 7216
rect 15384 6384 15436 6390
rect 15382 6352 15384 6361
rect 15436 6352 15438 6361
rect 15200 6316 15252 6322
rect 15488 6322 15516 7414
rect 15382 6287 15438 6296
rect 15476 6316 15528 6322
rect 15200 6258 15252 6264
rect 15476 6258 15528 6264
rect 15212 4758 15240 6258
rect 15488 5710 15516 6258
rect 15476 5704 15528 5710
rect 15476 5646 15528 5652
rect 15580 5642 15608 9064
rect 15672 8294 15700 9166
rect 15660 8288 15712 8294
rect 15764 8265 15792 10118
rect 15934 9616 15990 9625
rect 16040 9602 16068 10798
rect 16212 10736 16264 10742
rect 15990 9574 16068 9602
rect 16132 10696 16212 10724
rect 15934 9551 15936 9560
rect 15988 9551 15990 9560
rect 15936 9522 15988 9528
rect 15842 9480 15898 9489
rect 15842 9415 15898 9424
rect 15660 8230 15712 8236
rect 15750 8256 15806 8265
rect 15750 8191 15806 8200
rect 15752 7812 15804 7818
rect 15752 7754 15804 7760
rect 15660 7472 15712 7478
rect 15660 7414 15712 7420
rect 15672 6390 15700 7414
rect 15764 7410 15792 7754
rect 15752 7404 15804 7410
rect 15752 7346 15804 7352
rect 15660 6384 15712 6390
rect 15660 6326 15712 6332
rect 15672 5778 15700 6326
rect 15764 6322 15792 7346
rect 15752 6316 15804 6322
rect 15752 6258 15804 6264
rect 15856 5778 15884 9415
rect 16028 7880 16080 7886
rect 16028 7822 16080 7828
rect 16040 7750 16068 7822
rect 16028 7744 16080 7750
rect 16028 7686 16080 7692
rect 16040 7410 16068 7686
rect 16028 7404 16080 7410
rect 16028 7346 16080 7352
rect 16132 6361 16160 10696
rect 16212 10678 16264 10684
rect 16212 10600 16264 10606
rect 16212 10542 16264 10548
rect 16224 10198 16252 10542
rect 16212 10192 16264 10198
rect 16212 10134 16264 10140
rect 16224 9586 16252 10134
rect 16212 9580 16264 9586
rect 16212 9522 16264 9528
rect 16316 9450 16344 13330
rect 16396 12436 16448 12442
rect 16396 12378 16448 12384
rect 16408 11558 16436 12378
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 16396 11144 16448 11150
rect 16396 11086 16448 11092
rect 16408 9722 16436 11086
rect 16500 10742 16528 32438
rect 16672 22568 16724 22574
rect 16672 22510 16724 22516
rect 16580 21480 16632 21486
rect 16580 21422 16632 21428
rect 16592 20890 16620 21422
rect 16684 21010 16712 22510
rect 16764 22432 16816 22438
rect 16764 22374 16816 22380
rect 16672 21004 16724 21010
rect 16672 20946 16724 20952
rect 16776 20942 16804 22374
rect 16856 21480 16908 21486
rect 16856 21422 16908 21428
rect 16764 20936 16816 20942
rect 16592 20862 16712 20890
rect 16764 20878 16816 20884
rect 16684 20466 16712 20862
rect 16672 20460 16724 20466
rect 16672 20402 16724 20408
rect 16580 20256 16632 20262
rect 16580 20198 16632 20204
rect 16592 18766 16620 20198
rect 16580 18760 16632 18766
rect 16580 18702 16632 18708
rect 16684 17882 16712 20402
rect 16868 19854 16896 21422
rect 16856 19848 16908 19854
rect 16856 19790 16908 19796
rect 16868 19378 16896 19790
rect 16856 19372 16908 19378
rect 16856 19314 16908 19320
rect 16868 18290 16896 19314
rect 16856 18284 16908 18290
rect 16856 18226 16908 18232
rect 16672 17876 16724 17882
rect 16672 17818 16724 17824
rect 16580 17332 16632 17338
rect 16580 17274 16632 17280
rect 16672 17332 16724 17338
rect 16672 17274 16724 17280
rect 16592 16590 16620 17274
rect 16580 16584 16632 16590
rect 16580 16526 16632 16532
rect 16580 16448 16632 16454
rect 16580 16390 16632 16396
rect 16592 11370 16620 16390
rect 16684 16250 16712 17274
rect 16764 17128 16816 17134
rect 16764 17070 16816 17076
rect 16776 16726 16804 17070
rect 16764 16720 16816 16726
rect 16764 16662 16816 16668
rect 16868 16522 16896 18226
rect 16856 16516 16908 16522
rect 16856 16458 16908 16464
rect 16672 16244 16724 16250
rect 16672 16186 16724 16192
rect 16868 15978 16896 16458
rect 16960 16454 16988 33254
rect 16948 16448 17000 16454
rect 16948 16390 17000 16396
rect 16856 15972 16908 15978
rect 16856 15914 16908 15920
rect 16672 15496 16724 15502
rect 16672 15438 16724 15444
rect 16684 15026 16712 15438
rect 16868 15026 16896 15914
rect 16672 15020 16724 15026
rect 16672 14962 16724 14968
rect 16856 15020 16908 15026
rect 16856 14962 16908 14968
rect 16764 14952 16816 14958
rect 16764 14894 16816 14900
rect 16776 14346 16804 14894
rect 16764 14340 16816 14346
rect 16764 14282 16816 14288
rect 16868 13938 16896 14962
rect 16856 13932 16908 13938
rect 16856 13874 16908 13880
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 16672 12708 16724 12714
rect 16672 12650 16724 12656
rect 16684 12442 16712 12650
rect 16672 12436 16724 12442
rect 16672 12378 16724 12384
rect 16672 11756 16724 11762
rect 16672 11698 16724 11704
rect 16684 11665 16712 11698
rect 16670 11656 16726 11665
rect 16670 11591 16726 11600
rect 16592 11342 16712 11370
rect 16776 11354 16804 13262
rect 16868 11762 16896 13874
rect 17052 11801 17080 56850
rect 17328 34134 17356 60998
rect 17420 45490 17448 61066
rect 17868 60512 17920 60518
rect 17868 60454 17920 60460
rect 17880 60178 17908 60454
rect 17868 60172 17920 60178
rect 17868 60114 17920 60120
rect 17592 60036 17644 60042
rect 17592 59978 17644 59984
rect 17500 59968 17552 59974
rect 17500 59910 17552 59916
rect 17512 50289 17540 59910
rect 17604 59566 17632 59978
rect 18248 59702 18276 61270
rect 18708 61198 18736 63294
rect 19246 63200 19302 64000
rect 19982 63322 20038 64000
rect 19812 63294 20038 63322
rect 18696 61192 18748 61198
rect 18696 61134 18748 61140
rect 18880 61124 18932 61130
rect 18880 61066 18932 61072
rect 18420 60580 18472 60586
rect 18420 60522 18472 60528
rect 18432 60110 18460 60522
rect 18420 60104 18472 60110
rect 18420 60046 18472 60052
rect 18604 60104 18656 60110
rect 18604 60046 18656 60052
rect 18236 59696 18288 59702
rect 18236 59638 18288 59644
rect 17960 59628 18012 59634
rect 17960 59570 18012 59576
rect 17592 59560 17644 59566
rect 17592 59502 17644 59508
rect 17972 58886 18000 59570
rect 18616 59401 18644 60046
rect 18602 59392 18658 59401
rect 18602 59327 18658 59336
rect 17960 58880 18012 58886
rect 17960 58822 18012 58828
rect 17868 51536 17920 51542
rect 17868 51478 17920 51484
rect 17498 50280 17554 50289
rect 17498 50215 17554 50224
rect 17880 48278 17908 51478
rect 18604 49088 18656 49094
rect 18604 49030 18656 49036
rect 17868 48272 17920 48278
rect 17868 48214 17920 48220
rect 17408 45484 17460 45490
rect 17408 45426 17460 45432
rect 17684 45280 17736 45286
rect 17684 45222 17736 45228
rect 17316 34128 17368 34134
rect 17316 34070 17368 34076
rect 17132 33856 17184 33862
rect 17132 33798 17184 33804
rect 17144 33658 17172 33798
rect 17132 33652 17184 33658
rect 17132 33594 17184 33600
rect 17696 30666 17724 45222
rect 18616 40458 18644 49030
rect 18604 40452 18656 40458
rect 18604 40394 18656 40400
rect 18788 37188 18840 37194
rect 18788 37130 18840 37136
rect 18800 36786 18828 37130
rect 18892 36854 18920 61066
rect 19260 60874 19288 63200
rect 19432 61668 19484 61674
rect 19432 61610 19484 61616
rect 19260 60846 19380 60874
rect 19352 60790 19380 60846
rect 19340 60784 19392 60790
rect 19340 60726 19392 60732
rect 19248 60036 19300 60042
rect 19248 59978 19300 59984
rect 19260 59566 19288 59978
rect 19444 59650 19472 61610
rect 19812 61198 19840 63294
rect 19982 63200 20038 63294
rect 20718 63200 20774 64000
rect 21454 63322 21510 64000
rect 21284 63294 21510 63322
rect 20732 61198 20760 63200
rect 21180 61600 21232 61606
rect 21180 61542 21232 61548
rect 19800 61192 19852 61198
rect 19800 61134 19852 61140
rect 20720 61192 20772 61198
rect 20720 61134 20772 61140
rect 20444 61124 20496 61130
rect 20444 61066 20496 61072
rect 21088 61124 21140 61130
rect 21088 61066 21140 61072
rect 19574 60956 19882 60965
rect 19574 60954 19580 60956
rect 19636 60954 19660 60956
rect 19716 60954 19740 60956
rect 19796 60954 19820 60956
rect 19876 60954 19882 60956
rect 19636 60902 19638 60954
rect 19818 60902 19820 60954
rect 19574 60900 19580 60902
rect 19636 60900 19660 60902
rect 19716 60900 19740 60902
rect 19796 60900 19820 60902
rect 19876 60900 19882 60902
rect 19574 60891 19882 60900
rect 20260 60308 20312 60314
rect 20260 60250 20312 60256
rect 19984 60104 20036 60110
rect 19984 60046 20036 60052
rect 19574 59868 19882 59877
rect 19574 59866 19580 59868
rect 19636 59866 19660 59868
rect 19716 59866 19740 59868
rect 19796 59866 19820 59868
rect 19876 59866 19882 59868
rect 19636 59814 19638 59866
rect 19818 59814 19820 59866
rect 19574 59812 19580 59814
rect 19636 59812 19660 59814
rect 19716 59812 19740 59814
rect 19796 59812 19820 59814
rect 19876 59812 19882 59814
rect 19574 59803 19882 59812
rect 19444 59622 19748 59650
rect 19996 59634 20024 60046
rect 19248 59560 19300 59566
rect 19248 59502 19300 59508
rect 19524 59152 19576 59158
rect 19524 59094 19576 59100
rect 19536 58970 19564 59094
rect 19720 59022 19748 59622
rect 19984 59628 20036 59634
rect 19984 59570 20036 59576
rect 20168 59424 20220 59430
rect 20168 59366 20220 59372
rect 19352 58942 19564 58970
rect 19708 59016 19760 59022
rect 19708 58958 19760 58964
rect 19156 38480 19208 38486
rect 19156 38422 19208 38428
rect 18880 36848 18932 36854
rect 18880 36790 18932 36796
rect 18420 36780 18472 36786
rect 18420 36722 18472 36728
rect 18788 36780 18840 36786
rect 18788 36722 18840 36728
rect 17684 30660 17736 30666
rect 17684 30602 17736 30608
rect 17960 30592 18012 30598
rect 17960 30534 18012 30540
rect 17972 30394 18000 30534
rect 17960 30388 18012 30394
rect 17960 30330 18012 30336
rect 17224 25900 17276 25906
rect 17224 25842 17276 25848
rect 17236 25498 17264 25842
rect 18432 25838 18460 36722
rect 18880 30252 18932 30258
rect 18880 30194 18932 30200
rect 18972 30252 19024 30258
rect 18972 30194 19024 30200
rect 18892 27062 18920 30194
rect 18984 29578 19012 30194
rect 18972 29572 19024 29578
rect 18972 29514 19024 29520
rect 18880 27056 18932 27062
rect 18880 26998 18932 27004
rect 18420 25832 18472 25838
rect 18420 25774 18472 25780
rect 17224 25492 17276 25498
rect 17224 25434 17276 25440
rect 18788 23248 18840 23254
rect 18788 23190 18840 23196
rect 17868 23112 17920 23118
rect 17868 23054 17920 23060
rect 17880 22710 17908 23054
rect 18236 23044 18288 23050
rect 18236 22986 18288 22992
rect 17960 22976 18012 22982
rect 17960 22918 18012 22924
rect 17868 22704 17920 22710
rect 17868 22646 17920 22652
rect 17972 22642 18000 22918
rect 18248 22778 18276 22986
rect 18236 22772 18288 22778
rect 18236 22714 18288 22720
rect 17960 22636 18012 22642
rect 17960 22578 18012 22584
rect 18144 22636 18196 22642
rect 18144 22578 18196 22584
rect 18328 22636 18380 22642
rect 18328 22578 18380 22584
rect 17132 22024 17184 22030
rect 17132 21966 17184 21972
rect 17144 16726 17172 21966
rect 18156 21962 18184 22578
rect 18144 21956 18196 21962
rect 18144 21898 18196 21904
rect 18052 21548 18104 21554
rect 18052 21490 18104 21496
rect 17316 21344 17368 21350
rect 17316 21286 17368 21292
rect 17224 20936 17276 20942
rect 17224 20878 17276 20884
rect 17236 20398 17264 20878
rect 17224 20392 17276 20398
rect 17224 20334 17276 20340
rect 17328 17882 17356 21286
rect 17960 21004 18012 21010
rect 17960 20946 18012 20952
rect 17868 20460 17920 20466
rect 17868 20402 17920 20408
rect 17592 20324 17644 20330
rect 17592 20266 17644 20272
rect 17604 18902 17632 20266
rect 17776 19372 17828 19378
rect 17776 19314 17828 19320
rect 17592 18896 17644 18902
rect 17592 18838 17644 18844
rect 17316 17876 17368 17882
rect 17316 17818 17368 17824
rect 17788 17542 17816 19314
rect 17880 19174 17908 20402
rect 17972 19310 18000 20946
rect 17960 19304 18012 19310
rect 17960 19246 18012 19252
rect 17868 19168 17920 19174
rect 17868 19110 17920 19116
rect 17880 18358 17908 19110
rect 18064 18834 18092 21490
rect 18156 20806 18184 21898
rect 18340 21690 18368 22578
rect 18328 21684 18380 21690
rect 18328 21626 18380 21632
rect 18800 21554 18828 23190
rect 19168 22094 19196 38422
rect 19352 37874 19380 58942
rect 19984 58880 20036 58886
rect 19984 58822 20036 58828
rect 19574 58780 19882 58789
rect 19574 58778 19580 58780
rect 19636 58778 19660 58780
rect 19716 58778 19740 58780
rect 19796 58778 19820 58780
rect 19876 58778 19882 58780
rect 19636 58726 19638 58778
rect 19818 58726 19820 58778
rect 19574 58724 19580 58726
rect 19636 58724 19660 58726
rect 19716 58724 19740 58726
rect 19796 58724 19820 58726
rect 19876 58724 19882 58726
rect 19574 58715 19882 58724
rect 19574 57692 19882 57701
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57627 19882 57636
rect 19574 56604 19882 56613
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56539 19882 56548
rect 19574 55516 19882 55525
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55451 19882 55460
rect 19574 54428 19882 54437
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54363 19882 54372
rect 19574 53340 19882 53349
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53275 19882 53284
rect 19574 52252 19882 52261
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52187 19882 52196
rect 19574 51164 19882 51173
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51099 19882 51108
rect 19574 50076 19882 50085
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50011 19882 50020
rect 19574 48988 19882 48997
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48923 19882 48932
rect 19574 47900 19882 47909
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47835 19882 47844
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 19996 41414 20024 58822
rect 19996 41386 20116 41414
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 19432 38412 19484 38418
rect 19432 38354 19484 38360
rect 19984 38412 20036 38418
rect 19984 38354 20036 38360
rect 19444 37890 19472 38354
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 19444 37874 19748 37890
rect 19340 37868 19392 37874
rect 19444 37868 19760 37874
rect 19444 37862 19708 37868
rect 19340 37810 19392 37816
rect 19708 37810 19760 37816
rect 19340 37256 19392 37262
rect 19340 37198 19392 37204
rect 19248 37120 19300 37126
rect 19248 37062 19300 37068
rect 19260 35766 19288 37062
rect 19352 36650 19380 37198
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19432 36780 19484 36786
rect 19432 36722 19484 36728
rect 19340 36644 19392 36650
rect 19340 36586 19392 36592
rect 19352 35834 19380 36586
rect 19340 35828 19392 35834
rect 19340 35770 19392 35776
rect 19248 35760 19300 35766
rect 19248 35702 19300 35708
rect 19260 31482 19288 35702
rect 19340 35556 19392 35562
rect 19340 35498 19392 35504
rect 19352 34746 19380 35498
rect 19340 34740 19392 34746
rect 19340 34682 19392 34688
rect 19444 34610 19472 36722
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19996 34678 20024 38354
rect 20088 36854 20116 41386
rect 20180 38350 20208 59366
rect 20272 51338 20300 60250
rect 20456 60110 20484 61066
rect 20904 61056 20956 61062
rect 20904 60998 20956 61004
rect 20628 60580 20680 60586
rect 20628 60522 20680 60528
rect 20536 60512 20588 60518
rect 20536 60454 20588 60460
rect 20548 60110 20576 60454
rect 20444 60104 20496 60110
rect 20444 60046 20496 60052
rect 20536 60104 20588 60110
rect 20536 60046 20588 60052
rect 20260 51332 20312 51338
rect 20260 51274 20312 51280
rect 20444 51264 20496 51270
rect 20444 51206 20496 51212
rect 20456 41414 20484 51206
rect 20456 41386 20576 41414
rect 20548 38350 20576 41386
rect 20640 38418 20668 60522
rect 20720 60308 20772 60314
rect 20720 60250 20772 60256
rect 20732 60110 20760 60250
rect 20720 60104 20772 60110
rect 20720 60046 20772 60052
rect 20720 52420 20772 52426
rect 20720 52362 20772 52368
rect 20732 52018 20760 52362
rect 20720 52012 20772 52018
rect 20720 51954 20772 51960
rect 20732 45558 20760 51954
rect 20720 45552 20772 45558
rect 20720 45494 20772 45500
rect 20732 41414 20760 45494
rect 20732 41386 20852 41414
rect 20628 38412 20680 38418
rect 20628 38354 20680 38360
rect 20168 38344 20220 38350
rect 20168 38286 20220 38292
rect 20536 38344 20588 38350
rect 20536 38286 20588 38292
rect 20168 38208 20220 38214
rect 20168 38150 20220 38156
rect 20076 36848 20128 36854
rect 20076 36790 20128 36796
rect 20180 36718 20208 38150
rect 20824 38026 20852 41386
rect 20916 40186 20944 60998
rect 21100 59634 21128 61066
rect 21088 59628 21140 59634
rect 21088 59570 21140 59576
rect 21192 59430 21220 61542
rect 21284 61198 21312 63294
rect 21454 63200 21510 63294
rect 22190 63322 22246 64000
rect 22926 63322 22982 64000
rect 23662 63322 23718 64000
rect 22190 63294 22416 63322
rect 22190 63200 22246 63294
rect 22100 61328 22152 61334
rect 22100 61270 22152 61276
rect 21272 61192 21324 61198
rect 21272 61134 21324 61140
rect 22112 60722 22140 61270
rect 22388 61198 22416 63294
rect 22926 63294 23244 63322
rect 22926 63200 22982 63294
rect 22836 61260 22888 61266
rect 22836 61202 22888 61208
rect 22376 61192 22428 61198
rect 22376 61134 22428 61140
rect 22744 61124 22796 61130
rect 22744 61066 22796 61072
rect 22756 60761 22784 61066
rect 22742 60752 22798 60761
rect 22100 60716 22152 60722
rect 22100 60658 22152 60664
rect 22560 60716 22612 60722
rect 22742 60687 22798 60696
rect 22560 60658 22612 60664
rect 22468 60512 22520 60518
rect 22468 60454 22520 60460
rect 22098 60344 22154 60353
rect 21836 60302 22098 60330
rect 21364 60240 21416 60246
rect 21364 60182 21416 60188
rect 21272 60036 21324 60042
rect 21272 59978 21324 59984
rect 21180 59424 21232 59430
rect 21180 59366 21232 59372
rect 21284 55214 21312 59978
rect 21192 55186 21312 55214
rect 21192 51406 21220 55186
rect 21180 51400 21232 51406
rect 21180 51342 21232 51348
rect 21192 45554 21220 51342
rect 21100 45526 21220 45554
rect 20904 40180 20956 40186
rect 20904 40122 20956 40128
rect 20996 40044 21048 40050
rect 20996 39986 21048 39992
rect 20824 37998 20944 38026
rect 20718 37904 20774 37913
rect 20260 37868 20312 37874
rect 20916 37874 20944 37998
rect 20718 37839 20774 37848
rect 20812 37868 20864 37874
rect 20260 37810 20312 37816
rect 20272 37398 20300 37810
rect 20444 37732 20496 37738
rect 20444 37674 20496 37680
rect 20352 37664 20404 37670
rect 20352 37606 20404 37612
rect 20260 37392 20312 37398
rect 20260 37334 20312 37340
rect 20260 36848 20312 36854
rect 20260 36790 20312 36796
rect 20168 36712 20220 36718
rect 20168 36654 20220 36660
rect 20076 36576 20128 36582
rect 20076 36518 20128 36524
rect 20088 35494 20116 36518
rect 20168 36168 20220 36174
rect 20168 36110 20220 36116
rect 20180 35834 20208 36110
rect 20168 35828 20220 35834
rect 20168 35770 20220 35776
rect 20076 35488 20128 35494
rect 20076 35430 20128 35436
rect 19984 34672 20036 34678
rect 19984 34614 20036 34620
rect 19432 34604 19484 34610
rect 19432 34546 19484 34552
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 20272 31958 20300 36790
rect 20260 31952 20312 31958
rect 20260 31894 20312 31900
rect 20364 31754 20392 37606
rect 20456 36174 20484 37674
rect 20628 37664 20680 37670
rect 20628 37606 20680 37612
rect 20536 37256 20588 37262
rect 20536 37198 20588 37204
rect 20548 36854 20576 37198
rect 20536 36848 20588 36854
rect 20536 36790 20588 36796
rect 20640 36310 20668 37606
rect 20732 37466 20760 37839
rect 20812 37810 20864 37816
rect 20904 37868 20956 37874
rect 20904 37810 20956 37816
rect 20824 37466 20852 37810
rect 20720 37460 20772 37466
rect 20720 37402 20772 37408
rect 20812 37460 20864 37466
rect 20812 37402 20864 37408
rect 21008 37194 21036 39986
rect 21100 38282 21128 45526
rect 21180 40928 21232 40934
rect 21180 40870 21232 40876
rect 21192 40118 21220 40870
rect 21180 40112 21232 40118
rect 21180 40054 21232 40060
rect 21088 38276 21140 38282
rect 21088 38218 21140 38224
rect 21088 37868 21140 37874
rect 21088 37810 21140 37816
rect 21100 37330 21128 37810
rect 21272 37732 21324 37738
rect 21272 37674 21324 37680
rect 21088 37324 21140 37330
rect 21088 37266 21140 37272
rect 20996 37188 21048 37194
rect 20996 37130 21048 37136
rect 20996 36780 21048 36786
rect 20996 36722 21048 36728
rect 21008 36310 21036 36722
rect 20628 36304 20680 36310
rect 20628 36246 20680 36252
rect 20996 36304 21048 36310
rect 20996 36246 21048 36252
rect 20720 36236 20772 36242
rect 20720 36178 20772 36184
rect 20444 36168 20496 36174
rect 20444 36110 20496 36116
rect 20364 31726 20484 31754
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19248 31476 19300 31482
rect 19248 31418 19300 31424
rect 19260 30258 19288 31418
rect 19340 30796 19392 30802
rect 19340 30738 19392 30744
rect 19352 30394 19380 30738
rect 20352 30660 20404 30666
rect 20352 30602 20404 30608
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19340 30388 19392 30394
rect 19340 30330 19392 30336
rect 19248 30252 19300 30258
rect 19248 30194 19300 30200
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19340 22500 19392 22506
rect 19340 22442 19392 22448
rect 19076 22066 19196 22094
rect 18788 21548 18840 21554
rect 18788 21490 18840 21496
rect 18144 20800 18196 20806
rect 18144 20742 18196 20748
rect 18880 20596 18932 20602
rect 18880 20538 18932 20544
rect 18510 20496 18566 20505
rect 18510 20431 18512 20440
rect 18564 20431 18566 20440
rect 18512 20402 18564 20408
rect 18052 18828 18104 18834
rect 18052 18770 18104 18776
rect 17868 18352 17920 18358
rect 17868 18294 17920 18300
rect 17776 17536 17828 17542
rect 17776 17478 17828 17484
rect 18892 16998 18920 20538
rect 18144 16992 18196 16998
rect 18144 16934 18196 16940
rect 18880 16992 18932 16998
rect 18880 16934 18932 16940
rect 17132 16720 17184 16726
rect 17132 16662 17184 16668
rect 17408 16720 17460 16726
rect 17408 16662 17460 16668
rect 17224 15360 17276 15366
rect 17224 15302 17276 15308
rect 17236 13394 17264 15302
rect 17316 13524 17368 13530
rect 17316 13466 17368 13472
rect 17224 13388 17276 13394
rect 17224 13330 17276 13336
rect 17236 12986 17264 13330
rect 17224 12980 17276 12986
rect 17224 12922 17276 12928
rect 17328 12850 17356 13466
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 17420 12782 17448 16662
rect 17960 16448 18012 16454
rect 17960 16390 18012 16396
rect 18052 16448 18104 16454
rect 18052 16390 18104 16396
rect 17684 16108 17736 16114
rect 17684 16050 17736 16056
rect 17592 14340 17644 14346
rect 17592 14282 17644 14288
rect 17408 12776 17460 12782
rect 17408 12718 17460 12724
rect 17420 11898 17448 12718
rect 17408 11892 17460 11898
rect 17408 11834 17460 11840
rect 17038 11792 17094 11801
rect 16856 11756 16908 11762
rect 17038 11727 17094 11736
rect 17408 11756 17460 11762
rect 16856 11698 16908 11704
rect 16684 11234 16712 11342
rect 16764 11348 16816 11354
rect 16764 11290 16816 11296
rect 16684 11206 16804 11234
rect 16580 11144 16632 11150
rect 16580 11086 16632 11092
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 16488 10736 16540 10742
rect 16488 10678 16540 10684
rect 16488 10600 16540 10606
rect 16488 10542 16540 10548
rect 16500 10062 16528 10542
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 16396 9716 16448 9722
rect 16396 9658 16448 9664
rect 16500 9450 16528 9998
rect 16304 9444 16356 9450
rect 16304 9386 16356 9392
rect 16488 9444 16540 9450
rect 16488 9386 16540 9392
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16224 6662 16252 9114
rect 16500 8022 16528 9386
rect 16592 8634 16620 11086
rect 16684 10062 16712 11086
rect 16672 10056 16724 10062
rect 16672 9998 16724 10004
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 16684 8498 16712 9998
rect 16672 8492 16724 8498
rect 16672 8434 16724 8440
rect 16684 8022 16712 8434
rect 16488 8016 16540 8022
rect 16488 7958 16540 7964
rect 16672 8016 16724 8022
rect 16672 7958 16724 7964
rect 16304 7948 16356 7954
rect 16304 7890 16356 7896
rect 16316 7857 16344 7890
rect 16302 7848 16358 7857
rect 16302 7783 16358 7792
rect 16776 7750 16804 11206
rect 16854 11112 16910 11121
rect 16854 11047 16910 11056
rect 16764 7744 16816 7750
rect 16764 7686 16816 7692
rect 16776 7546 16804 7686
rect 16764 7540 16816 7546
rect 16764 7482 16816 7488
rect 16304 7472 16356 7478
rect 16304 7414 16356 7420
rect 16316 7342 16344 7414
rect 16304 7336 16356 7342
rect 16304 7278 16356 7284
rect 16212 6656 16264 6662
rect 16212 6598 16264 6604
rect 16118 6352 16174 6361
rect 16118 6287 16174 6296
rect 16212 6316 16264 6322
rect 16316 6304 16344 7278
rect 16868 7154 16896 11047
rect 17052 10742 17080 11727
rect 17408 11698 17460 11704
rect 17420 11529 17448 11698
rect 17406 11520 17462 11529
rect 17406 11455 17462 11464
rect 17604 11150 17632 14282
rect 17592 11144 17644 11150
rect 17592 11086 17644 11092
rect 17132 11076 17184 11082
rect 17132 11018 17184 11024
rect 17040 10736 17092 10742
rect 17040 10678 17092 10684
rect 17144 10606 17172 11018
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 17132 10600 17184 10606
rect 17132 10542 17184 10548
rect 17040 8968 17092 8974
rect 17040 8910 17092 8916
rect 17052 8673 17080 8910
rect 17038 8664 17094 8673
rect 17038 8599 17094 8608
rect 17052 8566 17080 8599
rect 17040 8560 17092 8566
rect 17040 8502 17092 8508
rect 17144 8498 17172 10542
rect 17224 8628 17276 8634
rect 17224 8570 17276 8576
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 17144 7410 17172 8434
rect 17236 7886 17264 8570
rect 17328 8430 17356 10610
rect 17696 10305 17724 16050
rect 17868 15904 17920 15910
rect 17868 15846 17920 15852
rect 17776 14272 17828 14278
rect 17776 14214 17828 14220
rect 17788 14006 17816 14214
rect 17776 14000 17828 14006
rect 17776 13942 17828 13948
rect 17880 13530 17908 15846
rect 17972 15094 18000 16390
rect 18064 15570 18092 16390
rect 18052 15564 18104 15570
rect 18052 15506 18104 15512
rect 18156 15162 18184 16934
rect 18420 15360 18472 15366
rect 18420 15302 18472 15308
rect 18144 15156 18196 15162
rect 18144 15098 18196 15104
rect 17960 15088 18012 15094
rect 17960 15030 18012 15036
rect 18328 15088 18380 15094
rect 18328 15030 18380 15036
rect 18052 14408 18104 14414
rect 18052 14350 18104 14356
rect 17960 13728 18012 13734
rect 17960 13670 18012 13676
rect 17868 13524 17920 13530
rect 17868 13466 17920 13472
rect 17868 13388 17920 13394
rect 17868 13330 17920 13336
rect 17776 12980 17828 12986
rect 17776 12922 17828 12928
rect 17788 11830 17816 12922
rect 17880 12918 17908 13330
rect 17972 13025 18000 13670
rect 17958 13016 18014 13025
rect 17958 12951 18014 12960
rect 17868 12912 17920 12918
rect 17868 12854 17920 12860
rect 17868 12096 17920 12102
rect 17868 12038 17920 12044
rect 17776 11824 17828 11830
rect 17776 11766 17828 11772
rect 17880 11257 17908 12038
rect 18064 11354 18092 14350
rect 18236 13864 18288 13870
rect 18236 13806 18288 13812
rect 18144 13388 18196 13394
rect 18144 13330 18196 13336
rect 18156 12986 18184 13330
rect 18144 12980 18196 12986
rect 18144 12922 18196 12928
rect 18144 12232 18196 12238
rect 18144 12174 18196 12180
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 17866 11248 17922 11257
rect 17866 11183 17868 11192
rect 17920 11183 17922 11192
rect 17960 11212 18012 11218
rect 17868 11154 17920 11160
rect 17960 11154 18012 11160
rect 17972 11098 18000 11154
rect 17880 11070 18000 11098
rect 17774 10432 17830 10441
rect 17774 10367 17830 10376
rect 17682 10296 17738 10305
rect 17682 10231 17738 10240
rect 17684 10192 17736 10198
rect 17684 10134 17736 10140
rect 17408 10056 17460 10062
rect 17408 9998 17460 10004
rect 17420 9722 17448 9998
rect 17408 9716 17460 9722
rect 17408 9658 17460 9664
rect 17316 8424 17368 8430
rect 17316 8366 17368 8372
rect 17328 7954 17356 8366
rect 17420 8294 17448 9658
rect 17592 9580 17644 9586
rect 17592 9522 17644 9528
rect 17500 9512 17552 9518
rect 17500 9454 17552 9460
rect 17512 8906 17540 9454
rect 17604 9042 17632 9522
rect 17592 9036 17644 9042
rect 17592 8978 17644 8984
rect 17500 8900 17552 8906
rect 17500 8842 17552 8848
rect 17512 8537 17540 8842
rect 17498 8528 17554 8537
rect 17498 8463 17554 8472
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17500 8016 17552 8022
rect 17500 7958 17552 7964
rect 17592 8016 17644 8022
rect 17592 7958 17644 7964
rect 17316 7948 17368 7954
rect 17316 7890 17368 7896
rect 17224 7880 17276 7886
rect 17224 7822 17276 7828
rect 17236 7478 17264 7822
rect 17224 7472 17276 7478
rect 17224 7414 17276 7420
rect 17132 7404 17184 7410
rect 17132 7346 17184 7352
rect 17040 7336 17092 7342
rect 17040 7278 17092 7284
rect 17052 7154 17080 7278
rect 17328 7274 17356 7890
rect 17408 7880 17460 7886
rect 17408 7822 17460 7828
rect 17316 7268 17368 7274
rect 17316 7210 17368 7216
rect 16868 7126 17080 7154
rect 17222 7032 17278 7041
rect 17222 6967 17278 6976
rect 16264 6276 16344 6304
rect 17040 6316 17092 6322
rect 16212 6258 16264 6264
rect 17040 6258 17092 6264
rect 16224 5846 16252 6258
rect 16396 6248 16448 6254
rect 16396 6190 16448 6196
rect 16212 5840 16264 5846
rect 16212 5782 16264 5788
rect 15660 5772 15712 5778
rect 15660 5714 15712 5720
rect 15844 5772 15896 5778
rect 15844 5714 15896 5720
rect 16408 5710 16436 6190
rect 16856 5840 16908 5846
rect 16856 5782 16908 5788
rect 16396 5704 16448 5710
rect 16396 5646 16448 5652
rect 16868 5642 16896 5782
rect 17052 5710 17080 6258
rect 17040 5704 17092 5710
rect 17092 5664 17172 5692
rect 17040 5646 17092 5652
rect 15568 5636 15620 5642
rect 15568 5578 15620 5584
rect 16856 5636 16908 5642
rect 16856 5578 16908 5584
rect 17144 5166 17172 5664
rect 17132 5160 17184 5166
rect 17132 5102 17184 5108
rect 16672 5024 16724 5030
rect 16672 4966 16724 4972
rect 15200 4752 15252 4758
rect 15200 4694 15252 4700
rect 15660 4752 15712 4758
rect 15660 4694 15712 4700
rect 15672 3534 15700 4694
rect 16396 4616 16448 4622
rect 16396 4558 16448 4564
rect 16580 4616 16632 4622
rect 16580 4558 16632 4564
rect 16120 4072 16172 4078
rect 16120 4014 16172 4020
rect 15936 3664 15988 3670
rect 15936 3606 15988 3612
rect 15108 3528 15160 3534
rect 15108 3470 15160 3476
rect 15660 3528 15712 3534
rect 15660 3470 15712 3476
rect 15568 3460 15620 3466
rect 15568 3402 15620 3408
rect 15292 3052 15344 3058
rect 15292 2994 15344 3000
rect 15016 2304 15068 2310
rect 15016 2246 15068 2252
rect 15028 800 15056 2246
rect 15304 800 15332 2994
rect 15580 800 15608 3402
rect 15672 3058 15700 3470
rect 15948 3194 15976 3606
rect 15936 3188 15988 3194
rect 15936 3130 15988 3136
rect 15660 3052 15712 3058
rect 15660 2994 15712 3000
rect 15752 2372 15804 2378
rect 15752 2314 15804 2320
rect 15764 1170 15792 2314
rect 15764 1142 15884 1170
rect 15856 800 15884 1142
rect 16132 800 16160 4014
rect 16408 800 16436 4558
rect 16592 4282 16620 4558
rect 16580 4276 16632 4282
rect 16580 4218 16632 4224
rect 16580 3460 16632 3466
rect 16580 3402 16632 3408
rect 16592 2854 16620 3402
rect 16580 2848 16632 2854
rect 16580 2790 16632 2796
rect 16684 800 16712 4966
rect 16946 4856 17002 4865
rect 16946 4791 17002 4800
rect 16960 4146 16988 4791
rect 17236 4486 17264 6967
rect 17420 6798 17448 7822
rect 17512 7478 17540 7958
rect 17500 7472 17552 7478
rect 17500 7414 17552 7420
rect 17408 6792 17460 6798
rect 17408 6734 17460 6740
rect 17420 5778 17448 6734
rect 17512 6730 17540 7414
rect 17500 6724 17552 6730
rect 17500 6666 17552 6672
rect 17408 5772 17460 5778
rect 17408 5714 17460 5720
rect 17420 5234 17448 5714
rect 17408 5228 17460 5234
rect 17408 5170 17460 5176
rect 17500 4820 17552 4826
rect 17500 4762 17552 4768
rect 17316 4752 17368 4758
rect 17316 4694 17368 4700
rect 17328 4486 17356 4694
rect 17224 4480 17276 4486
rect 17224 4422 17276 4428
rect 17316 4480 17368 4486
rect 17316 4422 17368 4428
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 16764 3936 16816 3942
rect 16764 3878 16816 3884
rect 16776 2961 16804 3878
rect 17512 3534 17540 4762
rect 17604 4146 17632 7958
rect 17592 4140 17644 4146
rect 17592 4082 17644 4088
rect 17224 3528 17276 3534
rect 17224 3470 17276 3476
rect 17500 3528 17552 3534
rect 17500 3470 17552 3476
rect 16762 2952 16818 2961
rect 16762 2887 16818 2896
rect 16948 2916 17000 2922
rect 16948 2858 17000 2864
rect 16856 2848 16908 2854
rect 16856 2790 16908 2796
rect 16868 2514 16896 2790
rect 16856 2508 16908 2514
rect 16856 2450 16908 2456
rect 16960 800 16988 2858
rect 17236 800 17264 3470
rect 17696 3040 17724 10134
rect 17788 8022 17816 10367
rect 17880 10198 17908 11070
rect 17960 10736 18012 10742
rect 17960 10678 18012 10684
rect 17868 10192 17920 10198
rect 17868 10134 17920 10140
rect 17972 8566 18000 10678
rect 18052 8934 18104 8940
rect 18052 8876 18104 8882
rect 17960 8560 18012 8566
rect 17960 8502 18012 8508
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 17880 8362 17908 8434
rect 17868 8356 17920 8362
rect 17868 8298 17920 8304
rect 17776 8016 17828 8022
rect 17776 7958 17828 7964
rect 17880 7834 17908 8298
rect 17972 7886 18000 8502
rect 17788 7806 17908 7834
rect 17960 7880 18012 7886
rect 17960 7822 18012 7828
rect 17788 6798 17816 7806
rect 17960 7744 18012 7750
rect 17960 7686 18012 7692
rect 17868 7472 17920 7478
rect 17868 7414 17920 7420
rect 17972 7426 18000 7686
rect 18064 7546 18092 8876
rect 18052 7540 18104 7546
rect 18052 7482 18104 7488
rect 17880 7342 17908 7414
rect 17972 7398 18092 7426
rect 17868 7336 17920 7342
rect 17868 7278 17920 7284
rect 17776 6792 17828 6798
rect 17776 6734 17828 6740
rect 17880 6610 17908 7278
rect 18064 7274 18092 7398
rect 18052 7268 18104 7274
rect 18052 7210 18104 7216
rect 17960 6792 18012 6798
rect 17960 6734 18012 6740
rect 17788 6582 17908 6610
rect 17788 6390 17816 6582
rect 17868 6452 17920 6458
rect 17868 6394 17920 6400
rect 17776 6384 17828 6390
rect 17776 6326 17828 6332
rect 17788 5710 17816 6326
rect 17776 5704 17828 5710
rect 17776 5646 17828 5652
rect 17774 4992 17830 5001
rect 17774 4927 17830 4936
rect 17788 3466 17816 4927
rect 17880 4622 17908 6394
rect 17972 6322 18000 6734
rect 17960 6316 18012 6322
rect 17960 6258 18012 6264
rect 18064 5234 18092 7210
rect 18156 6934 18184 12174
rect 18144 6928 18196 6934
rect 18144 6870 18196 6876
rect 18144 6656 18196 6662
rect 18144 6598 18196 6604
rect 18156 5778 18184 6598
rect 18144 5772 18196 5778
rect 18144 5714 18196 5720
rect 18052 5228 18104 5234
rect 18052 5170 18104 5176
rect 17868 4616 17920 4622
rect 17868 4558 17920 4564
rect 18052 4548 18104 4554
rect 18052 4490 18104 4496
rect 17958 3904 18014 3913
rect 17958 3839 18014 3848
rect 17972 3738 18000 3839
rect 17960 3732 18012 3738
rect 17960 3674 18012 3680
rect 17776 3460 17828 3466
rect 17776 3402 17828 3408
rect 17776 3052 17828 3058
rect 17696 3012 17776 3040
rect 17776 2994 17828 3000
rect 18064 2938 18092 4490
rect 18144 3936 18196 3942
rect 18144 3878 18196 3884
rect 18156 3126 18184 3878
rect 18248 3126 18276 13806
rect 18340 4622 18368 15030
rect 18432 14822 18460 15302
rect 18420 14816 18472 14822
rect 18420 14758 18472 14764
rect 18694 13832 18750 13841
rect 18694 13767 18750 13776
rect 18420 13456 18472 13462
rect 18418 13424 18420 13433
rect 18472 13424 18474 13433
rect 18418 13359 18474 13368
rect 18708 12434 18736 13767
rect 18880 13524 18932 13530
rect 18880 13466 18932 13472
rect 18432 12406 18736 12434
rect 18328 4616 18380 4622
rect 18328 4558 18380 4564
rect 18432 3942 18460 12406
rect 18512 12368 18564 12374
rect 18512 12310 18564 12316
rect 18696 12368 18748 12374
rect 18696 12310 18748 12316
rect 18524 8401 18552 12310
rect 18708 12238 18736 12310
rect 18892 12238 18920 13466
rect 18696 12232 18748 12238
rect 18696 12174 18748 12180
rect 18880 12232 18932 12238
rect 18880 12174 18932 12180
rect 18708 11558 18736 12174
rect 18892 11830 18920 12174
rect 18972 12096 19024 12102
rect 18972 12038 19024 12044
rect 18880 11824 18932 11830
rect 18880 11766 18932 11772
rect 18984 11642 19012 12038
rect 18892 11626 19012 11642
rect 18880 11620 19012 11626
rect 18932 11614 19012 11620
rect 18880 11562 18932 11568
rect 18696 11552 18748 11558
rect 18696 11494 18748 11500
rect 18972 10600 19024 10606
rect 18892 10560 18972 10588
rect 18696 10124 18748 10130
rect 18696 10066 18748 10072
rect 18788 10124 18840 10130
rect 18788 10066 18840 10072
rect 18604 9716 18656 9722
rect 18604 9658 18656 9664
rect 18510 8392 18566 8401
rect 18510 8327 18566 8336
rect 18512 8288 18564 8294
rect 18512 8230 18564 8236
rect 18524 7750 18552 8230
rect 18512 7744 18564 7750
rect 18512 7686 18564 7692
rect 18616 7528 18644 9658
rect 18708 8022 18736 10066
rect 18800 9722 18828 10066
rect 18788 9716 18840 9722
rect 18788 9658 18840 9664
rect 18788 9512 18840 9518
rect 18788 9454 18840 9460
rect 18800 9042 18828 9454
rect 18788 9036 18840 9042
rect 18788 8978 18840 8984
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 18696 8016 18748 8022
rect 18696 7958 18748 7964
rect 18524 7500 18644 7528
rect 18524 6798 18552 7500
rect 18602 7440 18658 7449
rect 18602 7375 18658 7384
rect 18616 6866 18644 7375
rect 18604 6860 18656 6866
rect 18604 6802 18656 6808
rect 18512 6792 18564 6798
rect 18512 6734 18564 6740
rect 18512 6656 18564 6662
rect 18512 6598 18564 6604
rect 18604 6656 18656 6662
rect 18604 6598 18656 6604
rect 18524 6390 18552 6598
rect 18512 6384 18564 6390
rect 18512 6326 18564 6332
rect 18512 6248 18564 6254
rect 18512 6190 18564 6196
rect 18524 5574 18552 6190
rect 18616 5574 18644 6598
rect 18708 6186 18736 7958
rect 18800 6254 18828 8774
rect 18788 6248 18840 6254
rect 18788 6190 18840 6196
rect 18696 6180 18748 6186
rect 18696 6122 18748 6128
rect 18892 5681 18920 10560
rect 18972 10542 19024 10548
rect 18972 9920 19024 9926
rect 18972 9862 19024 9868
rect 18984 8362 19012 9862
rect 19076 8838 19104 22066
rect 19352 20992 19380 22442
rect 20260 22432 20312 22438
rect 20260 22374 20312 22380
rect 19720 21962 20116 21978
rect 20272 21962 20300 22374
rect 19432 21956 19484 21962
rect 19432 21898 19484 21904
rect 19708 21956 20116 21962
rect 19760 21950 20116 21956
rect 19708 21898 19760 21904
rect 19260 20964 19380 20992
rect 19444 20992 19472 21898
rect 19800 21888 19852 21894
rect 19852 21848 20024 21876
rect 19800 21830 19852 21836
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19996 21690 20024 21848
rect 19708 21684 19760 21690
rect 19708 21626 19760 21632
rect 19984 21684 20036 21690
rect 19984 21626 20036 21632
rect 19524 21004 19576 21010
rect 19444 20964 19524 20992
rect 19260 20482 19288 20964
rect 19340 20868 19392 20874
rect 19340 20810 19392 20816
rect 19352 20602 19380 20810
rect 19340 20596 19392 20602
rect 19340 20538 19392 20544
rect 19260 20466 19380 20482
rect 19260 20460 19392 20466
rect 19260 20454 19340 20460
rect 19340 20402 19392 20408
rect 19352 20210 19380 20402
rect 19444 20398 19472 20964
rect 19524 20946 19576 20952
rect 19720 20806 19748 21626
rect 20088 21622 20116 21950
rect 20260 21956 20312 21962
rect 20260 21898 20312 21904
rect 20168 21888 20220 21894
rect 20168 21830 20220 21836
rect 20076 21616 20128 21622
rect 20076 21558 20128 21564
rect 19984 21344 20036 21350
rect 19984 21286 20036 21292
rect 20076 21344 20128 21350
rect 20076 21286 20128 21292
rect 19708 20800 19760 20806
rect 19708 20742 19760 20748
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19800 20596 19852 20602
rect 19800 20538 19852 20544
rect 19432 20392 19484 20398
rect 19432 20334 19484 20340
rect 19812 20262 19840 20538
rect 19800 20256 19852 20262
rect 19352 20182 19472 20210
rect 19800 20198 19852 20204
rect 19156 19984 19208 19990
rect 19156 19926 19208 19932
rect 19168 19378 19196 19926
rect 19340 19712 19392 19718
rect 19340 19654 19392 19660
rect 19156 19372 19208 19378
rect 19156 19314 19208 19320
rect 19248 18284 19300 18290
rect 19248 18226 19300 18232
rect 19260 16114 19288 18226
rect 19352 17882 19380 19654
rect 19444 18902 19472 20182
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19432 18896 19484 18902
rect 19432 18838 19484 18844
rect 19444 18306 19472 18838
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19444 18278 19564 18306
rect 19432 18216 19484 18222
rect 19432 18158 19484 18164
rect 19340 17876 19392 17882
rect 19340 17818 19392 17824
rect 19444 16250 19472 18158
rect 19536 17678 19564 18278
rect 19708 17876 19760 17882
rect 19708 17818 19760 17824
rect 19524 17672 19576 17678
rect 19524 17614 19576 17620
rect 19720 17610 19748 17818
rect 19996 17678 20024 21286
rect 20088 20874 20116 21286
rect 20180 20942 20208 21830
rect 20168 20936 20220 20942
rect 20168 20878 20220 20884
rect 20076 20868 20128 20874
rect 20076 20810 20128 20816
rect 20260 20800 20312 20806
rect 20260 20742 20312 20748
rect 20076 20256 20128 20262
rect 20076 20198 20128 20204
rect 19984 17672 20036 17678
rect 19984 17614 20036 17620
rect 19708 17604 19760 17610
rect 19708 17546 19760 17552
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 20088 16590 20116 20198
rect 20168 19712 20220 19718
rect 20168 19654 20220 19660
rect 20180 19378 20208 19654
rect 20168 19372 20220 19378
rect 20168 19314 20220 19320
rect 20076 16584 20128 16590
rect 20076 16526 20128 16532
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19432 16244 19484 16250
rect 19432 16186 19484 16192
rect 19340 16176 19392 16182
rect 19340 16118 19392 16124
rect 19248 16108 19300 16114
rect 19248 16050 19300 16056
rect 19248 15428 19300 15434
rect 19248 15370 19300 15376
rect 19156 15360 19208 15366
rect 19156 15302 19208 15308
rect 19168 12442 19196 15302
rect 19260 14958 19288 15370
rect 19248 14952 19300 14958
rect 19248 14894 19300 14900
rect 19248 14476 19300 14482
rect 19248 14418 19300 14424
rect 19260 13410 19288 14418
rect 19352 13530 19380 16118
rect 19432 16040 19484 16046
rect 19432 15982 19484 15988
rect 19444 14890 19472 15982
rect 19616 15904 19668 15910
rect 19616 15846 19668 15852
rect 20076 15904 20128 15910
rect 20076 15846 20128 15852
rect 19628 15502 19656 15846
rect 19616 15496 19668 15502
rect 20088 15484 20116 15846
rect 20272 15638 20300 20742
rect 20260 15632 20312 15638
rect 20260 15574 20312 15580
rect 20168 15496 20220 15502
rect 20088 15456 20168 15484
rect 19616 15438 19668 15444
rect 20168 15438 20220 15444
rect 20076 15360 20128 15366
rect 20076 15302 20128 15308
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 20088 15094 20116 15302
rect 20076 15088 20128 15094
rect 20076 15030 20128 15036
rect 19432 14884 19484 14890
rect 19432 14826 19484 14832
rect 19524 14816 19576 14822
rect 19524 14758 19576 14764
rect 19432 14612 19484 14618
rect 19432 14554 19484 14560
rect 19444 13734 19472 14554
rect 19536 14550 19564 14758
rect 19524 14544 19576 14550
rect 19524 14486 19576 14492
rect 19800 14408 19852 14414
rect 19614 14376 19670 14385
rect 19852 14356 20116 14362
rect 19800 14350 20116 14356
rect 19812 14334 20116 14350
rect 19614 14311 19616 14320
rect 19668 14311 19670 14320
rect 19616 14282 19668 14288
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19432 13728 19484 13734
rect 19432 13670 19484 13676
rect 19340 13524 19392 13530
rect 19340 13466 19392 13472
rect 19800 13524 19852 13530
rect 19800 13466 19852 13472
rect 19260 13382 19380 13410
rect 19156 12436 19208 12442
rect 19156 12378 19208 12384
rect 19156 11688 19208 11694
rect 19156 11630 19208 11636
rect 19246 11656 19302 11665
rect 19168 10062 19196 11630
rect 19246 11591 19248 11600
rect 19300 11591 19302 11600
rect 19248 11562 19300 11568
rect 19352 11354 19380 13382
rect 19432 13252 19484 13258
rect 19432 13194 19484 13200
rect 19444 12968 19472 13194
rect 19812 13190 19840 13466
rect 20088 13394 20116 14334
rect 20076 13388 20128 13394
rect 20076 13330 20128 13336
rect 19800 13184 19852 13190
rect 19800 13126 19852 13132
rect 19984 13184 20036 13190
rect 20036 13144 20116 13172
rect 19984 13126 20036 13132
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19444 12940 19564 12968
rect 19536 12714 19564 12940
rect 19616 12912 19668 12918
rect 19616 12854 19668 12860
rect 19432 12708 19484 12714
rect 19432 12650 19484 12656
rect 19524 12708 19576 12714
rect 19524 12650 19576 12656
rect 19444 12374 19472 12650
rect 19522 12608 19578 12617
rect 19522 12543 19578 12552
rect 19432 12368 19484 12374
rect 19432 12310 19484 12316
rect 19444 12238 19472 12310
rect 19432 12232 19484 12238
rect 19432 12174 19484 12180
rect 19536 12084 19564 12543
rect 19628 12238 19656 12854
rect 19616 12232 19668 12238
rect 19616 12174 19668 12180
rect 19984 12164 20036 12170
rect 19984 12106 20036 12112
rect 19444 12056 19564 12084
rect 19444 11898 19472 12056
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19996 11937 20024 12106
rect 19982 11928 20038 11937
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 19892 11892 19944 11898
rect 20088 11898 20116 13144
rect 20180 12617 20208 15438
rect 20166 12608 20222 12617
rect 20166 12543 20222 12552
rect 20364 11914 20392 30602
rect 20456 28422 20484 31726
rect 20444 28416 20496 28422
rect 20444 28358 20496 28364
rect 20732 27146 20760 36178
rect 21008 34474 21036 36246
rect 21100 35698 21128 37266
rect 21088 35692 21140 35698
rect 21088 35634 21140 35640
rect 20996 34468 21048 34474
rect 20996 34410 21048 34416
rect 21008 33504 21036 34410
rect 21284 33930 21312 37674
rect 21376 33998 21404 60182
rect 21836 60110 21864 60302
rect 22098 60279 22154 60288
rect 22098 60208 22154 60217
rect 22098 60143 22154 60152
rect 22112 60110 22140 60143
rect 22480 60110 22508 60454
rect 22572 60353 22600 60658
rect 22558 60344 22614 60353
rect 22558 60279 22614 60288
rect 22652 60240 22704 60246
rect 22652 60182 22704 60188
rect 21824 60104 21876 60110
rect 21824 60046 21876 60052
rect 22008 60104 22060 60110
rect 22008 60046 22060 60052
rect 22100 60104 22152 60110
rect 22100 60046 22152 60052
rect 22376 60104 22428 60110
rect 22376 60046 22428 60052
rect 22468 60104 22520 60110
rect 22468 60046 22520 60052
rect 21640 59968 21692 59974
rect 21640 59910 21692 59916
rect 21456 59696 21508 59702
rect 21456 59638 21508 59644
rect 21468 59430 21496 59638
rect 21456 59424 21508 59430
rect 21456 59366 21508 59372
rect 21468 59022 21496 59366
rect 21456 59016 21508 59022
rect 21456 58958 21508 58964
rect 21468 44334 21496 58958
rect 21456 44328 21508 44334
rect 21456 44270 21508 44276
rect 21364 33992 21416 33998
rect 21364 33934 21416 33940
rect 21272 33924 21324 33930
rect 21272 33866 21324 33872
rect 21088 33516 21140 33522
rect 21008 33476 21088 33504
rect 21088 33458 21140 33464
rect 20904 33312 20956 33318
rect 20904 33254 20956 33260
rect 20916 33114 20944 33254
rect 20904 33108 20956 33114
rect 20904 33050 20956 33056
rect 21284 31278 21312 33866
rect 21468 33590 21496 44270
rect 21548 34128 21600 34134
rect 21546 34096 21548 34105
rect 21600 34096 21602 34105
rect 21546 34031 21602 34040
rect 21548 33992 21600 33998
rect 21548 33934 21600 33940
rect 21456 33584 21508 33590
rect 21456 33526 21508 33532
rect 21468 33425 21496 33526
rect 21454 33416 21510 33425
rect 21454 33351 21510 33360
rect 21272 31272 21324 31278
rect 21272 31214 21324 31220
rect 21560 29730 21588 33934
rect 21652 30190 21680 59910
rect 22020 59673 22048 60046
rect 22006 59664 22062 59673
rect 22006 59599 22062 59608
rect 22100 59628 22152 59634
rect 22100 59570 22152 59576
rect 22112 56914 22140 59570
rect 22388 59498 22416 60046
rect 22376 59492 22428 59498
rect 22376 59434 22428 59440
rect 22100 56908 22152 56914
rect 22100 56850 22152 56856
rect 22468 40452 22520 40458
rect 22468 40394 22520 40400
rect 21732 39840 21784 39846
rect 21732 39782 21784 39788
rect 21744 38350 21772 39782
rect 22284 39568 22336 39574
rect 22284 39510 22336 39516
rect 21732 38344 21784 38350
rect 21732 38286 21784 38292
rect 21824 38208 21876 38214
rect 21824 38150 21876 38156
rect 22008 38208 22060 38214
rect 22008 38150 22060 38156
rect 21732 34196 21784 34202
rect 21732 34138 21784 34144
rect 21744 33114 21772 34138
rect 21732 33108 21784 33114
rect 21732 33050 21784 33056
rect 21744 31754 21772 33050
rect 21836 32910 21864 38150
rect 21916 37256 21968 37262
rect 21916 37198 21968 37204
rect 21824 32904 21876 32910
rect 21824 32846 21876 32852
rect 21732 31748 21784 31754
rect 21732 31690 21784 31696
rect 21824 31204 21876 31210
rect 21824 31146 21876 31152
rect 21640 30184 21692 30190
rect 21640 30126 21692 30132
rect 21560 29702 21680 29730
rect 21548 29640 21600 29646
rect 21548 29582 21600 29588
rect 21560 29306 21588 29582
rect 21548 29300 21600 29306
rect 21548 29242 21600 29248
rect 20732 27118 20852 27146
rect 20720 26920 20772 26926
rect 20720 26862 20772 26868
rect 20732 25265 20760 26862
rect 20718 25256 20774 25265
rect 20718 25191 20774 25200
rect 20824 22506 20852 27118
rect 21652 22710 21680 29702
rect 21836 29578 21864 31146
rect 21928 29646 21956 37198
rect 22020 32434 22048 38150
rect 22192 36168 22244 36174
rect 22192 36110 22244 36116
rect 22204 35562 22232 36110
rect 22192 35556 22244 35562
rect 22192 35498 22244 35504
rect 22296 35086 22324 39510
rect 22480 36174 22508 40394
rect 22560 37800 22612 37806
rect 22558 37768 22560 37777
rect 22612 37768 22614 37777
rect 22558 37703 22614 37712
rect 22468 36168 22520 36174
rect 22468 36110 22520 36116
rect 22284 35080 22336 35086
rect 22284 35022 22336 35028
rect 22376 34672 22428 34678
rect 22376 34614 22428 34620
rect 22192 34128 22244 34134
rect 22192 34070 22244 34076
rect 22204 33522 22232 34070
rect 22284 33652 22336 33658
rect 22284 33594 22336 33600
rect 22192 33516 22244 33522
rect 22192 33458 22244 33464
rect 22192 32836 22244 32842
rect 22192 32778 22244 32784
rect 22100 32768 22152 32774
rect 22100 32710 22152 32716
rect 22008 32428 22060 32434
rect 22008 32370 22060 32376
rect 21916 29640 21968 29646
rect 21916 29582 21968 29588
rect 21824 29572 21876 29578
rect 21824 29514 21876 29520
rect 21732 29164 21784 29170
rect 21732 29106 21784 29112
rect 21640 22704 21692 22710
rect 21640 22646 21692 22652
rect 20812 22500 20864 22506
rect 20812 22442 20864 22448
rect 20996 22160 21048 22166
rect 20996 22102 21048 22108
rect 21008 22030 21036 22102
rect 20996 22024 21048 22030
rect 20996 21966 21048 21972
rect 21456 21684 21508 21690
rect 21456 21626 21508 21632
rect 20812 21616 20864 21622
rect 20812 21558 20864 21564
rect 20824 20058 20852 21558
rect 21468 20466 21496 21626
rect 21456 20460 21508 20466
rect 21456 20402 21508 20408
rect 20812 20052 20864 20058
rect 20812 19994 20864 20000
rect 21468 19990 21496 20402
rect 21456 19984 21508 19990
rect 21456 19926 21508 19932
rect 20812 19848 20864 19854
rect 20812 19790 20864 19796
rect 20720 19304 20772 19310
rect 20720 19246 20772 19252
rect 20732 17202 20760 19246
rect 20824 18902 20852 19790
rect 21468 19242 21496 19926
rect 21456 19236 21508 19242
rect 21456 19178 21508 19184
rect 20812 18896 20864 18902
rect 20812 18838 20864 18844
rect 20996 18692 21048 18698
rect 20996 18634 21048 18640
rect 20902 18592 20958 18601
rect 20902 18527 20958 18536
rect 20916 18426 20944 18527
rect 21008 18426 21036 18634
rect 20904 18420 20956 18426
rect 20904 18362 20956 18368
rect 20996 18420 21048 18426
rect 20996 18362 21048 18368
rect 21638 18320 21694 18329
rect 21638 18255 21640 18264
rect 21692 18255 21694 18264
rect 21640 18226 21692 18232
rect 21272 17332 21324 17338
rect 21272 17274 21324 17280
rect 21284 17202 21312 17274
rect 20720 17196 20772 17202
rect 20720 17138 20772 17144
rect 21088 17196 21140 17202
rect 21088 17138 21140 17144
rect 21272 17196 21324 17202
rect 21272 17138 21324 17144
rect 20996 17128 21048 17134
rect 20996 17070 21048 17076
rect 20444 17060 20496 17066
rect 20444 17002 20496 17008
rect 20456 16250 20484 17002
rect 21008 16998 21036 17070
rect 20996 16992 21048 16998
rect 20996 16934 21048 16940
rect 20444 16244 20496 16250
rect 20444 16186 20496 16192
rect 20718 16008 20774 16017
rect 20718 15943 20774 15952
rect 20904 15972 20956 15978
rect 20442 15192 20498 15201
rect 20442 15127 20498 15136
rect 19982 11863 20038 11872
rect 20076 11892 20128 11898
rect 19892 11834 19944 11840
rect 20076 11834 20128 11840
rect 20272 11886 20392 11914
rect 19800 11756 19852 11762
rect 19800 11698 19852 11704
rect 19812 11665 19840 11698
rect 19798 11656 19854 11665
rect 19708 11620 19760 11626
rect 19798 11591 19854 11600
rect 19708 11562 19760 11568
rect 19524 11552 19576 11558
rect 19524 11494 19576 11500
rect 19340 11348 19392 11354
rect 19340 11290 19392 11296
rect 19536 11218 19564 11494
rect 19720 11393 19748 11562
rect 19706 11384 19762 11393
rect 19706 11319 19762 11328
rect 19524 11212 19576 11218
rect 19524 11154 19576 11160
rect 19904 11150 19932 11834
rect 20088 11626 20116 11834
rect 20272 11778 20300 11886
rect 20180 11750 20300 11778
rect 20076 11620 20128 11626
rect 20076 11562 20128 11568
rect 20074 11520 20130 11529
rect 20074 11455 20130 11464
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19892 11144 19944 11150
rect 19892 11086 19944 11092
rect 19444 10606 19472 11086
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19614 10704 19670 10713
rect 19614 10639 19670 10648
rect 19432 10600 19484 10606
rect 19432 10542 19484 10548
rect 19340 10192 19392 10198
rect 19340 10134 19392 10140
rect 19156 10056 19208 10062
rect 19156 9998 19208 10004
rect 19156 9512 19208 9518
rect 19156 9454 19208 9460
rect 19168 9081 19196 9454
rect 19246 9344 19302 9353
rect 19246 9279 19302 9288
rect 19154 9072 19210 9081
rect 19154 9007 19210 9016
rect 19064 8832 19116 8838
rect 19064 8774 19116 8780
rect 19154 8800 19210 8809
rect 19154 8735 19210 8744
rect 19168 8634 19196 8735
rect 19260 8634 19288 9279
rect 19156 8628 19208 8634
rect 19156 8570 19208 8576
rect 19248 8628 19300 8634
rect 19248 8570 19300 8576
rect 19352 8480 19380 10134
rect 19444 10062 19472 10542
rect 19524 10532 19576 10538
rect 19524 10474 19576 10480
rect 19536 10266 19564 10474
rect 19524 10260 19576 10266
rect 19524 10202 19576 10208
rect 19432 10056 19484 10062
rect 19432 9998 19484 10004
rect 19444 9518 19472 9998
rect 19628 9994 19656 10639
rect 19798 10296 19854 10305
rect 19798 10231 19854 10240
rect 19812 10198 19840 10231
rect 19800 10192 19852 10198
rect 19800 10134 19852 10140
rect 19616 9988 19668 9994
rect 19616 9930 19668 9936
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19432 9512 19484 9518
rect 19432 9454 19484 9460
rect 19444 8616 19472 9454
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19892 8628 19944 8634
rect 19444 8588 19564 8616
rect 19352 8452 19472 8480
rect 19444 8378 19472 8452
rect 18972 8356 19024 8362
rect 18972 8298 19024 8304
rect 19352 8350 19472 8378
rect 19064 8288 19116 8294
rect 19248 8288 19300 8294
rect 19064 8230 19116 8236
rect 19168 8236 19248 8242
rect 19168 8230 19300 8236
rect 19076 8106 19104 8230
rect 18984 8078 19104 8106
rect 19168 8214 19288 8230
rect 18984 7585 19012 8078
rect 19168 8022 19196 8214
rect 19156 8016 19208 8022
rect 19156 7958 19208 7964
rect 19064 7880 19116 7886
rect 19064 7822 19116 7828
rect 18970 7576 19026 7585
rect 18970 7511 19026 7520
rect 19076 7478 19104 7822
rect 19352 7750 19380 8350
rect 19536 8294 19564 8588
rect 19892 8570 19944 8576
rect 19904 8362 19932 8570
rect 19984 8424 20036 8430
rect 19984 8366 20036 8372
rect 19892 8356 19944 8362
rect 19892 8298 19944 8304
rect 19444 8266 19564 8294
rect 19444 7954 19472 8266
rect 19996 8129 20024 8366
rect 19982 8120 20038 8129
rect 19982 8055 20038 8064
rect 19432 7948 19484 7954
rect 19432 7890 19484 7896
rect 19340 7744 19392 7750
rect 19154 7712 19210 7721
rect 19340 7686 19392 7692
rect 19154 7647 19210 7656
rect 19168 7562 19196 7647
rect 19168 7534 19380 7562
rect 19064 7472 19116 7478
rect 19064 7414 19116 7420
rect 18972 7404 19024 7410
rect 18972 7346 19024 7352
rect 18984 6866 19012 7346
rect 19064 7336 19116 7342
rect 19064 7278 19116 7284
rect 19154 7304 19210 7313
rect 19076 7177 19104 7278
rect 19154 7239 19156 7248
rect 19208 7239 19210 7248
rect 19156 7210 19208 7216
rect 19062 7168 19118 7177
rect 19062 7103 19118 7112
rect 18972 6860 19024 6866
rect 18972 6802 19024 6808
rect 18984 5710 19012 6802
rect 19352 6798 19380 7534
rect 19444 7410 19472 7890
rect 19984 7880 20036 7886
rect 19984 7822 20036 7828
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19524 7472 19576 7478
rect 19522 7440 19524 7449
rect 19576 7440 19578 7449
rect 19432 7404 19484 7410
rect 19522 7375 19578 7384
rect 19432 7346 19484 7352
rect 19340 6792 19392 6798
rect 19340 6734 19392 6740
rect 19444 6780 19472 7346
rect 19892 7336 19944 7342
rect 19890 7304 19892 7313
rect 19944 7304 19946 7313
rect 19996 7274 20024 7822
rect 19890 7239 19946 7248
rect 19984 7268 20036 7274
rect 19984 7210 20036 7216
rect 19616 6792 19668 6798
rect 19444 6752 19616 6780
rect 19248 6316 19300 6322
rect 19248 6258 19300 6264
rect 19340 6316 19392 6322
rect 19340 6258 19392 6264
rect 19062 6216 19118 6225
rect 19062 6151 19118 6160
rect 18972 5704 19024 5710
rect 18878 5672 18934 5681
rect 18972 5646 19024 5652
rect 18878 5607 18934 5616
rect 18512 5568 18564 5574
rect 18512 5510 18564 5516
rect 18604 5568 18656 5574
rect 18604 5510 18656 5516
rect 18616 5370 18644 5510
rect 18604 5364 18656 5370
rect 18604 5306 18656 5312
rect 18970 4720 19026 4729
rect 18880 4684 18932 4690
rect 18970 4655 18972 4664
rect 18880 4626 18932 4632
rect 19024 4655 19026 4664
rect 18972 4626 19024 4632
rect 18604 4140 18656 4146
rect 18604 4082 18656 4088
rect 18512 4072 18564 4078
rect 18512 4014 18564 4020
rect 18420 3936 18472 3942
rect 18420 3878 18472 3884
rect 18524 3738 18552 4014
rect 18512 3732 18564 3738
rect 18512 3674 18564 3680
rect 18418 3632 18474 3641
rect 18418 3567 18474 3576
rect 18432 3534 18460 3567
rect 18420 3528 18472 3534
rect 18420 3470 18472 3476
rect 18144 3120 18196 3126
rect 18144 3062 18196 3068
rect 18236 3120 18288 3126
rect 18236 3062 18288 3068
rect 17960 2916 18012 2922
rect 18064 2910 18368 2938
rect 17960 2858 18012 2864
rect 17972 2774 18000 2858
rect 17972 2746 18092 2774
rect 17498 2680 17554 2689
rect 17408 2644 17460 2650
rect 17498 2615 17554 2624
rect 17408 2586 17460 2592
rect 17316 2440 17368 2446
rect 17316 2382 17368 2388
rect 17328 1766 17356 2382
rect 17316 1760 17368 1766
rect 17316 1702 17368 1708
rect 17420 1306 17448 2586
rect 17512 2446 17540 2615
rect 17776 2508 17828 2514
rect 17776 2450 17828 2456
rect 17500 2440 17552 2446
rect 17500 2382 17552 2388
rect 17420 1278 17540 1306
rect 17512 800 17540 1278
rect 17788 800 17816 2450
rect 18064 800 18092 2746
rect 18340 800 18368 2910
rect 18420 2440 18472 2446
rect 18420 2382 18472 2388
rect 18432 2038 18460 2382
rect 18420 2032 18472 2038
rect 18420 1974 18472 1980
rect 18616 800 18644 4082
rect 18788 3936 18840 3942
rect 18788 3878 18840 3884
rect 18800 3466 18828 3878
rect 18788 3460 18840 3466
rect 18788 3402 18840 3408
rect 18892 800 18920 4626
rect 19076 4146 19104 6151
rect 19260 5250 19288 6258
rect 19352 5370 19380 6258
rect 19444 6254 19472 6752
rect 19616 6734 19668 6740
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19524 6384 19576 6390
rect 19524 6326 19576 6332
rect 19800 6384 19852 6390
rect 19800 6326 19852 6332
rect 19432 6248 19484 6254
rect 19432 6190 19484 6196
rect 19444 5710 19472 6190
rect 19536 5817 19564 6326
rect 19616 5840 19668 5846
rect 19522 5808 19578 5817
rect 19812 5828 19840 6326
rect 19668 5800 19840 5828
rect 19616 5782 19668 5788
rect 19522 5743 19578 5752
rect 19432 5704 19484 5710
rect 19432 5646 19484 5652
rect 19616 5704 19668 5710
rect 19668 5664 20024 5692
rect 19616 5646 19668 5652
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19340 5364 19392 5370
rect 19340 5306 19392 5312
rect 19430 5264 19486 5273
rect 19260 5234 19380 5250
rect 19260 5228 19392 5234
rect 19260 5222 19340 5228
rect 19430 5199 19486 5208
rect 19340 5170 19392 5176
rect 19444 4706 19472 5199
rect 19892 5160 19944 5166
rect 19892 5102 19944 5108
rect 19904 4758 19932 5102
rect 19352 4678 19472 4706
rect 19892 4752 19944 4758
rect 19892 4694 19944 4700
rect 19352 4457 19380 4678
rect 19432 4616 19484 4622
rect 19430 4584 19432 4593
rect 19484 4584 19486 4593
rect 19430 4519 19486 4528
rect 19890 4584 19946 4593
rect 19890 4519 19892 4528
rect 19944 4519 19946 4528
rect 19892 4490 19944 4496
rect 19338 4448 19394 4457
rect 19338 4383 19394 4392
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19338 4312 19394 4321
rect 19574 4315 19882 4324
rect 19338 4247 19340 4256
rect 19392 4247 19394 4256
rect 19340 4218 19392 4224
rect 19524 4208 19576 4214
rect 19522 4176 19524 4185
rect 19576 4176 19578 4185
rect 19064 4140 19116 4146
rect 19522 4111 19578 4120
rect 19616 4140 19668 4146
rect 19064 4082 19116 4088
rect 19800 4140 19852 4146
rect 19668 4100 19800 4128
rect 19616 4082 19668 4088
rect 19800 4082 19852 4088
rect 19996 4078 20024 5664
rect 20088 4622 20116 11455
rect 20180 7750 20208 11750
rect 20352 11620 20404 11626
rect 20352 11562 20404 11568
rect 20364 11354 20392 11562
rect 20260 11348 20312 11354
rect 20260 11290 20312 11296
rect 20352 11348 20404 11354
rect 20352 11290 20404 11296
rect 20272 8362 20300 11290
rect 20350 8664 20406 8673
rect 20350 8599 20406 8608
rect 20364 8498 20392 8599
rect 20352 8492 20404 8498
rect 20352 8434 20404 8440
rect 20260 8356 20312 8362
rect 20260 8298 20312 8304
rect 20456 7834 20484 15127
rect 20628 14816 20680 14822
rect 20628 14758 20680 14764
rect 20536 12300 20588 12306
rect 20536 12242 20588 12248
rect 20548 11762 20576 12242
rect 20536 11756 20588 11762
rect 20536 11698 20588 11704
rect 20640 11370 20668 14758
rect 20732 14657 20760 15943
rect 20904 15914 20956 15920
rect 20916 15745 20944 15914
rect 20902 15736 20958 15745
rect 20902 15671 20958 15680
rect 20718 14648 20774 14657
rect 20718 14583 20774 14592
rect 20812 14544 20864 14550
rect 20812 14486 20864 14492
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 20732 13530 20760 13874
rect 20824 13870 20852 14486
rect 20904 14272 20956 14278
rect 20904 14214 20956 14220
rect 20812 13864 20864 13870
rect 20812 13806 20864 13812
rect 20720 13524 20772 13530
rect 20720 13466 20772 13472
rect 20916 12782 20944 14214
rect 20812 12776 20864 12782
rect 20812 12718 20864 12724
rect 20904 12776 20956 12782
rect 20904 12718 20956 12724
rect 20824 11626 20852 12718
rect 20904 12232 20956 12238
rect 20904 12174 20956 12180
rect 20916 12102 20944 12174
rect 20904 12096 20956 12102
rect 20904 12038 20956 12044
rect 20904 11892 20956 11898
rect 20904 11834 20956 11840
rect 20812 11620 20864 11626
rect 20812 11562 20864 11568
rect 20640 11342 20760 11370
rect 20628 11280 20680 11286
rect 20548 11240 20628 11268
rect 20548 10674 20576 11240
rect 20628 11222 20680 11228
rect 20732 11098 20760 11342
rect 20640 11070 20760 11098
rect 20640 10742 20668 11070
rect 20628 10736 20680 10742
rect 20916 10690 20944 11834
rect 20628 10678 20680 10684
rect 20536 10668 20588 10674
rect 20536 10610 20588 10616
rect 20732 10662 20944 10690
rect 20732 10588 20760 10662
rect 20640 10560 20760 10588
rect 20536 9920 20588 9926
rect 20536 9862 20588 9868
rect 20272 7806 20484 7834
rect 20168 7744 20220 7750
rect 20168 7686 20220 7692
rect 20272 7562 20300 7806
rect 20352 7744 20404 7750
rect 20352 7686 20404 7692
rect 20180 7534 20300 7562
rect 20076 4616 20128 4622
rect 20076 4558 20128 4564
rect 19432 4072 19484 4078
rect 19430 4040 19432 4049
rect 19984 4072 20036 4078
rect 19484 4040 19486 4049
rect 18972 4004 19024 4010
rect 19984 4014 20036 4020
rect 19430 3975 19486 3984
rect 18972 3946 19024 3952
rect 18984 3602 19012 3946
rect 19432 3936 19484 3942
rect 19260 3896 19380 3924
rect 19260 3738 19288 3896
rect 19248 3732 19300 3738
rect 19248 3674 19300 3680
rect 18972 3596 19024 3602
rect 18972 3538 19024 3544
rect 19156 2848 19208 2854
rect 19156 2790 19208 2796
rect 19168 800 19196 2790
rect 19352 1986 19380 3896
rect 19616 3936 19668 3942
rect 19484 3884 19616 3890
rect 19432 3878 19668 3884
rect 19444 3862 19656 3878
rect 19522 3632 19578 3641
rect 19522 3567 19524 3576
rect 19576 3567 19578 3576
rect 19996 3584 20024 4014
rect 19996 3556 20116 3584
rect 19524 3538 19576 3544
rect 19904 3466 20024 3482
rect 20088 3466 20116 3556
rect 19904 3460 20036 3466
rect 19904 3454 19984 3460
rect 19524 3392 19576 3398
rect 19904 3380 19932 3454
rect 19984 3402 20036 3408
rect 20076 3460 20128 3466
rect 20076 3402 20128 3408
rect 19576 3352 19932 3380
rect 19524 3334 19576 3340
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19708 3052 19760 3058
rect 20088 3040 20116 3402
rect 19760 3012 20116 3040
rect 19708 2994 19760 3000
rect 19524 2916 19576 2922
rect 19524 2858 19576 2864
rect 19536 2650 19564 2858
rect 19890 2680 19946 2689
rect 19432 2644 19484 2650
rect 19432 2586 19484 2592
rect 19524 2644 19576 2650
rect 19890 2615 19946 2624
rect 19524 2586 19576 2592
rect 19444 2530 19472 2586
rect 19444 2502 19564 2530
rect 19536 2310 19564 2502
rect 19904 2446 19932 2615
rect 19892 2440 19944 2446
rect 19892 2382 19944 2388
rect 20076 2372 20128 2378
rect 20076 2314 20128 2320
rect 19432 2304 19484 2310
rect 19432 2246 19484 2252
rect 19524 2304 19576 2310
rect 19524 2246 19576 2252
rect 19444 2106 19472 2246
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19432 2100 19484 2106
rect 19432 2042 19484 2048
rect 19706 2000 19762 2009
rect 19352 1958 19472 1986
rect 19444 800 19472 1958
rect 19706 1935 19762 1944
rect 19720 800 19748 1935
rect 20088 1170 20116 2314
rect 20180 1766 20208 7534
rect 20364 7426 20392 7686
rect 20364 7398 20484 7426
rect 20260 5704 20312 5710
rect 20260 5646 20312 5652
rect 20272 5234 20300 5646
rect 20260 5228 20312 5234
rect 20260 5170 20312 5176
rect 20352 3732 20404 3738
rect 20352 3674 20404 3680
rect 20260 2848 20312 2854
rect 20260 2790 20312 2796
rect 20168 1760 20220 1766
rect 20168 1702 20220 1708
rect 19996 1142 20116 1170
rect 19996 800 20024 1142
rect 20272 800 20300 2790
rect 20364 1714 20392 3674
rect 20456 2310 20484 7398
rect 20548 7002 20576 9862
rect 20536 6996 20588 7002
rect 20536 6938 20588 6944
rect 20640 6225 20668 10560
rect 21008 10062 21036 16934
rect 21100 16522 21128 17138
rect 21088 16516 21140 16522
rect 21088 16458 21140 16464
rect 21100 15978 21128 16458
rect 21180 16108 21232 16114
rect 21180 16050 21232 16056
rect 21456 16108 21508 16114
rect 21456 16050 21508 16056
rect 21088 15972 21140 15978
rect 21088 15914 21140 15920
rect 21100 15502 21128 15914
rect 21088 15496 21140 15502
rect 21088 15438 21140 15444
rect 21088 14272 21140 14278
rect 21088 14214 21140 14220
rect 21100 14074 21128 14214
rect 21088 14068 21140 14074
rect 21088 14010 21140 14016
rect 21100 13326 21128 14010
rect 21088 13320 21140 13326
rect 21088 13262 21140 13268
rect 21088 13184 21140 13190
rect 21088 13126 21140 13132
rect 21100 11914 21128 13126
rect 21192 12434 21220 16050
rect 21468 15638 21496 16050
rect 21546 15872 21602 15881
rect 21546 15807 21602 15816
rect 21456 15632 21508 15638
rect 21456 15574 21508 15580
rect 21454 14376 21510 14385
rect 21454 14311 21456 14320
rect 21508 14311 21510 14320
rect 21456 14282 21508 14288
rect 21468 13938 21496 14282
rect 21456 13932 21508 13938
rect 21456 13874 21508 13880
rect 21456 12640 21508 12646
rect 21456 12582 21508 12588
rect 21192 12406 21404 12434
rect 21270 12200 21326 12209
rect 21270 12135 21326 12144
rect 21100 11886 21220 11914
rect 21088 11824 21140 11830
rect 21088 11766 21140 11772
rect 21100 11354 21128 11766
rect 21088 11348 21140 11354
rect 21088 11290 21140 11296
rect 21192 10470 21220 11886
rect 21180 10464 21232 10470
rect 21100 10412 21180 10418
rect 21100 10406 21232 10412
rect 21100 10390 21220 10406
rect 21100 10266 21128 10390
rect 21088 10260 21140 10266
rect 21088 10202 21140 10208
rect 20996 10056 21048 10062
rect 20996 9998 21048 10004
rect 21180 9580 21232 9586
rect 21180 9522 21232 9528
rect 21088 9512 21140 9518
rect 21088 9454 21140 9460
rect 21100 9382 21128 9454
rect 21088 9376 21140 9382
rect 21088 9318 21140 9324
rect 21100 9178 21128 9318
rect 21088 9172 21140 9178
rect 21088 9114 21140 9120
rect 21192 8838 21220 9522
rect 21284 9178 21312 12135
rect 21272 9172 21324 9178
rect 21272 9114 21324 9120
rect 21180 8832 21232 8838
rect 21180 8774 21232 8780
rect 21086 8392 21142 8401
rect 21086 8327 21142 8336
rect 20812 8288 20864 8294
rect 20812 8230 20864 8236
rect 20824 8022 20852 8230
rect 20812 8016 20864 8022
rect 20812 7958 20864 7964
rect 20720 7948 20772 7954
rect 20720 7890 20772 7896
rect 20732 6934 20760 7890
rect 21100 7274 21128 8327
rect 21180 7404 21232 7410
rect 21180 7346 21232 7352
rect 21088 7268 21140 7274
rect 21088 7210 21140 7216
rect 21192 7002 21220 7346
rect 21272 7200 21324 7206
rect 21272 7142 21324 7148
rect 21284 7002 21312 7142
rect 21180 6996 21232 7002
rect 21180 6938 21232 6944
rect 21272 6996 21324 7002
rect 21272 6938 21324 6944
rect 20720 6928 20772 6934
rect 20720 6870 20772 6876
rect 21180 6860 21232 6866
rect 21180 6802 21232 6808
rect 21192 6730 21220 6802
rect 21180 6724 21232 6730
rect 21180 6666 21232 6672
rect 20720 6656 20772 6662
rect 20720 6598 20772 6604
rect 20626 6216 20682 6225
rect 20626 6151 20682 6160
rect 20732 6118 20760 6598
rect 20720 6112 20772 6118
rect 20720 6054 20772 6060
rect 21088 5568 21140 5574
rect 21088 5510 21140 5516
rect 20904 5296 20956 5302
rect 20902 5264 20904 5273
rect 20956 5264 20958 5273
rect 20628 5228 20680 5234
rect 20902 5199 20958 5208
rect 20628 5170 20680 5176
rect 20640 5030 20668 5170
rect 20628 5024 20680 5030
rect 20628 4966 20680 4972
rect 20810 4584 20866 4593
rect 20810 4519 20866 4528
rect 20536 4480 20588 4486
rect 20536 4422 20588 4428
rect 20548 4214 20576 4422
rect 20536 4208 20588 4214
rect 20536 4150 20588 4156
rect 20718 3768 20774 3777
rect 20718 3703 20720 3712
rect 20772 3703 20774 3712
rect 20720 3674 20772 3680
rect 20628 2916 20680 2922
rect 20628 2858 20680 2864
rect 20640 2582 20668 2858
rect 20628 2576 20680 2582
rect 20628 2518 20680 2524
rect 20444 2304 20496 2310
rect 20444 2246 20496 2252
rect 20364 1686 20576 1714
rect 20548 800 20576 1686
rect 20824 800 20852 4519
rect 21100 4185 21128 5510
rect 21192 4690 21220 6666
rect 21376 6186 21404 12406
rect 21468 11393 21496 12582
rect 21454 11384 21510 11393
rect 21454 11319 21510 11328
rect 21560 8906 21588 15807
rect 21640 14408 21692 14414
rect 21640 14350 21692 14356
rect 21652 14006 21680 14350
rect 21640 14000 21692 14006
rect 21640 13942 21692 13948
rect 21744 11121 21772 29106
rect 21928 22094 21956 29582
rect 21836 22066 21956 22094
rect 21836 16402 21864 22066
rect 22112 22030 22140 32710
rect 22008 22024 22060 22030
rect 22008 21966 22060 21972
rect 22100 22024 22152 22030
rect 22100 21966 22152 21972
rect 22020 21690 22048 21966
rect 22100 21888 22152 21894
rect 22100 21830 22152 21836
rect 22008 21684 22060 21690
rect 22008 21626 22060 21632
rect 22112 20534 22140 21830
rect 22100 20528 22152 20534
rect 22100 20470 22152 20476
rect 22008 20392 22060 20398
rect 22008 20334 22060 20340
rect 22020 19378 22048 20334
rect 22204 19786 22232 32778
rect 22296 32502 22324 33594
rect 22388 33522 22416 34614
rect 22376 33516 22428 33522
rect 22376 33458 22428 33464
rect 22560 33516 22612 33522
rect 22560 33458 22612 33464
rect 22572 32858 22600 33458
rect 22664 33402 22692 60182
rect 22848 60110 22876 61202
rect 23216 60722 23244 63294
rect 23662 63294 23888 63322
rect 23662 63200 23718 63294
rect 23860 61198 23888 63294
rect 24398 63200 24454 64000
rect 25134 63200 25190 64000
rect 25870 63322 25926 64000
rect 25870 63294 26188 63322
rect 25870 63200 25926 63294
rect 23848 61192 23900 61198
rect 23848 61134 23900 61140
rect 23480 60852 23532 60858
rect 23480 60794 23532 60800
rect 23756 60852 23808 60858
rect 23756 60794 23808 60800
rect 23296 60784 23348 60790
rect 23296 60726 23348 60732
rect 23204 60716 23256 60722
rect 23204 60658 23256 60664
rect 22928 60512 22980 60518
rect 22928 60454 22980 60460
rect 22836 60104 22888 60110
rect 22836 60046 22888 60052
rect 22742 59664 22798 59673
rect 22742 59599 22744 59608
rect 22796 59599 22798 59608
rect 22744 59570 22796 59576
rect 22836 54596 22888 54602
rect 22836 54538 22888 54544
rect 22848 53961 22876 54538
rect 22834 53952 22890 53961
rect 22834 53887 22890 53896
rect 22940 38962 22968 60454
rect 23308 59634 23336 60726
rect 23388 60512 23440 60518
rect 23388 60454 23440 60460
rect 23400 60246 23428 60454
rect 23388 60240 23440 60246
rect 23388 60182 23440 60188
rect 23492 60110 23520 60794
rect 23768 60110 23796 60794
rect 24412 60790 24440 63200
rect 25148 61198 25176 63200
rect 26160 62098 26188 63294
rect 26606 63200 26662 64000
rect 27342 63322 27398 64000
rect 27342 63294 27568 63322
rect 27342 63200 27398 63294
rect 26160 62070 26280 62098
rect 26252 61198 26280 62070
rect 26620 61198 26648 63200
rect 25136 61192 25188 61198
rect 25136 61134 25188 61140
rect 26240 61192 26292 61198
rect 26240 61134 26292 61140
rect 26608 61192 26660 61198
rect 26608 61134 26660 61140
rect 24768 61124 24820 61130
rect 24768 61066 24820 61072
rect 24400 60784 24452 60790
rect 24400 60726 24452 60732
rect 23480 60104 23532 60110
rect 23480 60046 23532 60052
rect 23756 60104 23808 60110
rect 23756 60046 23808 60052
rect 23940 60104 23992 60110
rect 23940 60046 23992 60052
rect 23572 60036 23624 60042
rect 23572 59978 23624 59984
rect 23388 59696 23440 59702
rect 23386 59664 23388 59673
rect 23440 59664 23442 59673
rect 23296 59628 23348 59634
rect 23386 59599 23442 59608
rect 23296 59570 23348 59576
rect 23480 59492 23532 59498
rect 23480 59434 23532 59440
rect 23492 53446 23520 59434
rect 23584 56438 23612 59978
rect 23664 59628 23716 59634
rect 23664 59570 23716 59576
rect 23676 59430 23704 59570
rect 23664 59424 23716 59430
rect 23664 59366 23716 59372
rect 23572 56432 23624 56438
rect 23572 56374 23624 56380
rect 23848 56160 23900 56166
rect 23848 56102 23900 56108
rect 23480 53440 23532 53446
rect 23480 53382 23532 53388
rect 23480 45484 23532 45490
rect 23480 45426 23532 45432
rect 23296 40384 23348 40390
rect 23296 40326 23348 40332
rect 23308 39030 23336 40326
rect 23492 40186 23520 45426
rect 23480 40180 23532 40186
rect 23480 40122 23532 40128
rect 23756 40044 23808 40050
rect 23756 39986 23808 39992
rect 23572 39364 23624 39370
rect 23572 39306 23624 39312
rect 23296 39024 23348 39030
rect 23296 38966 23348 38972
rect 22928 38956 22980 38962
rect 22928 38898 22980 38904
rect 23204 38956 23256 38962
rect 23204 38898 23256 38904
rect 23112 38820 23164 38826
rect 23112 38762 23164 38768
rect 23020 38548 23072 38554
rect 23020 38490 23072 38496
rect 22928 38344 22980 38350
rect 22928 38286 22980 38292
rect 22940 37942 22968 38286
rect 23032 38214 23060 38490
rect 23020 38208 23072 38214
rect 23020 38150 23072 38156
rect 23032 38010 23060 38150
rect 23020 38004 23072 38010
rect 23020 37946 23072 37952
rect 22928 37936 22980 37942
rect 22926 37904 22928 37913
rect 22980 37904 22982 37913
rect 22926 37839 22982 37848
rect 23020 37868 23072 37874
rect 23020 37810 23072 37816
rect 23032 37777 23060 37810
rect 23018 37768 23074 37777
rect 23018 37703 23074 37712
rect 23124 37398 23152 38762
rect 23112 37392 23164 37398
rect 23112 37334 23164 37340
rect 22744 36032 22796 36038
rect 22744 35974 22796 35980
rect 22756 35290 22784 35974
rect 22744 35284 22796 35290
rect 22744 35226 22796 35232
rect 23020 34944 23072 34950
rect 23020 34886 23072 34892
rect 22836 34604 22888 34610
rect 22836 34546 22888 34552
rect 22742 34096 22798 34105
rect 22742 34031 22798 34040
rect 22756 33862 22784 34031
rect 22744 33856 22796 33862
rect 22744 33798 22796 33804
rect 22848 33522 22876 34546
rect 23032 33998 23060 34886
rect 23020 33992 23072 33998
rect 23020 33934 23072 33940
rect 22836 33516 22888 33522
rect 22836 33458 22888 33464
rect 22664 33374 22876 33402
rect 22652 33312 22704 33318
rect 22652 33254 22704 33260
rect 22664 33046 22692 33254
rect 22652 33040 22704 33046
rect 22652 32982 22704 32988
rect 22572 32830 22692 32858
rect 22284 32496 22336 32502
rect 22284 32438 22336 32444
rect 22284 30660 22336 30666
rect 22284 30602 22336 30608
rect 22296 30258 22324 30602
rect 22284 30252 22336 30258
rect 22284 30194 22336 30200
rect 22560 30252 22612 30258
rect 22560 30194 22612 30200
rect 22468 30184 22520 30190
rect 22468 30126 22520 30132
rect 22480 21690 22508 30126
rect 22572 29850 22600 30194
rect 22560 29844 22612 29850
rect 22560 29786 22612 29792
rect 22664 28558 22692 32830
rect 22744 32224 22796 32230
rect 22744 32166 22796 32172
rect 22756 31822 22784 32166
rect 22744 31816 22796 31822
rect 22744 31758 22796 31764
rect 22744 31272 22796 31278
rect 22744 31214 22796 31220
rect 22756 29578 22784 31214
rect 22744 29572 22796 29578
rect 22744 29514 22796 29520
rect 22652 28552 22704 28558
rect 22652 28494 22704 28500
rect 22848 28150 22876 33374
rect 22928 31952 22980 31958
rect 22928 31894 22980 31900
rect 22836 28144 22888 28150
rect 22836 28086 22888 28092
rect 22836 27328 22888 27334
rect 22836 27270 22888 27276
rect 22848 26994 22876 27270
rect 22836 26988 22888 26994
rect 22836 26930 22888 26936
rect 22558 25528 22614 25537
rect 22558 25463 22560 25472
rect 22612 25463 22614 25472
rect 22560 25434 22612 25440
rect 22560 22976 22612 22982
rect 22560 22918 22612 22924
rect 22284 21684 22336 21690
rect 22284 21626 22336 21632
rect 22468 21684 22520 21690
rect 22468 21626 22520 21632
rect 22296 21418 22324 21626
rect 22572 21434 22600 22918
rect 22940 22094 22968 31894
rect 23124 31754 23152 37334
rect 23216 36310 23244 38898
rect 23480 36576 23532 36582
rect 23480 36518 23532 36524
rect 23492 36378 23520 36518
rect 23480 36372 23532 36378
rect 23480 36314 23532 36320
rect 23204 36304 23256 36310
rect 23204 36246 23256 36252
rect 23296 36168 23348 36174
rect 23296 36110 23348 36116
rect 23388 36168 23440 36174
rect 23388 36110 23440 36116
rect 23308 35222 23336 36110
rect 23400 35630 23428 36110
rect 23584 36106 23612 39306
rect 23572 36100 23624 36106
rect 23572 36042 23624 36048
rect 23388 35624 23440 35630
rect 23388 35566 23440 35572
rect 23296 35216 23348 35222
rect 23296 35158 23348 35164
rect 23204 35012 23256 35018
rect 23204 34954 23256 34960
rect 23216 34474 23244 34954
rect 23204 34468 23256 34474
rect 23204 34410 23256 34416
rect 23572 34468 23624 34474
rect 23572 34410 23624 34416
rect 23296 33380 23348 33386
rect 23296 33322 23348 33328
rect 23204 32904 23256 32910
rect 23204 32846 23256 32852
rect 23032 31726 23152 31754
rect 23032 29646 23060 31726
rect 23216 30734 23244 32846
rect 23308 31958 23336 33322
rect 23296 31952 23348 31958
rect 23296 31894 23348 31900
rect 23296 31680 23348 31686
rect 23296 31622 23348 31628
rect 23308 30938 23336 31622
rect 23296 30932 23348 30938
rect 23296 30874 23348 30880
rect 23584 30734 23612 34410
rect 23768 31754 23796 39986
rect 23860 37618 23888 56102
rect 23952 53106 23980 60046
rect 24400 59968 24452 59974
rect 24400 59910 24452 59916
rect 24216 56432 24268 56438
rect 24216 56374 24268 56380
rect 24032 56296 24084 56302
rect 24032 56238 24084 56244
rect 23940 53100 23992 53106
rect 23940 53042 23992 53048
rect 23940 52896 23992 52902
rect 23940 52838 23992 52844
rect 23952 37806 23980 52838
rect 23940 37800 23992 37806
rect 23940 37742 23992 37748
rect 23860 37590 23980 37618
rect 23848 36712 23900 36718
rect 23848 36654 23900 36660
rect 23860 36378 23888 36654
rect 23848 36372 23900 36378
rect 23848 36314 23900 36320
rect 23676 31726 23796 31754
rect 23112 30728 23164 30734
rect 23112 30670 23164 30676
rect 23204 30728 23256 30734
rect 23204 30670 23256 30676
rect 23572 30728 23624 30734
rect 23572 30670 23624 30676
rect 23124 29850 23152 30670
rect 23112 29844 23164 29850
rect 23112 29786 23164 29792
rect 23020 29640 23072 29646
rect 23020 29582 23072 29588
rect 23032 29170 23060 29582
rect 23020 29164 23072 29170
rect 23020 29106 23072 29112
rect 23112 28076 23164 28082
rect 23112 28018 23164 28024
rect 23020 27872 23072 27878
rect 23020 27814 23072 27820
rect 23032 27470 23060 27814
rect 23020 27464 23072 27470
rect 23020 27406 23072 27412
rect 23124 25770 23152 28018
rect 23216 26994 23244 30670
rect 23388 29572 23440 29578
rect 23388 29514 23440 29520
rect 23296 28552 23348 28558
rect 23296 28494 23348 28500
rect 23308 28014 23336 28494
rect 23296 28008 23348 28014
rect 23296 27950 23348 27956
rect 23296 27464 23348 27470
rect 23296 27406 23348 27412
rect 23204 26988 23256 26994
rect 23204 26930 23256 26936
rect 23112 25764 23164 25770
rect 23112 25706 23164 25712
rect 23308 25702 23336 27406
rect 23400 27402 23428 29514
rect 23584 28150 23612 30670
rect 23572 28144 23624 28150
rect 23572 28086 23624 28092
rect 23388 27396 23440 27402
rect 23388 27338 23440 27344
rect 23296 25696 23348 25702
rect 23296 25638 23348 25644
rect 23400 23186 23428 27338
rect 23388 23180 23440 23186
rect 23388 23122 23440 23128
rect 23584 22094 23612 28086
rect 23676 27674 23704 31726
rect 23664 27668 23716 27674
rect 23664 27610 23716 27616
rect 22388 21418 22600 21434
rect 22284 21412 22336 21418
rect 22284 21354 22336 21360
rect 22376 21412 22600 21418
rect 22428 21406 22600 21412
rect 22664 22066 22968 22094
rect 23492 22066 23612 22094
rect 22376 21354 22428 21360
rect 22296 19854 22324 21354
rect 22284 19848 22336 19854
rect 22284 19790 22336 19796
rect 22192 19780 22244 19786
rect 22192 19722 22244 19728
rect 22008 19372 22060 19378
rect 22008 19314 22060 19320
rect 22020 18698 22048 19314
rect 22100 18964 22152 18970
rect 22100 18906 22152 18912
rect 22008 18692 22060 18698
rect 22008 18634 22060 18640
rect 21836 16374 21956 16402
rect 21824 16244 21876 16250
rect 21824 16186 21876 16192
rect 21836 16046 21864 16186
rect 21824 16040 21876 16046
rect 21824 15982 21876 15988
rect 21928 15881 21956 16374
rect 22020 16046 22048 18634
rect 22112 18426 22140 18906
rect 22192 18692 22244 18698
rect 22192 18634 22244 18640
rect 22100 18420 22152 18426
rect 22100 18362 22152 18368
rect 22204 18358 22232 18634
rect 22284 18624 22336 18630
rect 22284 18566 22336 18572
rect 22192 18352 22244 18358
rect 22192 18294 22244 18300
rect 22296 18290 22324 18566
rect 22388 18358 22416 21354
rect 22558 21312 22614 21321
rect 22664 21298 22692 22066
rect 22836 22024 22888 22030
rect 22836 21966 22888 21972
rect 22744 21684 22796 21690
rect 22744 21626 22796 21632
rect 22614 21270 22692 21298
rect 22558 21247 22614 21256
rect 22466 18456 22522 18465
rect 22466 18391 22522 18400
rect 22376 18352 22428 18358
rect 22376 18294 22428 18300
rect 22284 18284 22336 18290
rect 22284 18226 22336 18232
rect 22480 16658 22508 18391
rect 22468 16652 22520 16658
rect 22468 16594 22520 16600
rect 22192 16584 22244 16590
rect 22192 16526 22244 16532
rect 22008 16040 22060 16046
rect 22008 15982 22060 15988
rect 21914 15872 21970 15881
rect 21914 15807 21970 15816
rect 22020 15162 22048 15982
rect 22008 15156 22060 15162
rect 22008 15098 22060 15104
rect 22020 14482 22048 15098
rect 21824 14476 21876 14482
rect 21824 14418 21876 14424
rect 22008 14476 22060 14482
rect 22008 14418 22060 14424
rect 21836 13938 21864 14418
rect 21824 13932 21876 13938
rect 21824 13874 21876 13880
rect 22204 13841 22232 16526
rect 22284 16448 22336 16454
rect 22284 16390 22336 16396
rect 22190 13832 22246 13841
rect 21824 13796 21876 13802
rect 22190 13767 22246 13776
rect 21824 13738 21876 13744
rect 21836 12481 21864 13738
rect 22192 13728 22244 13734
rect 22192 13670 22244 13676
rect 22008 13184 22060 13190
rect 22008 13126 22060 13132
rect 21822 12472 21878 12481
rect 21822 12407 21878 12416
rect 21730 11112 21786 11121
rect 21730 11047 21786 11056
rect 21916 10532 21968 10538
rect 21916 10474 21968 10480
rect 21640 10192 21692 10198
rect 21928 10169 21956 10474
rect 21914 10160 21970 10169
rect 21640 10134 21692 10140
rect 21652 9994 21680 10134
rect 21744 10130 21864 10146
rect 21744 10124 21876 10130
rect 21744 10118 21824 10124
rect 21640 9988 21692 9994
rect 21640 9930 21692 9936
rect 21744 9586 21772 10118
rect 21914 10095 21970 10104
rect 21824 10066 21876 10072
rect 21824 9988 21876 9994
rect 21824 9930 21876 9936
rect 21732 9580 21784 9586
rect 21732 9522 21784 9528
rect 21548 8900 21600 8906
rect 21548 8842 21600 8848
rect 21456 7744 21508 7750
rect 21456 7686 21508 7692
rect 21468 7546 21496 7686
rect 21456 7540 21508 7546
rect 21456 7482 21508 7488
rect 21546 7304 21602 7313
rect 21546 7239 21602 7248
rect 21560 7206 21588 7239
rect 21456 7200 21508 7206
rect 21456 7142 21508 7148
rect 21548 7200 21600 7206
rect 21548 7142 21600 7148
rect 21468 6662 21496 7142
rect 21744 6866 21772 9522
rect 21732 6860 21784 6866
rect 21732 6802 21784 6808
rect 21456 6656 21508 6662
rect 21456 6598 21508 6604
rect 21364 6180 21416 6186
rect 21364 6122 21416 6128
rect 21376 5166 21404 6122
rect 21456 6112 21508 6118
rect 21456 6054 21508 6060
rect 21468 5710 21496 6054
rect 21836 5760 21864 9930
rect 21744 5732 21864 5760
rect 21456 5704 21508 5710
rect 21456 5646 21508 5652
rect 21364 5160 21416 5166
rect 21468 5137 21496 5646
rect 21364 5102 21416 5108
rect 21454 5128 21510 5137
rect 21376 4706 21404 5102
rect 21454 5063 21510 5072
rect 21180 4684 21232 4690
rect 21376 4678 21496 4706
rect 21180 4626 21232 4632
rect 21086 4176 21142 4185
rect 20996 4140 21048 4146
rect 21086 4111 21142 4120
rect 20996 4082 21048 4088
rect 21008 3670 21036 4082
rect 21192 4049 21220 4626
rect 21364 4616 21416 4622
rect 21364 4558 21416 4564
rect 21178 4040 21234 4049
rect 21178 3975 21234 3984
rect 20996 3664 21048 3670
rect 20902 3632 20958 3641
rect 20996 3606 21048 3612
rect 21192 3602 21220 3975
rect 21376 3942 21404 4558
rect 21468 4486 21496 4678
rect 21456 4480 21508 4486
rect 21456 4422 21508 4428
rect 21364 3936 21416 3942
rect 21364 3878 21416 3884
rect 20902 3567 20958 3576
rect 21180 3596 21232 3602
rect 20916 3466 20944 3567
rect 21180 3538 21232 3544
rect 20904 3460 20956 3466
rect 20904 3402 20956 3408
rect 20916 2854 20944 3402
rect 21088 3392 21140 3398
rect 21088 3334 21140 3340
rect 21456 3392 21508 3398
rect 21456 3334 21508 3340
rect 20904 2848 20956 2854
rect 20904 2790 20956 2796
rect 20996 2440 21048 2446
rect 20994 2408 20996 2417
rect 21048 2408 21050 2417
rect 20994 2343 21050 2352
rect 21100 800 21128 3334
rect 21468 3126 21496 3334
rect 21456 3120 21508 3126
rect 21456 3062 21508 3068
rect 21744 2961 21772 5732
rect 21822 5672 21878 5681
rect 21822 5607 21878 5616
rect 21836 3466 21864 5607
rect 22020 4622 22048 13126
rect 22204 11665 22232 13670
rect 22296 11694 22324 16390
rect 22466 16008 22522 16017
rect 22466 15943 22522 15952
rect 22376 13932 22428 13938
rect 22376 13874 22428 13880
rect 22388 11898 22416 13874
rect 22480 12434 22508 15943
rect 22572 12850 22600 21247
rect 22756 21026 22784 21626
rect 22664 20998 22784 21026
rect 22664 17898 22692 20998
rect 22744 20936 22796 20942
rect 22744 20878 22796 20884
rect 22756 20058 22784 20878
rect 22744 20052 22796 20058
rect 22744 19994 22796 20000
rect 22664 17870 22784 17898
rect 22652 17740 22704 17746
rect 22652 17682 22704 17688
rect 22664 17338 22692 17682
rect 22652 17332 22704 17338
rect 22652 17274 22704 17280
rect 22756 16402 22784 17870
rect 22848 16590 22876 21966
rect 23492 21554 23520 22066
rect 23480 21548 23532 21554
rect 23480 21490 23532 21496
rect 23020 21412 23072 21418
rect 23020 21354 23072 21360
rect 23032 20942 23060 21354
rect 23020 20936 23072 20942
rect 23020 20878 23072 20884
rect 22836 16584 22888 16590
rect 22836 16526 22888 16532
rect 22664 16374 22784 16402
rect 22664 15366 22692 16374
rect 22836 16176 22888 16182
rect 22836 16118 22888 16124
rect 22652 15360 22704 15366
rect 22652 15302 22704 15308
rect 22560 12844 22612 12850
rect 22560 12786 22612 12792
rect 22480 12406 22600 12434
rect 22376 11892 22428 11898
rect 22376 11834 22428 11840
rect 22284 11688 22336 11694
rect 22190 11656 22246 11665
rect 22284 11630 22336 11636
rect 22190 11591 22246 11600
rect 22100 10464 22152 10470
rect 22100 10406 22152 10412
rect 22112 10169 22140 10406
rect 22098 10160 22154 10169
rect 22098 10095 22154 10104
rect 22284 10124 22336 10130
rect 22284 10066 22336 10072
rect 22296 8430 22324 10066
rect 22468 8968 22520 8974
rect 22466 8936 22468 8945
rect 22520 8936 22522 8945
rect 22466 8871 22522 8880
rect 22376 8492 22428 8498
rect 22376 8434 22428 8440
rect 22284 8424 22336 8430
rect 22284 8366 22336 8372
rect 22284 7744 22336 7750
rect 22284 7686 22336 7692
rect 22296 6730 22324 7686
rect 22388 7177 22416 8434
rect 22374 7168 22430 7177
rect 22374 7103 22430 7112
rect 22284 6724 22336 6730
rect 22284 6666 22336 6672
rect 22374 5536 22430 5545
rect 22374 5471 22430 5480
rect 22388 4622 22416 5471
rect 22468 5160 22520 5166
rect 22468 5102 22520 5108
rect 22008 4616 22060 4622
rect 22008 4558 22060 4564
rect 22376 4616 22428 4622
rect 22376 4558 22428 4564
rect 22376 4276 22428 4282
rect 22376 4218 22428 4224
rect 22388 4146 22416 4218
rect 22376 4140 22428 4146
rect 22376 4082 22428 4088
rect 22376 3596 22428 3602
rect 22376 3538 22428 3544
rect 21824 3460 21876 3466
rect 21824 3402 21876 3408
rect 22282 3224 22338 3233
rect 22282 3159 22338 3168
rect 22296 3058 22324 3159
rect 22388 3058 22416 3538
rect 21916 3052 21968 3058
rect 21916 2994 21968 3000
rect 22284 3052 22336 3058
rect 22284 2994 22336 3000
rect 22376 3052 22428 3058
rect 22376 2994 22428 3000
rect 21730 2952 21786 2961
rect 21730 2887 21786 2896
rect 21364 2644 21416 2650
rect 21364 2586 21416 2592
rect 21376 800 21404 2586
rect 21640 2304 21692 2310
rect 21640 2246 21692 2252
rect 21652 800 21680 2246
rect 21928 800 21956 2994
rect 22192 2916 22244 2922
rect 22192 2858 22244 2864
rect 22008 2848 22060 2854
rect 22008 2790 22060 2796
rect 22020 2514 22048 2790
rect 22008 2508 22060 2514
rect 22008 2450 22060 2456
rect 22204 800 22232 2858
rect 22480 800 22508 5102
rect 22572 2774 22600 12406
rect 22744 11892 22796 11898
rect 22744 11834 22796 11840
rect 22756 11082 22784 11834
rect 22744 11076 22796 11082
rect 22744 11018 22796 11024
rect 22650 8936 22706 8945
rect 22650 8871 22706 8880
rect 22664 6322 22692 8871
rect 22742 8800 22798 8809
rect 22742 8735 22798 8744
rect 22756 8634 22784 8735
rect 22744 8628 22796 8634
rect 22744 8570 22796 8576
rect 22652 6316 22704 6322
rect 22652 6258 22704 6264
rect 22744 4548 22796 4554
rect 22744 4490 22796 4496
rect 22572 2746 22692 2774
rect 22664 2446 22692 2746
rect 22652 2440 22704 2446
rect 22652 2382 22704 2388
rect 22756 800 22784 4490
rect 22848 2038 22876 16118
rect 22928 14272 22980 14278
rect 22928 14214 22980 14220
rect 22940 6662 22968 14214
rect 23032 14006 23060 20878
rect 23492 20806 23520 21490
rect 23480 20800 23532 20806
rect 23480 20742 23532 20748
rect 23204 20256 23256 20262
rect 23204 20198 23256 20204
rect 23216 19854 23244 20198
rect 23204 19848 23256 19854
rect 23204 19790 23256 19796
rect 23112 19780 23164 19786
rect 23112 19722 23164 19728
rect 23020 14000 23072 14006
rect 23020 13942 23072 13948
rect 23020 13864 23072 13870
rect 23020 13806 23072 13812
rect 23032 12986 23060 13806
rect 23020 12980 23072 12986
rect 23020 12922 23072 12928
rect 23020 12844 23072 12850
rect 23020 12786 23072 12792
rect 23032 12374 23060 12786
rect 23020 12368 23072 12374
rect 23020 12310 23072 12316
rect 23020 12096 23072 12102
rect 23020 12038 23072 12044
rect 23032 11762 23060 12038
rect 23020 11756 23072 11762
rect 23020 11698 23072 11704
rect 23018 11656 23074 11665
rect 23018 11591 23074 11600
rect 23032 11150 23060 11591
rect 23124 11150 23152 19722
rect 23216 17746 23244 19790
rect 23480 19236 23532 19242
rect 23480 19178 23532 19184
rect 23388 19168 23440 19174
rect 23308 19116 23388 19122
rect 23308 19110 23440 19116
rect 23308 19094 23428 19110
rect 23308 18222 23336 19094
rect 23492 18766 23520 19178
rect 23480 18760 23532 18766
rect 23480 18702 23532 18708
rect 23388 18624 23440 18630
rect 23388 18566 23440 18572
rect 23400 18329 23428 18566
rect 23572 18420 23624 18426
rect 23572 18362 23624 18368
rect 23386 18320 23442 18329
rect 23584 18290 23612 18362
rect 23386 18255 23442 18264
rect 23572 18284 23624 18290
rect 23572 18226 23624 18232
rect 23296 18216 23348 18222
rect 23296 18158 23348 18164
rect 23480 18216 23532 18222
rect 23480 18158 23532 18164
rect 23388 18148 23440 18154
rect 23388 18090 23440 18096
rect 23400 17882 23428 18090
rect 23388 17876 23440 17882
rect 23388 17818 23440 17824
rect 23204 17740 23256 17746
rect 23204 17682 23256 17688
rect 23492 17678 23520 18158
rect 23584 18086 23612 18226
rect 23572 18080 23624 18086
rect 23572 18022 23624 18028
rect 23480 17672 23532 17678
rect 23480 17614 23532 17620
rect 23388 16652 23440 16658
rect 23388 16594 23440 16600
rect 23204 16584 23256 16590
rect 23204 16526 23256 16532
rect 23216 15552 23244 16526
rect 23400 16454 23428 16594
rect 23388 16448 23440 16454
rect 23388 16390 23440 16396
rect 23400 16114 23428 16390
rect 23388 16108 23440 16114
rect 23388 16050 23440 16056
rect 23492 15978 23520 17614
rect 23676 17610 23704 27610
rect 23848 21888 23900 21894
rect 23848 21830 23900 21836
rect 23860 20942 23888 21830
rect 23848 20936 23900 20942
rect 23848 20878 23900 20884
rect 23756 19712 23808 19718
rect 23756 19654 23808 19660
rect 23768 19242 23796 19654
rect 23756 19236 23808 19242
rect 23756 19178 23808 19184
rect 23664 17604 23716 17610
rect 23716 17564 23796 17592
rect 23664 17546 23716 17552
rect 23664 16992 23716 16998
rect 23664 16934 23716 16940
rect 23572 16652 23624 16658
rect 23572 16594 23624 16600
rect 23584 16182 23612 16594
rect 23572 16176 23624 16182
rect 23572 16118 23624 16124
rect 23480 15972 23532 15978
rect 23480 15914 23532 15920
rect 23572 15904 23624 15910
rect 23572 15846 23624 15852
rect 23480 15632 23532 15638
rect 23480 15574 23532 15580
rect 23216 15524 23336 15552
rect 23204 15428 23256 15434
rect 23204 15370 23256 15376
rect 23216 13802 23244 15370
rect 23308 14090 23336 15524
rect 23386 15464 23442 15473
rect 23386 15399 23442 15408
rect 23400 15366 23428 15399
rect 23492 15366 23520 15574
rect 23584 15570 23612 15846
rect 23572 15564 23624 15570
rect 23572 15506 23624 15512
rect 23388 15360 23440 15366
rect 23388 15302 23440 15308
rect 23480 15360 23532 15366
rect 23480 15302 23532 15308
rect 23308 14062 23428 14090
rect 23204 13796 23256 13802
rect 23204 13738 23256 13744
rect 23216 12238 23244 13738
rect 23400 13258 23428 14062
rect 23572 13932 23624 13938
rect 23572 13874 23624 13880
rect 23480 13388 23532 13394
rect 23480 13330 23532 13336
rect 23388 13252 23440 13258
rect 23388 13194 23440 13200
rect 23492 12986 23520 13330
rect 23480 12980 23532 12986
rect 23480 12922 23532 12928
rect 23480 12436 23532 12442
rect 23480 12378 23532 12384
rect 23388 12368 23440 12374
rect 23388 12310 23440 12316
rect 23296 12300 23348 12306
rect 23296 12242 23348 12248
rect 23204 12232 23256 12238
rect 23204 12174 23256 12180
rect 23308 12102 23336 12242
rect 23296 12096 23348 12102
rect 23296 12038 23348 12044
rect 23294 11928 23350 11937
rect 23294 11863 23350 11872
rect 23020 11144 23072 11150
rect 23020 11086 23072 11092
rect 23112 11144 23164 11150
rect 23112 11086 23164 11092
rect 23032 10169 23060 11086
rect 23124 10441 23152 11086
rect 23110 10432 23166 10441
rect 23110 10367 23166 10376
rect 23308 10282 23336 11863
rect 23400 10742 23428 12310
rect 23492 11898 23520 12378
rect 23480 11892 23532 11898
rect 23480 11834 23532 11840
rect 23388 10736 23440 10742
rect 23388 10678 23440 10684
rect 23216 10254 23336 10282
rect 23018 10160 23074 10169
rect 23018 10095 23074 10104
rect 23020 9716 23072 9722
rect 23020 9658 23072 9664
rect 23032 9466 23060 9658
rect 23032 9438 23152 9466
rect 23020 9376 23072 9382
rect 23020 9318 23072 9324
rect 23032 8838 23060 9318
rect 23020 8832 23072 8838
rect 23020 8774 23072 8780
rect 23032 8294 23060 8774
rect 23124 8514 23152 9438
rect 23216 8616 23244 10254
rect 23400 9897 23428 10678
rect 23480 10600 23532 10606
rect 23480 10542 23532 10548
rect 23492 10198 23520 10542
rect 23480 10192 23532 10198
rect 23480 10134 23532 10140
rect 23386 9888 23442 9897
rect 23386 9823 23442 9832
rect 23386 9752 23442 9761
rect 23386 9687 23442 9696
rect 23400 9353 23428 9687
rect 23584 9654 23612 13874
rect 23676 10985 23704 16934
rect 23768 12238 23796 17564
rect 23848 16584 23900 16590
rect 23848 16526 23900 16532
rect 23860 14346 23888 16526
rect 23848 14340 23900 14346
rect 23848 14282 23900 14288
rect 23952 14006 23980 37590
rect 24044 36786 24072 56238
rect 24124 51604 24176 51610
rect 24124 51546 24176 51552
rect 24136 37806 24164 51546
rect 24228 45490 24256 56374
rect 24412 56370 24440 59910
rect 24492 59424 24544 59430
rect 24492 59366 24544 59372
rect 24400 56364 24452 56370
rect 24400 56306 24452 56312
rect 24308 55684 24360 55690
rect 24308 55626 24360 55632
rect 24216 45484 24268 45490
rect 24216 45426 24268 45432
rect 24124 37800 24176 37806
rect 24124 37742 24176 37748
rect 24032 36780 24084 36786
rect 24032 36722 24084 36728
rect 24136 35698 24164 37742
rect 24124 35692 24176 35698
rect 24124 35634 24176 35640
rect 24032 33924 24084 33930
rect 24032 33866 24084 33872
rect 24044 16402 24072 33866
rect 24136 31346 24164 35634
rect 24124 31340 24176 31346
rect 24124 31282 24176 31288
rect 24216 31340 24268 31346
rect 24216 31282 24268 31288
rect 24136 30122 24164 31282
rect 24228 30938 24256 31282
rect 24216 30932 24268 30938
rect 24216 30874 24268 30880
rect 24124 30116 24176 30122
rect 24124 30058 24176 30064
rect 24136 16998 24164 30058
rect 24320 20618 24348 55626
rect 24400 37664 24452 37670
rect 24400 37606 24452 37612
rect 24412 31754 24440 37606
rect 24504 33998 24532 59366
rect 24780 56370 24808 61066
rect 25412 61056 25464 61062
rect 25412 60998 25464 61004
rect 27344 61056 27396 61062
rect 27344 60998 27396 61004
rect 25228 60512 25280 60518
rect 25228 60454 25280 60460
rect 24768 56364 24820 56370
rect 24768 56306 24820 56312
rect 24860 54800 24912 54806
rect 24860 54742 24912 54748
rect 24584 53440 24636 53446
rect 24584 53382 24636 53388
rect 24596 53106 24624 53382
rect 24584 53100 24636 53106
rect 24584 53042 24636 53048
rect 24596 51074 24624 53042
rect 24596 51046 24716 51074
rect 24584 36576 24636 36582
rect 24584 36518 24636 36524
rect 24596 36174 24624 36518
rect 24584 36168 24636 36174
rect 24584 36110 24636 36116
rect 24688 35766 24716 51046
rect 24768 38752 24820 38758
rect 24768 38694 24820 38700
rect 24780 36174 24808 38694
rect 24768 36168 24820 36174
rect 24768 36110 24820 36116
rect 24676 35760 24728 35766
rect 24676 35702 24728 35708
rect 24872 35086 24900 54742
rect 24952 53508 25004 53514
rect 24952 53450 25004 53456
rect 24964 53242 24992 53450
rect 24952 53236 25004 53242
rect 24952 53178 25004 53184
rect 24964 52698 24992 53178
rect 24952 52692 25004 52698
rect 24952 52634 25004 52640
rect 25240 37942 25268 60454
rect 25320 56364 25372 56370
rect 25320 56306 25372 56312
rect 25332 55758 25360 56306
rect 25320 55752 25372 55758
rect 25320 55694 25372 55700
rect 25332 54806 25360 55694
rect 25320 54800 25372 54806
rect 25320 54742 25372 54748
rect 25424 47666 25452 60998
rect 26884 60172 26936 60178
rect 26884 60114 26936 60120
rect 26896 56914 26924 60114
rect 26884 56908 26936 56914
rect 26884 56850 26936 56856
rect 25688 55752 25740 55758
rect 25688 55694 25740 55700
rect 25700 54670 25728 55694
rect 25688 54664 25740 54670
rect 25688 54606 25740 54612
rect 27356 48929 27384 60998
rect 27540 60790 27568 63294
rect 28078 63200 28134 64000
rect 28814 63200 28870 64000
rect 29550 63322 29606 64000
rect 29550 63294 29868 63322
rect 29550 63200 29606 63294
rect 28092 61198 28120 63200
rect 28448 61668 28500 61674
rect 28448 61610 28500 61616
rect 28080 61192 28132 61198
rect 28080 61134 28132 61140
rect 28172 61124 28224 61130
rect 28172 61066 28224 61072
rect 27528 60784 27580 60790
rect 27528 60726 27580 60732
rect 28184 60110 28212 61066
rect 28356 61056 28408 61062
rect 28356 60998 28408 61004
rect 28080 60104 28132 60110
rect 28080 60046 28132 60052
rect 28172 60104 28224 60110
rect 28172 60046 28224 60052
rect 28092 54534 28120 60046
rect 28080 54528 28132 54534
rect 28080 54470 28132 54476
rect 27342 48920 27398 48929
rect 27342 48855 27398 48864
rect 25412 47660 25464 47666
rect 25412 47602 25464 47608
rect 26240 47592 26292 47598
rect 26240 47534 26292 47540
rect 25320 40180 25372 40186
rect 25320 40122 25372 40128
rect 25228 37936 25280 37942
rect 25228 37878 25280 37884
rect 25332 37874 25360 40122
rect 26148 38208 26200 38214
rect 26148 38150 26200 38156
rect 26160 38010 26188 38150
rect 26148 38004 26200 38010
rect 26148 37946 26200 37952
rect 25320 37868 25372 37874
rect 25320 37810 25372 37816
rect 24952 36032 25004 36038
rect 24952 35974 25004 35980
rect 24860 35080 24912 35086
rect 24860 35022 24912 35028
rect 24872 34649 24900 35022
rect 24858 34640 24914 34649
rect 24858 34575 24914 34584
rect 24492 33992 24544 33998
rect 24964 33946 24992 35974
rect 25332 33998 25360 37810
rect 25504 36780 25556 36786
rect 25504 36722 25556 36728
rect 25412 36100 25464 36106
rect 25412 36042 25464 36048
rect 24492 33934 24544 33940
rect 24872 33930 24992 33946
rect 25320 33992 25372 33998
rect 25320 33934 25372 33940
rect 24860 33924 24992 33930
rect 24912 33918 24992 33924
rect 24860 33866 24912 33872
rect 24768 32904 24820 32910
rect 24768 32846 24820 32852
rect 24412 31726 24532 31754
rect 24320 20590 24440 20618
rect 24308 20460 24360 20466
rect 24308 20402 24360 20408
rect 24216 20256 24268 20262
rect 24216 20198 24268 20204
rect 24228 19378 24256 20198
rect 24320 20058 24348 20402
rect 24308 20052 24360 20058
rect 24308 19994 24360 20000
rect 24216 19372 24268 19378
rect 24216 19314 24268 19320
rect 24308 19372 24360 19378
rect 24308 19314 24360 19320
rect 24320 18426 24348 19314
rect 24308 18420 24360 18426
rect 24308 18362 24360 18368
rect 24412 17241 24440 20590
rect 24398 17232 24454 17241
rect 24398 17167 24454 17176
rect 24124 16992 24176 16998
rect 24124 16934 24176 16940
rect 24504 16590 24532 31726
rect 24584 31476 24636 31482
rect 24584 31418 24636 31424
rect 24596 31346 24624 31418
rect 24584 31340 24636 31346
rect 24584 31282 24636 31288
rect 24780 31210 24808 32846
rect 24768 31204 24820 31210
rect 24768 31146 24820 31152
rect 24860 30592 24912 30598
rect 24860 30534 24912 30540
rect 24872 29617 24900 30534
rect 24858 29608 24914 29617
rect 24858 29543 24914 29552
rect 24964 29510 24992 33918
rect 25228 33856 25280 33862
rect 25228 33798 25280 33804
rect 25240 33046 25268 33798
rect 25228 33040 25280 33046
rect 25228 32982 25280 32988
rect 24952 29504 25004 29510
rect 24952 29446 25004 29452
rect 24952 22772 25004 22778
rect 24952 22714 25004 22720
rect 24584 22636 24636 22642
rect 24584 22578 24636 22584
rect 24596 17882 24624 22578
rect 24676 22500 24728 22506
rect 24676 22442 24728 22448
rect 24584 17876 24636 17882
rect 24584 17818 24636 17824
rect 24584 17740 24636 17746
rect 24584 17682 24636 17688
rect 24596 17202 24624 17682
rect 24584 17196 24636 17202
rect 24584 17138 24636 17144
rect 24492 16584 24544 16590
rect 24492 16526 24544 16532
rect 24044 16374 24440 16402
rect 24124 16244 24176 16250
rect 24124 16186 24176 16192
rect 24032 15972 24084 15978
rect 24032 15914 24084 15920
rect 24044 14822 24072 15914
rect 24032 14816 24084 14822
rect 24032 14758 24084 14764
rect 23940 14000 23992 14006
rect 23940 13942 23992 13948
rect 23940 13524 23992 13530
rect 23940 13466 23992 13472
rect 23848 13320 23900 13326
rect 23848 13262 23900 13268
rect 23860 13161 23888 13262
rect 23846 13152 23902 13161
rect 23846 13087 23902 13096
rect 23756 12232 23808 12238
rect 23756 12174 23808 12180
rect 23756 11620 23808 11626
rect 23952 11608 23980 13466
rect 24044 13326 24072 14758
rect 24032 13320 24084 13326
rect 24032 13262 24084 13268
rect 24030 12064 24086 12073
rect 24030 11999 24086 12008
rect 23808 11580 23980 11608
rect 23756 11562 23808 11568
rect 23768 11150 23796 11562
rect 24044 11558 24072 11999
rect 24032 11552 24084 11558
rect 24032 11494 24084 11500
rect 23848 11280 23900 11286
rect 23848 11222 23900 11228
rect 23756 11144 23808 11150
rect 23756 11086 23808 11092
rect 23662 10976 23718 10985
rect 23662 10911 23718 10920
rect 23676 10470 23704 10911
rect 23664 10464 23716 10470
rect 23664 10406 23716 10412
rect 23664 10260 23716 10266
rect 23664 10202 23716 10208
rect 23676 9994 23704 10202
rect 23664 9988 23716 9994
rect 23664 9930 23716 9936
rect 23572 9648 23624 9654
rect 23572 9590 23624 9596
rect 23480 9512 23532 9518
rect 23480 9454 23532 9460
rect 23386 9344 23442 9353
rect 23386 9279 23442 9288
rect 23492 9330 23520 9454
rect 23570 9344 23626 9353
rect 23492 9302 23570 9330
rect 23388 8900 23440 8906
rect 23388 8842 23440 8848
rect 23296 8628 23348 8634
rect 23216 8588 23296 8616
rect 23296 8570 23348 8576
rect 23124 8486 23244 8514
rect 23020 8288 23072 8294
rect 23020 8230 23072 8236
rect 23032 7750 23060 8230
rect 23020 7744 23072 7750
rect 23020 7686 23072 7692
rect 23112 7744 23164 7750
rect 23112 7686 23164 7692
rect 22928 6656 22980 6662
rect 22928 6598 22980 6604
rect 23124 5914 23152 7686
rect 23112 5908 23164 5914
rect 23112 5850 23164 5856
rect 23216 5794 23244 8486
rect 23296 6724 23348 6730
rect 23296 6666 23348 6672
rect 23124 5778 23244 5794
rect 23112 5772 23244 5778
rect 23164 5766 23244 5772
rect 23112 5714 23164 5720
rect 23204 5704 23256 5710
rect 23204 5646 23256 5652
rect 23020 4072 23072 4078
rect 23020 4014 23072 4020
rect 22836 2032 22888 2038
rect 22836 1974 22888 1980
rect 23032 800 23060 4014
rect 23216 3942 23244 5646
rect 23308 5642 23336 6666
rect 23400 5914 23428 8842
rect 23492 7834 23520 9302
rect 23570 9279 23626 9288
rect 23664 9172 23716 9178
rect 23664 9114 23716 9120
rect 23572 9104 23624 9110
rect 23572 9046 23624 9052
rect 23584 8294 23612 9046
rect 23676 8974 23704 9114
rect 23664 8968 23716 8974
rect 23664 8910 23716 8916
rect 23572 8288 23624 8294
rect 23572 8230 23624 8236
rect 23768 7954 23796 11086
rect 23860 9353 23888 11222
rect 23938 11112 23994 11121
rect 23938 11047 23940 11056
rect 23992 11047 23994 11056
rect 23940 11018 23992 11024
rect 23940 9580 23992 9586
rect 23940 9522 23992 9528
rect 23952 9382 23980 9522
rect 23940 9376 23992 9382
rect 23846 9344 23902 9353
rect 23940 9318 23992 9324
rect 23846 9279 23902 9288
rect 23848 8832 23900 8838
rect 23848 8774 23900 8780
rect 23860 8634 23888 8774
rect 23848 8628 23900 8634
rect 23848 8570 23900 8576
rect 23952 8430 23980 9318
rect 24044 9110 24072 11494
rect 24032 9104 24084 9110
rect 24032 9046 24084 9052
rect 24136 8974 24164 16186
rect 24216 16176 24268 16182
rect 24216 16118 24268 16124
rect 24124 8968 24176 8974
rect 24124 8910 24176 8916
rect 24032 8900 24084 8906
rect 24032 8842 24084 8848
rect 23940 8424 23992 8430
rect 23940 8366 23992 8372
rect 23756 7948 23808 7954
rect 23756 7890 23808 7896
rect 23492 7806 23612 7834
rect 23480 7744 23532 7750
rect 23480 7686 23532 7692
rect 23492 7546 23520 7686
rect 23480 7540 23532 7546
rect 23480 7482 23532 7488
rect 23388 5908 23440 5914
rect 23388 5850 23440 5856
rect 23296 5636 23348 5642
rect 23296 5578 23348 5584
rect 23386 5400 23442 5409
rect 23386 5335 23442 5344
rect 23400 5234 23428 5335
rect 23388 5228 23440 5234
rect 23388 5170 23440 5176
rect 23584 5137 23612 7806
rect 23664 5636 23716 5642
rect 23664 5578 23716 5584
rect 23570 5128 23626 5137
rect 23570 5063 23626 5072
rect 23676 5001 23704 5578
rect 23662 4992 23718 5001
rect 23662 4927 23718 4936
rect 23768 4758 23796 7890
rect 24044 7886 24072 8842
rect 24122 8800 24178 8809
rect 24122 8735 24178 8744
rect 24136 8498 24164 8735
rect 24124 8492 24176 8498
rect 24124 8434 24176 8440
rect 24228 8242 24256 16118
rect 24412 15586 24440 16374
rect 24412 15558 24624 15586
rect 24492 15496 24544 15502
rect 24492 15438 24544 15444
rect 24308 15020 24360 15026
rect 24308 14962 24360 14968
rect 24320 14346 24348 14962
rect 24400 14544 24452 14550
rect 24400 14486 24452 14492
rect 24308 14340 24360 14346
rect 24308 14282 24360 14288
rect 24412 14074 24440 14486
rect 24400 14068 24452 14074
rect 24400 14010 24452 14016
rect 24400 13864 24452 13870
rect 24398 13832 24400 13841
rect 24452 13832 24454 13841
rect 24398 13767 24454 13776
rect 24308 12096 24360 12102
rect 24306 12064 24308 12073
rect 24360 12064 24362 12073
rect 24306 11999 24362 12008
rect 24504 11665 24532 15438
rect 24596 13410 24624 15558
rect 24688 15450 24716 22442
rect 24860 22432 24912 22438
rect 24860 22374 24912 22380
rect 24872 19446 24900 22374
rect 24964 21690 24992 22714
rect 25044 21956 25096 21962
rect 25044 21898 25096 21904
rect 25056 21690 25084 21898
rect 24952 21684 25004 21690
rect 24952 21626 25004 21632
rect 25044 21684 25096 21690
rect 25044 21626 25096 21632
rect 25044 21480 25096 21486
rect 25044 21422 25096 21428
rect 24952 19848 25004 19854
rect 24950 19816 24952 19825
rect 25004 19816 25006 19825
rect 24950 19751 25006 19760
rect 24952 19712 25004 19718
rect 24952 19654 25004 19660
rect 24860 19440 24912 19446
rect 24860 19382 24912 19388
rect 24768 18760 24820 18766
rect 24768 18702 24820 18708
rect 24780 18465 24808 18702
rect 24766 18456 24822 18465
rect 24766 18391 24822 18400
rect 24768 18284 24820 18290
rect 24768 18226 24820 18232
rect 24780 16726 24808 18226
rect 24964 17678 24992 19654
rect 25056 17746 25084 21422
rect 25228 20800 25280 20806
rect 25228 20742 25280 20748
rect 25134 20496 25190 20505
rect 25134 20431 25190 20440
rect 25044 17740 25096 17746
rect 25044 17682 25096 17688
rect 24952 17672 25004 17678
rect 24952 17614 25004 17620
rect 24860 17536 24912 17542
rect 25044 17536 25096 17542
rect 24860 17478 24912 17484
rect 25042 17504 25044 17513
rect 25096 17504 25098 17513
rect 24768 16720 24820 16726
rect 24768 16662 24820 16668
rect 24872 16590 24900 17478
rect 25042 17439 25098 17448
rect 25148 17202 25176 20431
rect 25240 19334 25268 20742
rect 25424 20482 25452 36042
rect 25516 20618 25544 36722
rect 26252 35894 26280 47534
rect 26884 41472 26936 41478
rect 26884 41414 26936 41420
rect 26252 35866 26372 35894
rect 25596 22568 25648 22574
rect 25596 22510 25648 22516
rect 25608 21418 25636 22510
rect 26148 22092 26200 22098
rect 26148 22034 26200 22040
rect 25872 21888 25924 21894
rect 25872 21830 25924 21836
rect 25884 21570 25912 21830
rect 25884 21542 26004 21570
rect 25596 21412 25648 21418
rect 25596 21354 25648 21360
rect 25976 20806 26004 21542
rect 26160 21486 26188 22034
rect 26148 21480 26200 21486
rect 26148 21422 26200 21428
rect 26240 20936 26292 20942
rect 26240 20878 26292 20884
rect 25964 20800 26016 20806
rect 25964 20742 26016 20748
rect 25516 20590 25728 20618
rect 25424 20454 25636 20482
rect 25320 20392 25372 20398
rect 25320 20334 25372 20340
rect 25504 20392 25556 20398
rect 25504 20334 25556 20340
rect 25332 19854 25360 20334
rect 25412 19984 25464 19990
rect 25412 19926 25464 19932
rect 25320 19848 25372 19854
rect 25320 19790 25372 19796
rect 25240 19306 25360 19334
rect 25424 19310 25452 19926
rect 25516 19922 25544 20334
rect 25504 19916 25556 19922
rect 25504 19858 25556 19864
rect 25608 19802 25636 20454
rect 25516 19774 25636 19802
rect 25228 17264 25280 17270
rect 25226 17232 25228 17241
rect 25280 17232 25282 17241
rect 25136 17196 25188 17202
rect 25226 17167 25282 17176
rect 25136 17138 25188 17144
rect 24860 16584 24912 16590
rect 25332 16538 25360 19306
rect 25412 19304 25464 19310
rect 25412 19246 25464 19252
rect 25412 17264 25464 17270
rect 25412 17206 25464 17212
rect 24860 16526 24912 16532
rect 24964 16510 25360 16538
rect 24860 16448 24912 16454
rect 24858 16416 24860 16425
rect 24912 16416 24914 16425
rect 24858 16351 24914 16360
rect 24860 16040 24912 16046
rect 24860 15982 24912 15988
rect 24872 15706 24900 15982
rect 24860 15700 24912 15706
rect 24860 15642 24912 15648
rect 24964 15586 24992 16510
rect 25424 16454 25452 17206
rect 25044 16448 25096 16454
rect 25412 16448 25464 16454
rect 25044 16390 25096 16396
rect 25226 16416 25282 16425
rect 24872 15558 24992 15586
rect 24688 15434 24808 15450
rect 24688 15428 24820 15434
rect 24688 15422 24768 15428
rect 24688 15201 24716 15422
rect 24768 15370 24820 15376
rect 24674 15192 24730 15201
rect 24674 15127 24730 15136
rect 24768 15020 24820 15026
rect 24768 14962 24820 14968
rect 24596 13382 24716 13410
rect 24688 13326 24716 13382
rect 24676 13320 24728 13326
rect 24676 13262 24728 13268
rect 24780 12850 24808 14962
rect 24872 14600 24900 15558
rect 24952 15496 25004 15502
rect 24952 15438 25004 15444
rect 24964 14822 24992 15438
rect 24952 14816 25004 14822
rect 24952 14758 25004 14764
rect 24872 14572 24992 14600
rect 24860 14476 24912 14482
rect 24860 14418 24912 14424
rect 24872 13870 24900 14418
rect 24964 13938 24992 14572
rect 24952 13932 25004 13938
rect 24952 13874 25004 13880
rect 24860 13864 24912 13870
rect 24860 13806 24912 13812
rect 24768 12844 24820 12850
rect 24768 12786 24820 12792
rect 24768 12368 24820 12374
rect 24768 12310 24820 12316
rect 24780 12238 24808 12310
rect 24872 12306 24900 13806
rect 25056 13394 25084 16390
rect 25412 16390 25464 16396
rect 25226 16351 25282 16360
rect 25136 15360 25188 15366
rect 25136 15302 25188 15308
rect 25044 13388 25096 13394
rect 25044 13330 25096 13336
rect 25148 13326 25176 15302
rect 24952 13320 25004 13326
rect 24952 13262 25004 13268
rect 25136 13320 25188 13326
rect 25136 13262 25188 13268
rect 24964 13190 24992 13262
rect 24952 13184 25004 13190
rect 24952 13126 25004 13132
rect 25136 12980 25188 12986
rect 25136 12922 25188 12928
rect 25044 12436 25096 12442
rect 25044 12378 25096 12384
rect 24860 12300 24912 12306
rect 24860 12242 24912 12248
rect 25056 12238 25084 12378
rect 24584 12232 24636 12238
rect 24584 12174 24636 12180
rect 24768 12232 24820 12238
rect 24768 12174 24820 12180
rect 25044 12232 25096 12238
rect 25044 12174 25096 12180
rect 24490 11656 24546 11665
rect 24490 11591 24546 11600
rect 24596 11286 24624 12174
rect 24860 12096 24912 12102
rect 24860 12038 24912 12044
rect 24676 11688 24728 11694
rect 24676 11630 24728 11636
rect 24308 11280 24360 11286
rect 24584 11280 24636 11286
rect 24308 11222 24360 11228
rect 24398 11248 24454 11257
rect 24320 10470 24348 11222
rect 24584 11222 24636 11228
rect 24398 11183 24454 11192
rect 24308 10464 24360 10470
rect 24308 10406 24360 10412
rect 24308 9512 24360 9518
rect 24308 9454 24360 9460
rect 24320 9353 24348 9454
rect 24306 9344 24362 9353
rect 24306 9279 24362 9288
rect 24320 8673 24348 9279
rect 24412 9217 24440 11183
rect 24688 11150 24716 11630
rect 24768 11552 24820 11558
rect 24768 11494 24820 11500
rect 24492 11144 24544 11150
rect 24490 11112 24492 11121
rect 24676 11144 24728 11150
rect 24544 11112 24546 11121
rect 24676 11086 24728 11092
rect 24490 11047 24546 11056
rect 24584 11008 24636 11014
rect 24676 11008 24728 11014
rect 24584 10950 24636 10956
rect 24674 10976 24676 10985
rect 24728 10976 24730 10985
rect 24492 10464 24544 10470
rect 24492 10406 24544 10412
rect 24504 10266 24532 10406
rect 24492 10260 24544 10266
rect 24492 10202 24544 10208
rect 24398 9208 24454 9217
rect 24398 9143 24454 9152
rect 24400 9104 24452 9110
rect 24400 9046 24452 9052
rect 24306 8664 24362 8673
rect 24306 8599 24362 8608
rect 24136 8214 24256 8242
rect 24032 7880 24084 7886
rect 24032 7822 24084 7828
rect 23846 7168 23902 7177
rect 23846 7103 23902 7112
rect 23860 6934 23888 7103
rect 23848 6928 23900 6934
rect 23848 6870 23900 6876
rect 23756 4752 23808 4758
rect 23756 4694 23808 4700
rect 23572 4480 23624 4486
rect 23572 4422 23624 4428
rect 23756 4480 23808 4486
rect 23756 4422 23808 4428
rect 23940 4480 23992 4486
rect 23940 4422 23992 4428
rect 23584 4146 23612 4422
rect 23572 4140 23624 4146
rect 23572 4082 23624 4088
rect 23296 4072 23348 4078
rect 23296 4014 23348 4020
rect 23204 3936 23256 3942
rect 23204 3878 23256 3884
rect 23308 3534 23336 4014
rect 23768 3738 23796 4422
rect 23756 3732 23808 3738
rect 23756 3674 23808 3680
rect 23296 3528 23348 3534
rect 23296 3470 23348 3476
rect 23204 3460 23256 3466
rect 23204 3402 23256 3408
rect 23216 3194 23244 3402
rect 23664 3392 23716 3398
rect 23664 3334 23716 3340
rect 23204 3188 23256 3194
rect 23204 3130 23256 3136
rect 23676 3126 23704 3334
rect 23664 3120 23716 3126
rect 23664 3062 23716 3068
rect 23572 3052 23624 3058
rect 23572 2994 23624 3000
rect 23584 2961 23612 2994
rect 23952 2990 23980 4422
rect 24136 4282 24164 8214
rect 24216 5160 24268 5166
rect 24216 5102 24268 5108
rect 24124 4276 24176 4282
rect 24124 4218 24176 4224
rect 24124 3460 24176 3466
rect 24124 3402 24176 3408
rect 23940 2984 23992 2990
rect 23570 2952 23626 2961
rect 23940 2926 23992 2932
rect 23570 2887 23626 2896
rect 23848 2916 23900 2922
rect 23848 2858 23900 2864
rect 23296 2848 23348 2854
rect 23296 2790 23348 2796
rect 23388 2848 23440 2854
rect 23388 2790 23440 2796
rect 23308 800 23336 2790
rect 23400 2310 23428 2790
rect 23664 2440 23716 2446
rect 23664 2382 23716 2388
rect 23480 2372 23532 2378
rect 23532 2332 23612 2360
rect 23480 2314 23532 2320
rect 23388 2304 23440 2310
rect 23388 2246 23440 2252
rect 23584 800 23612 2332
rect 23676 1834 23704 2382
rect 23756 2372 23808 2378
rect 23756 2314 23808 2320
rect 23768 2038 23796 2314
rect 23756 2032 23808 2038
rect 23756 1974 23808 1980
rect 23664 1828 23716 1834
rect 23664 1770 23716 1776
rect 23860 800 23888 2858
rect 24136 800 24164 3402
rect 24228 2825 24256 5102
rect 24412 4593 24440 9046
rect 24504 8362 24532 10202
rect 24596 10062 24624 10950
rect 24674 10911 24730 10920
rect 24676 10464 24728 10470
rect 24676 10406 24728 10412
rect 24584 10056 24636 10062
rect 24584 9998 24636 10004
rect 24688 9722 24716 10406
rect 24780 10198 24808 11494
rect 24768 10192 24820 10198
rect 24768 10134 24820 10140
rect 24676 9716 24728 9722
rect 24676 9658 24728 9664
rect 24768 9376 24820 9382
rect 24768 9318 24820 9324
rect 24674 9072 24730 9081
rect 24674 9007 24730 9016
rect 24688 8401 24716 9007
rect 24674 8392 24730 8401
rect 24492 8356 24544 8362
rect 24674 8327 24730 8336
rect 24492 8298 24544 8304
rect 24676 6792 24728 6798
rect 24676 6734 24728 6740
rect 24688 6458 24716 6734
rect 24780 6730 24808 9318
rect 24768 6724 24820 6730
rect 24768 6666 24820 6672
rect 24676 6452 24728 6458
rect 24676 6394 24728 6400
rect 24872 5710 24900 12038
rect 24950 10840 25006 10849
rect 24950 10775 25006 10784
rect 25044 10804 25096 10810
rect 24964 10538 24992 10775
rect 25044 10746 25096 10752
rect 24952 10532 25004 10538
rect 24952 10474 25004 10480
rect 24952 9988 25004 9994
rect 24952 9930 25004 9936
rect 24964 9722 24992 9930
rect 24952 9716 25004 9722
rect 24952 9658 25004 9664
rect 25056 9674 25084 10746
rect 25148 10690 25176 12922
rect 25240 12306 25268 16351
rect 25318 15464 25374 15473
rect 25318 15399 25320 15408
rect 25372 15399 25374 15408
rect 25320 15370 25372 15376
rect 25516 15162 25544 19774
rect 25596 19440 25648 19446
rect 25596 19382 25648 19388
rect 25608 16998 25636 19382
rect 25596 16992 25648 16998
rect 25596 16934 25648 16940
rect 25700 15609 25728 20590
rect 25976 20505 26004 20742
rect 25962 20496 26018 20505
rect 26252 20466 26280 20878
rect 25962 20431 26018 20440
rect 26240 20460 26292 20466
rect 26240 20402 26292 20408
rect 25872 19780 25924 19786
rect 25872 19722 25924 19728
rect 25780 18760 25832 18766
rect 25780 18702 25832 18708
rect 25792 17542 25820 18702
rect 25780 17536 25832 17542
rect 25780 17478 25832 17484
rect 25686 15600 25742 15609
rect 25686 15535 25742 15544
rect 25504 15156 25556 15162
rect 25504 15098 25556 15104
rect 25700 15042 25728 15535
rect 25516 15014 25728 15042
rect 25412 14816 25464 14822
rect 25412 14758 25464 14764
rect 25424 14346 25452 14758
rect 25412 14340 25464 14346
rect 25412 14282 25464 14288
rect 25516 13852 25544 15014
rect 25688 14272 25740 14278
rect 25688 14214 25740 14220
rect 25700 13938 25728 14214
rect 25688 13932 25740 13938
rect 25688 13874 25740 13880
rect 25424 13824 25544 13852
rect 25424 13818 25452 13824
rect 25332 13790 25452 13818
rect 25228 12300 25280 12306
rect 25228 12242 25280 12248
rect 25240 11898 25268 12242
rect 25228 11892 25280 11898
rect 25228 11834 25280 11840
rect 25228 11756 25280 11762
rect 25228 11698 25280 11704
rect 25240 11354 25268 11698
rect 25228 11348 25280 11354
rect 25228 11290 25280 11296
rect 25148 10662 25268 10690
rect 25136 10260 25188 10266
rect 25136 10202 25188 10208
rect 25148 10062 25176 10202
rect 25136 10056 25188 10062
rect 25136 9998 25188 10004
rect 24964 8838 24992 9658
rect 25056 9646 25176 9674
rect 25044 9580 25096 9586
rect 25044 9522 25096 9528
rect 24952 8832 25004 8838
rect 24952 8774 25004 8780
rect 24950 8256 25006 8265
rect 24950 8191 25006 8200
rect 24964 7886 24992 8191
rect 24952 7880 25004 7886
rect 24952 7822 25004 7828
rect 25056 6322 25084 9522
rect 25148 8634 25176 9646
rect 25136 8628 25188 8634
rect 25136 8570 25188 8576
rect 25136 6656 25188 6662
rect 25136 6598 25188 6604
rect 25044 6316 25096 6322
rect 25044 6258 25096 6264
rect 24860 5704 24912 5710
rect 24860 5646 24912 5652
rect 24676 5024 24728 5030
rect 24676 4966 24728 4972
rect 24688 4826 24716 4966
rect 24676 4820 24728 4826
rect 24676 4762 24728 4768
rect 24492 4616 24544 4622
rect 24398 4584 24454 4593
rect 24492 4558 24544 4564
rect 24676 4616 24728 4622
rect 24676 4558 24728 4564
rect 24398 4519 24454 4528
rect 24504 4010 24532 4558
rect 24688 4282 24716 4558
rect 24676 4276 24728 4282
rect 24676 4218 24728 4224
rect 24872 4214 24900 5646
rect 25056 5386 25084 6258
rect 24964 5358 25084 5386
rect 24964 5234 24992 5358
rect 25148 5234 25176 6598
rect 24952 5228 25004 5234
rect 24952 5170 25004 5176
rect 25136 5228 25188 5234
rect 25136 5170 25188 5176
rect 24964 5030 24992 5170
rect 24952 5024 25004 5030
rect 24952 4966 25004 4972
rect 24964 4690 24992 4966
rect 25240 4758 25268 10662
rect 25332 10538 25360 13790
rect 25412 12844 25464 12850
rect 25412 12786 25464 12792
rect 25424 12442 25452 12786
rect 25504 12640 25556 12646
rect 25504 12582 25556 12588
rect 25516 12442 25544 12582
rect 25412 12436 25464 12442
rect 25412 12378 25464 12384
rect 25504 12436 25556 12442
rect 25504 12378 25556 12384
rect 25412 12164 25464 12170
rect 25412 12106 25464 12112
rect 25424 11830 25452 12106
rect 25516 12102 25544 12378
rect 25504 12096 25556 12102
rect 25504 12038 25556 12044
rect 25412 11824 25464 11830
rect 25412 11766 25464 11772
rect 25504 11756 25556 11762
rect 25504 11698 25556 11704
rect 25412 11688 25464 11694
rect 25412 11630 25464 11636
rect 25320 10532 25372 10538
rect 25320 10474 25372 10480
rect 25320 10192 25372 10198
rect 25320 10134 25372 10140
rect 25332 9217 25360 10134
rect 25424 9586 25452 11630
rect 25516 9586 25544 11698
rect 25596 11688 25648 11694
rect 25596 11630 25648 11636
rect 25608 10849 25636 11630
rect 25688 11280 25740 11286
rect 25688 11222 25740 11228
rect 25700 11082 25728 11222
rect 25688 11076 25740 11082
rect 25688 11018 25740 11024
rect 25594 10840 25650 10849
rect 25594 10775 25650 10784
rect 25792 9994 25820 17478
rect 25884 17270 25912 19722
rect 26056 19168 26108 19174
rect 26056 19110 26108 19116
rect 26068 18834 26096 19110
rect 26056 18828 26108 18834
rect 26056 18770 26108 18776
rect 26240 18148 26292 18154
rect 26240 18090 26292 18096
rect 26056 17740 26108 17746
rect 26108 17700 26188 17728
rect 26056 17682 26108 17688
rect 25872 17264 25924 17270
rect 25872 17206 25924 17212
rect 25964 17196 26016 17202
rect 25964 17138 26016 17144
rect 25976 16425 26004 17138
rect 25962 16416 26018 16425
rect 25962 16351 26018 16360
rect 25964 15428 26016 15434
rect 25964 15370 26016 15376
rect 25872 14952 25924 14958
rect 25872 14894 25924 14900
rect 25884 14414 25912 14894
rect 25976 14822 26004 15370
rect 26056 15156 26108 15162
rect 26056 15098 26108 15104
rect 25964 14816 26016 14822
rect 25964 14758 26016 14764
rect 25872 14408 25924 14414
rect 25872 14350 25924 14356
rect 25964 13796 26016 13802
rect 25964 13738 26016 13744
rect 25872 12640 25924 12646
rect 25872 12582 25924 12588
rect 25884 12238 25912 12582
rect 25872 12232 25924 12238
rect 25872 12174 25924 12180
rect 25976 10996 26004 13738
rect 26068 11529 26096 15098
rect 26160 14482 26188 17700
rect 26252 17678 26280 18090
rect 26240 17672 26292 17678
rect 26240 17614 26292 17620
rect 26252 16810 26280 17614
rect 26344 16946 26372 35866
rect 26896 26926 26924 41414
rect 26976 33924 27028 33930
rect 26976 33866 27028 33872
rect 26884 26920 26936 26926
rect 26884 26862 26936 26868
rect 26988 24138 27016 33866
rect 28368 27130 28396 60998
rect 28460 60110 28488 61610
rect 28828 60790 28856 63200
rect 29840 61198 29868 63294
rect 30286 63200 30342 64000
rect 31022 63322 31078 64000
rect 31022 63294 31248 63322
rect 31022 63200 31078 63294
rect 30104 61804 30156 61810
rect 30104 61746 30156 61752
rect 29828 61192 29880 61198
rect 29828 61134 29880 61140
rect 29920 61056 29972 61062
rect 29920 60998 29972 61004
rect 28816 60784 28868 60790
rect 28816 60726 28868 60732
rect 29000 60512 29052 60518
rect 29000 60454 29052 60460
rect 29828 60512 29880 60518
rect 29828 60454 29880 60460
rect 29012 60178 29040 60454
rect 29000 60172 29052 60178
rect 29000 60114 29052 60120
rect 28448 60104 28500 60110
rect 28448 60046 28500 60052
rect 28540 59968 28592 59974
rect 28540 59910 28592 59916
rect 28724 59968 28776 59974
rect 28724 59910 28776 59916
rect 28448 59628 28500 59634
rect 28448 59570 28500 59576
rect 28460 36854 28488 59570
rect 28552 59566 28580 59910
rect 28630 59664 28686 59673
rect 28630 59599 28686 59608
rect 28644 59566 28672 59599
rect 28540 59560 28592 59566
rect 28540 59502 28592 59508
rect 28632 59560 28684 59566
rect 28632 59502 28684 59508
rect 28736 54738 28764 59910
rect 29840 59634 29868 60454
rect 29736 59628 29788 59634
rect 29736 59570 29788 59576
rect 29828 59628 29880 59634
rect 29828 59570 29880 59576
rect 29748 59430 29776 59570
rect 29736 59424 29788 59430
rect 29736 59366 29788 59372
rect 29368 57044 29420 57050
rect 29368 56986 29420 56992
rect 29380 56370 29408 56986
rect 29368 56364 29420 56370
rect 29368 56306 29420 56312
rect 29736 56296 29788 56302
rect 29736 56238 29788 56244
rect 29000 56160 29052 56166
rect 29000 56102 29052 56108
rect 28724 54732 28776 54738
rect 28724 54674 28776 54680
rect 28448 36848 28500 36854
rect 28448 36790 28500 36796
rect 28356 27124 28408 27130
rect 28356 27066 28408 27072
rect 27804 26920 27856 26926
rect 27804 26862 27856 26868
rect 27252 26852 27304 26858
rect 27252 26794 27304 26800
rect 26700 24132 26752 24138
rect 26700 24074 26752 24080
rect 26976 24132 27028 24138
rect 26976 24074 27028 24080
rect 26712 23322 26740 24074
rect 26700 23316 26752 23322
rect 26700 23258 26752 23264
rect 26608 23180 26660 23186
rect 26608 23122 26660 23128
rect 26516 18760 26568 18766
rect 26516 18702 26568 18708
rect 26528 18601 26556 18702
rect 26514 18592 26570 18601
rect 26514 18527 26570 18536
rect 26516 18080 26568 18086
rect 26516 18022 26568 18028
rect 26528 17202 26556 18022
rect 26424 17196 26476 17202
rect 26424 17138 26476 17144
rect 26516 17196 26568 17202
rect 26516 17138 26568 17144
rect 26436 17048 26464 17138
rect 26436 17020 26556 17048
rect 26344 16918 26464 16946
rect 26252 16794 26372 16810
rect 26252 16788 26384 16794
rect 26252 16782 26332 16788
rect 26332 16730 26384 16736
rect 26240 16448 26292 16454
rect 26240 16390 26292 16396
rect 26148 14476 26200 14482
rect 26148 14418 26200 14424
rect 26160 13977 26188 14418
rect 26146 13968 26202 13977
rect 26146 13903 26202 13912
rect 26252 13734 26280 16390
rect 26344 15570 26372 16730
rect 26332 15564 26384 15570
rect 26332 15506 26384 15512
rect 26344 15094 26372 15506
rect 26332 15088 26384 15094
rect 26332 15030 26384 15036
rect 26332 14816 26384 14822
rect 26332 14758 26384 14764
rect 26344 14346 26372 14758
rect 26436 14482 26464 16918
rect 26424 14476 26476 14482
rect 26424 14418 26476 14424
rect 26332 14340 26384 14346
rect 26332 14282 26384 14288
rect 26240 13728 26292 13734
rect 26240 13670 26292 13676
rect 26148 12980 26200 12986
rect 26148 12922 26200 12928
rect 26240 12980 26292 12986
rect 26240 12922 26292 12928
rect 26160 12850 26188 12922
rect 26148 12844 26200 12850
rect 26148 12786 26200 12792
rect 26252 11762 26280 12922
rect 26240 11756 26292 11762
rect 26240 11698 26292 11704
rect 26054 11520 26110 11529
rect 26054 11455 26110 11464
rect 26148 11348 26200 11354
rect 26148 11290 26200 11296
rect 26056 11280 26108 11286
rect 26056 11222 26108 11228
rect 26068 11150 26096 11222
rect 26160 11150 26188 11290
rect 26056 11144 26108 11150
rect 26056 11086 26108 11092
rect 26148 11144 26200 11150
rect 26148 11086 26200 11092
rect 25976 10968 26188 10996
rect 25872 10668 25924 10674
rect 25872 10610 25924 10616
rect 25596 9988 25648 9994
rect 25596 9930 25648 9936
rect 25780 9988 25832 9994
rect 25780 9930 25832 9936
rect 25608 9761 25636 9930
rect 25778 9888 25834 9897
rect 25778 9823 25834 9832
rect 25594 9752 25650 9761
rect 25594 9687 25650 9696
rect 25412 9580 25464 9586
rect 25412 9522 25464 9528
rect 25504 9580 25556 9586
rect 25504 9522 25556 9528
rect 25318 9208 25374 9217
rect 25318 9143 25374 9152
rect 25332 8974 25360 9143
rect 25320 8968 25372 8974
rect 25320 8910 25372 8916
rect 25424 8430 25452 9522
rect 25516 9353 25544 9522
rect 25502 9344 25558 9353
rect 25502 9279 25558 9288
rect 25412 8424 25464 8430
rect 25412 8366 25464 8372
rect 25228 4752 25280 4758
rect 25228 4694 25280 4700
rect 24952 4684 25004 4690
rect 24952 4626 25004 4632
rect 25424 4622 25452 8366
rect 25412 4616 25464 4622
rect 25412 4558 25464 4564
rect 25516 4554 25544 9279
rect 25792 8974 25820 9823
rect 25884 9586 25912 10610
rect 25964 10600 26016 10606
rect 25964 10542 26016 10548
rect 25976 9586 26004 10542
rect 26056 10532 26108 10538
rect 26056 10474 26108 10480
rect 26068 10441 26096 10474
rect 26054 10432 26110 10441
rect 26054 10367 26110 10376
rect 25872 9580 25924 9586
rect 25872 9522 25924 9528
rect 25964 9580 26016 9586
rect 25964 9522 26016 9528
rect 25884 9110 25912 9522
rect 25872 9104 25924 9110
rect 25872 9046 25924 9052
rect 25688 8968 25740 8974
rect 25688 8910 25740 8916
rect 25780 8968 25832 8974
rect 25780 8910 25832 8916
rect 25700 7857 25728 8910
rect 25792 8430 25820 8910
rect 25780 8424 25832 8430
rect 25780 8366 25832 8372
rect 25686 7848 25742 7857
rect 25686 7783 25742 7792
rect 25688 7200 25740 7206
rect 25688 7142 25740 7148
rect 25596 6724 25648 6730
rect 25596 6666 25648 6672
rect 25608 6458 25636 6666
rect 25700 6458 25728 7142
rect 25596 6452 25648 6458
rect 25596 6394 25648 6400
rect 25688 6452 25740 6458
rect 25688 6394 25740 6400
rect 25884 5250 25912 9046
rect 25976 9042 26004 9522
rect 25964 9036 26016 9042
rect 25964 8978 26016 8984
rect 26160 8537 26188 10968
rect 26252 10130 26280 11698
rect 26240 10124 26292 10130
rect 26240 10066 26292 10072
rect 26344 8906 26372 14282
rect 26424 14068 26476 14074
rect 26528 14056 26556 17020
rect 26620 14414 26648 23122
rect 26976 20868 27028 20874
rect 26976 20810 27028 20816
rect 26700 20800 26752 20806
rect 26700 20742 26752 20748
rect 26712 20534 26740 20742
rect 26700 20528 26752 20534
rect 26700 20470 26752 20476
rect 26988 19530 27016 20810
rect 27160 20460 27212 20466
rect 27160 20402 27212 20408
rect 26804 19502 27016 19530
rect 26700 18896 26752 18902
rect 26700 18838 26752 18844
rect 26712 17678 26740 18838
rect 26804 18630 26832 19502
rect 26976 19372 27028 19378
rect 26976 19314 27028 19320
rect 26792 18624 26844 18630
rect 26792 18566 26844 18572
rect 26884 18624 26936 18630
rect 26884 18566 26936 18572
rect 26700 17672 26752 17678
rect 26700 17614 26752 17620
rect 26896 16998 26924 18566
rect 26988 18358 27016 19314
rect 27068 18896 27120 18902
rect 27068 18838 27120 18844
rect 26976 18352 27028 18358
rect 26976 18294 27028 18300
rect 27080 18290 27108 18838
rect 27172 18290 27200 20402
rect 27068 18284 27120 18290
rect 27068 18226 27120 18232
rect 27160 18284 27212 18290
rect 27160 18226 27212 18232
rect 27172 18154 27200 18226
rect 27160 18148 27212 18154
rect 27160 18090 27212 18096
rect 27264 17610 27292 26794
rect 27436 25492 27488 25498
rect 27436 25434 27488 25440
rect 27344 17808 27396 17814
rect 27344 17750 27396 17756
rect 27252 17604 27304 17610
rect 27252 17546 27304 17552
rect 27356 17338 27384 17750
rect 27344 17332 27396 17338
rect 27344 17274 27396 17280
rect 26884 16992 26936 16998
rect 26884 16934 26936 16940
rect 26884 16788 26936 16794
rect 26884 16730 26936 16736
rect 26792 16584 26844 16590
rect 26792 16526 26844 16532
rect 26804 16182 26832 16526
rect 26792 16176 26844 16182
rect 26792 16118 26844 16124
rect 26698 15328 26754 15337
rect 26698 15263 26754 15272
rect 26608 14408 26660 14414
rect 26608 14350 26660 14356
rect 26476 14028 26556 14056
rect 26424 14010 26476 14016
rect 26516 13932 26568 13938
rect 26516 13874 26568 13880
rect 26424 13864 26476 13870
rect 26424 13806 26476 13812
rect 26436 13530 26464 13806
rect 26424 13524 26476 13530
rect 26424 13466 26476 13472
rect 26528 12374 26556 13874
rect 26608 12640 26660 12646
rect 26608 12582 26660 12588
rect 26516 12368 26568 12374
rect 26516 12310 26568 12316
rect 26424 11756 26476 11762
rect 26424 11698 26476 11704
rect 26436 10810 26464 11698
rect 26424 10804 26476 10810
rect 26424 10746 26476 10752
rect 26528 10266 26556 12310
rect 26620 11370 26648 12582
rect 26712 11558 26740 15263
rect 26792 12164 26844 12170
rect 26792 12106 26844 12112
rect 26804 11898 26832 12106
rect 26896 12102 26924 16730
rect 27068 16652 27120 16658
rect 27068 16594 27120 16600
rect 27080 16454 27108 16594
rect 27068 16448 27120 16454
rect 27068 16390 27120 16396
rect 27080 16250 27108 16390
rect 27068 16244 27120 16250
rect 27068 16186 27120 16192
rect 27344 15564 27396 15570
rect 27344 15506 27396 15512
rect 27160 14476 27212 14482
rect 27160 14418 27212 14424
rect 27172 14278 27200 14418
rect 27252 14408 27304 14414
rect 27252 14350 27304 14356
rect 27160 14272 27212 14278
rect 27160 14214 27212 14220
rect 27264 13870 27292 14350
rect 27252 13864 27304 13870
rect 27252 13806 27304 13812
rect 27356 13530 27384 15506
rect 27344 13524 27396 13530
rect 27344 13466 27396 13472
rect 27068 12708 27120 12714
rect 27068 12650 27120 12656
rect 26974 12336 27030 12345
rect 26974 12271 26976 12280
rect 27028 12271 27030 12280
rect 26976 12242 27028 12248
rect 26884 12096 26936 12102
rect 26884 12038 26936 12044
rect 26792 11892 26844 11898
rect 26792 11834 26844 11840
rect 26700 11552 26752 11558
rect 26700 11494 26752 11500
rect 26620 11342 26740 11370
rect 26516 10260 26568 10266
rect 26516 10202 26568 10208
rect 26422 9616 26478 9625
rect 26422 9551 26478 9560
rect 26436 8974 26464 9551
rect 26424 8968 26476 8974
rect 26424 8910 26476 8916
rect 26332 8900 26384 8906
rect 26332 8842 26384 8848
rect 26146 8528 26202 8537
rect 26146 8463 26202 8472
rect 26240 8084 26292 8090
rect 26240 8026 26292 8032
rect 26252 6322 26280 8026
rect 26436 6730 26464 8910
rect 26528 8838 26556 10202
rect 26606 9616 26662 9625
rect 26606 9551 26662 9560
rect 26620 9518 26648 9551
rect 26608 9512 26660 9518
rect 26608 9454 26660 9460
rect 26516 8832 26568 8838
rect 26516 8774 26568 8780
rect 26712 8401 26740 11342
rect 26884 10124 26936 10130
rect 26884 10066 26936 10072
rect 26698 8392 26754 8401
rect 26698 8327 26754 8336
rect 26792 6860 26844 6866
rect 26792 6802 26844 6808
rect 26424 6724 26476 6730
rect 26424 6666 26476 6672
rect 26516 6656 26568 6662
rect 26516 6598 26568 6604
rect 26240 6316 26292 6322
rect 26240 6258 26292 6264
rect 26056 6248 26108 6254
rect 26056 6190 26108 6196
rect 26424 6248 26476 6254
rect 26424 6190 26476 6196
rect 26068 5370 26096 6190
rect 26240 5908 26292 5914
rect 26240 5850 26292 5856
rect 26252 5817 26280 5850
rect 26238 5808 26294 5817
rect 26238 5743 26294 5752
rect 26056 5364 26108 5370
rect 26056 5306 26108 5312
rect 26436 5302 26464 6190
rect 26528 5574 26556 6598
rect 26608 6316 26660 6322
rect 26608 6258 26660 6264
rect 26620 5846 26648 6258
rect 26608 5840 26660 5846
rect 26608 5782 26660 5788
rect 26608 5704 26660 5710
rect 26608 5646 26660 5652
rect 26516 5568 26568 5574
rect 26516 5510 26568 5516
rect 26424 5296 26476 5302
rect 25884 5222 26096 5250
rect 26424 5238 26476 5244
rect 25780 5024 25832 5030
rect 25780 4966 25832 4972
rect 25872 5024 25924 5030
rect 25872 4966 25924 4972
rect 25596 4820 25648 4826
rect 25596 4762 25648 4768
rect 25608 4554 25636 4762
rect 25504 4548 25556 4554
rect 25504 4490 25556 4496
rect 25596 4548 25648 4554
rect 25596 4490 25648 4496
rect 24860 4208 24912 4214
rect 24860 4150 24912 4156
rect 24676 4072 24728 4078
rect 24676 4014 24728 4020
rect 24492 4004 24544 4010
rect 24492 3946 24544 3952
rect 24214 2816 24270 2825
rect 24214 2751 24270 2760
rect 24400 2508 24452 2514
rect 24400 2450 24452 2456
rect 24412 800 24440 2450
rect 24688 800 24716 4014
rect 24872 3641 24900 4150
rect 24858 3632 24914 3641
rect 24858 3567 24914 3576
rect 25228 2916 25280 2922
rect 25228 2858 25280 2864
rect 24952 2372 25004 2378
rect 24952 2314 25004 2320
rect 24964 800 24992 2314
rect 25240 800 25268 2858
rect 25504 2372 25556 2378
rect 25504 2314 25556 2320
rect 25516 800 25544 2314
rect 25792 800 25820 4966
rect 25884 4758 25912 4966
rect 25872 4752 25924 4758
rect 25872 4694 25924 4700
rect 25964 4752 26016 4758
rect 25964 4694 26016 4700
rect 25976 4622 26004 4694
rect 25964 4616 26016 4622
rect 25964 4558 26016 4564
rect 25964 3936 26016 3942
rect 25964 3878 26016 3884
rect 25976 1034 26004 3878
rect 26068 1766 26096 5222
rect 26332 5160 26384 5166
rect 26332 5102 26384 5108
rect 26344 4758 26372 5102
rect 26332 4752 26384 4758
rect 26332 4694 26384 4700
rect 26436 4622 26464 5238
rect 26528 5166 26556 5510
rect 26516 5160 26568 5166
rect 26516 5102 26568 5108
rect 26424 4616 26476 4622
rect 26424 4558 26476 4564
rect 26240 4548 26292 4554
rect 26240 4490 26292 4496
rect 26252 2774 26280 4490
rect 26516 3528 26568 3534
rect 26516 3470 26568 3476
rect 26528 3126 26556 3470
rect 26516 3120 26568 3126
rect 26516 3062 26568 3068
rect 26424 2984 26476 2990
rect 26424 2926 26476 2932
rect 26252 2746 26372 2774
rect 26148 2304 26200 2310
rect 26148 2246 26200 2252
rect 26056 1760 26108 1766
rect 26056 1702 26108 1708
rect 26160 1426 26188 2246
rect 26148 1420 26200 1426
rect 26148 1362 26200 1368
rect 25976 1006 26096 1034
rect 26068 800 26096 1006
rect 26344 800 26372 2746
rect 26436 1562 26464 2926
rect 26424 1556 26476 1562
rect 26424 1498 26476 1504
rect 26620 800 26648 5646
rect 26700 3460 26752 3466
rect 26700 3402 26752 3408
rect 26712 1970 26740 3402
rect 26804 2650 26832 6802
rect 26896 6254 26924 10066
rect 27080 9178 27108 12650
rect 27356 12345 27384 13466
rect 27448 12850 27476 25434
rect 27528 21616 27580 21622
rect 27528 21558 27580 21564
rect 27540 21010 27568 21558
rect 27712 21548 27764 21554
rect 27712 21490 27764 21496
rect 27620 21140 27672 21146
rect 27620 21082 27672 21088
rect 27528 21004 27580 21010
rect 27528 20946 27580 20952
rect 27632 19922 27660 21082
rect 27724 20942 27752 21490
rect 27712 20936 27764 20942
rect 27712 20878 27764 20884
rect 27724 20602 27752 20878
rect 27712 20596 27764 20602
rect 27712 20538 27764 20544
rect 27620 19916 27672 19922
rect 27620 19858 27672 19864
rect 27620 17536 27672 17542
rect 27620 17478 27672 17484
rect 27528 17196 27580 17202
rect 27528 17138 27580 17144
rect 27540 16969 27568 17138
rect 27526 16960 27582 16969
rect 27526 16895 27582 16904
rect 27528 15360 27580 15366
rect 27632 15348 27660 17478
rect 27816 17270 27844 26862
rect 28460 26314 28488 36790
rect 29012 27577 29040 56102
rect 29748 55758 29776 56238
rect 29736 55752 29788 55758
rect 29736 55694 29788 55700
rect 29932 50454 29960 60998
rect 30012 60036 30064 60042
rect 30012 59978 30064 59984
rect 30024 59634 30052 59978
rect 30116 59702 30144 61746
rect 30300 60874 30328 63200
rect 31220 61198 31248 63294
rect 31758 63200 31814 64000
rect 32494 63322 32550 64000
rect 33230 63322 33286 64000
rect 33966 63322 34022 64000
rect 32494 63294 32904 63322
rect 32494 63200 32550 63294
rect 31772 61198 31800 63200
rect 32876 61198 32904 63294
rect 33230 63294 33548 63322
rect 33230 63200 33286 63294
rect 33416 61736 33468 61742
rect 33416 61678 33468 61684
rect 31208 61192 31260 61198
rect 31208 61134 31260 61140
rect 31760 61192 31812 61198
rect 31760 61134 31812 61140
rect 32864 61192 32916 61198
rect 32864 61134 32916 61140
rect 33140 61124 33192 61130
rect 33140 61066 33192 61072
rect 31300 61056 31352 61062
rect 31300 60998 31352 61004
rect 32588 61056 32640 61062
rect 32588 60998 32640 61004
rect 30300 60846 30420 60874
rect 30392 60790 30420 60846
rect 30380 60784 30432 60790
rect 30380 60726 30432 60732
rect 30564 60512 30616 60518
rect 30564 60454 30616 60460
rect 30196 60240 30248 60246
rect 30196 60182 30248 60188
rect 30104 59696 30156 59702
rect 30104 59638 30156 59644
rect 30208 59634 30236 60182
rect 30380 60104 30432 60110
rect 30378 60072 30380 60081
rect 30432 60072 30434 60081
rect 30378 60007 30434 60016
rect 30576 59634 30604 60454
rect 30656 60036 30708 60042
rect 30656 59978 30708 59984
rect 30668 59945 30696 59978
rect 31024 59968 31076 59974
rect 30654 59936 30710 59945
rect 31024 59910 31076 59916
rect 30654 59871 30710 59880
rect 30012 59628 30064 59634
rect 30012 59570 30064 59576
rect 30196 59628 30248 59634
rect 30196 59570 30248 59576
rect 30564 59628 30616 59634
rect 30564 59570 30616 59576
rect 30104 59560 30156 59566
rect 30656 59560 30708 59566
rect 30156 59508 30604 59514
rect 30104 59502 30604 59508
rect 30656 59502 30708 59508
rect 30116 59498 30604 59502
rect 30116 59492 30616 59498
rect 30116 59486 30564 59492
rect 30564 59434 30616 59440
rect 30288 59424 30340 59430
rect 30472 59424 30524 59430
rect 30340 59372 30472 59378
rect 30288 59366 30524 59372
rect 30300 59350 30512 59366
rect 30668 57050 30696 59502
rect 30656 57044 30708 57050
rect 30656 56986 30708 56992
rect 31036 55826 31064 59910
rect 31024 55820 31076 55826
rect 31024 55762 31076 55768
rect 29920 50448 29972 50454
rect 29920 50390 29972 50396
rect 29828 50380 29880 50386
rect 29828 50322 29880 50328
rect 29736 37868 29788 37874
rect 29736 37810 29788 37816
rect 29748 35766 29776 37810
rect 29736 35760 29788 35766
rect 29736 35702 29788 35708
rect 29184 32428 29236 32434
rect 29184 32370 29236 32376
rect 29092 30932 29144 30938
rect 29092 30874 29144 30880
rect 29104 28558 29132 30874
rect 29092 28552 29144 28558
rect 29092 28494 29144 28500
rect 28998 27568 29054 27577
rect 28998 27503 29054 27512
rect 28448 26308 28500 26314
rect 28448 26250 28500 26256
rect 28632 21956 28684 21962
rect 28632 21898 28684 21904
rect 28540 21888 28592 21894
rect 28540 21830 28592 21836
rect 27896 21480 27948 21486
rect 27896 21422 27948 21428
rect 27988 21480 28040 21486
rect 27988 21422 28040 21428
rect 27908 21146 27936 21422
rect 27896 21140 27948 21146
rect 27896 21082 27948 21088
rect 28000 21010 28028 21422
rect 28264 21412 28316 21418
rect 28264 21354 28316 21360
rect 27988 21004 28040 21010
rect 27988 20946 28040 20952
rect 27896 17672 27948 17678
rect 27896 17614 27948 17620
rect 27804 17264 27856 17270
rect 27804 17206 27856 17212
rect 27908 17202 27936 17614
rect 27896 17196 27948 17202
rect 27896 17138 27948 17144
rect 27896 16584 27948 16590
rect 27894 16552 27896 16561
rect 27948 16552 27950 16561
rect 27894 16487 27950 16496
rect 27908 16182 27936 16487
rect 27896 16176 27948 16182
rect 27896 16118 27948 16124
rect 28000 16046 28028 20946
rect 28172 20596 28224 20602
rect 28172 20538 28224 20544
rect 28184 17678 28212 20538
rect 28276 20330 28304 21354
rect 28356 21344 28408 21350
rect 28356 21286 28408 21292
rect 28368 21010 28396 21286
rect 28356 21004 28408 21010
rect 28356 20946 28408 20952
rect 28448 20800 28500 20806
rect 28448 20742 28500 20748
rect 28264 20324 28316 20330
rect 28264 20266 28316 20272
rect 28356 19168 28408 19174
rect 28356 19110 28408 19116
rect 28368 18970 28396 19110
rect 28356 18964 28408 18970
rect 28356 18906 28408 18912
rect 28264 18828 28316 18834
rect 28264 18770 28316 18776
rect 28356 18828 28408 18834
rect 28356 18770 28408 18776
rect 28276 18290 28304 18770
rect 28368 18698 28396 18770
rect 28356 18692 28408 18698
rect 28356 18634 28408 18640
rect 28264 18284 28316 18290
rect 28264 18226 28316 18232
rect 28080 17672 28132 17678
rect 28080 17614 28132 17620
rect 28172 17672 28224 17678
rect 28172 17614 28224 17620
rect 27712 16040 27764 16046
rect 27712 15982 27764 15988
rect 27988 16040 28040 16046
rect 27988 15982 28040 15988
rect 27724 15910 27752 15982
rect 27712 15904 27764 15910
rect 27712 15846 27764 15852
rect 27580 15320 27660 15348
rect 27528 15302 27580 15308
rect 27540 15094 27568 15302
rect 27528 15088 27580 15094
rect 27528 15030 27580 15036
rect 27540 13938 27568 15030
rect 27620 15020 27672 15026
rect 27620 14962 27672 14968
rect 27896 15020 27948 15026
rect 27896 14962 27948 14968
rect 27632 14618 27660 14962
rect 27712 14952 27764 14958
rect 27712 14894 27764 14900
rect 27724 14618 27752 14894
rect 27620 14612 27672 14618
rect 27620 14554 27672 14560
rect 27712 14612 27764 14618
rect 27712 14554 27764 14560
rect 27528 13932 27580 13938
rect 27528 13874 27580 13880
rect 27908 13530 27936 14962
rect 28000 14958 28028 15982
rect 27988 14952 28040 14958
rect 27988 14894 28040 14900
rect 27988 14340 28040 14346
rect 27988 14282 28040 14288
rect 28000 13954 28028 14282
rect 28092 14074 28120 17614
rect 28170 17368 28226 17377
rect 28170 17303 28226 17312
rect 28080 14068 28132 14074
rect 28080 14010 28132 14016
rect 28000 13926 28120 13954
rect 27896 13524 27948 13530
rect 27896 13466 27948 13472
rect 27618 13152 27674 13161
rect 27618 13087 27674 13096
rect 27632 12850 27660 13087
rect 27804 12912 27856 12918
rect 27804 12854 27856 12860
rect 27436 12844 27488 12850
rect 27436 12786 27488 12792
rect 27620 12844 27672 12850
rect 27620 12786 27672 12792
rect 27342 12336 27398 12345
rect 27342 12271 27398 12280
rect 27342 11792 27398 11801
rect 27342 11727 27398 11736
rect 27356 11694 27384 11727
rect 27448 11694 27476 12786
rect 27712 12640 27764 12646
rect 27712 12582 27764 12588
rect 27344 11688 27396 11694
rect 27344 11630 27396 11636
rect 27436 11688 27488 11694
rect 27436 11630 27488 11636
rect 27724 11200 27752 12582
rect 27816 11354 27844 12854
rect 27804 11348 27856 11354
rect 27804 11290 27856 11296
rect 27632 11172 27752 11200
rect 27342 11112 27398 11121
rect 27342 11047 27398 11056
rect 27252 10532 27304 10538
rect 27252 10474 27304 10480
rect 27264 10441 27292 10474
rect 27250 10432 27306 10441
rect 27250 10367 27306 10376
rect 27264 10062 27292 10367
rect 27252 10056 27304 10062
rect 27252 9998 27304 10004
rect 27158 9344 27214 9353
rect 27158 9279 27214 9288
rect 27068 9172 27120 9178
rect 27068 9114 27120 9120
rect 26976 8832 27028 8838
rect 26976 8774 27028 8780
rect 26884 6248 26936 6254
rect 26884 6190 26936 6196
rect 26884 5160 26936 5166
rect 26884 5102 26936 5108
rect 26896 3398 26924 5102
rect 26884 3392 26936 3398
rect 26884 3334 26936 3340
rect 26792 2644 26844 2650
rect 26792 2586 26844 2592
rect 26884 2304 26936 2310
rect 26884 2246 26936 2252
rect 26700 1964 26752 1970
rect 26700 1906 26752 1912
rect 26896 800 26924 2246
rect 26988 1970 27016 8774
rect 27080 6866 27108 9114
rect 27172 8498 27200 9279
rect 27160 8492 27212 8498
rect 27160 8434 27212 8440
rect 27172 7002 27200 8434
rect 27160 6996 27212 7002
rect 27160 6938 27212 6944
rect 27068 6860 27120 6866
rect 27068 6802 27120 6808
rect 27160 6316 27212 6322
rect 27160 6258 27212 6264
rect 27172 5953 27200 6258
rect 27158 5944 27214 5953
rect 27158 5879 27214 5888
rect 27264 5234 27292 9998
rect 27356 8022 27384 11047
rect 27632 10742 27660 11172
rect 27802 11112 27858 11121
rect 27712 11076 27764 11082
rect 27802 11047 27858 11056
rect 27712 11018 27764 11024
rect 27620 10736 27672 10742
rect 27620 10678 27672 10684
rect 27632 10112 27660 10678
rect 27448 10084 27660 10112
rect 27448 9042 27476 10084
rect 27618 10024 27674 10033
rect 27618 9959 27620 9968
rect 27672 9959 27674 9968
rect 27620 9930 27672 9936
rect 27620 9580 27672 9586
rect 27724 9568 27752 11018
rect 27816 10606 27844 11047
rect 27804 10600 27856 10606
rect 27804 10542 27856 10548
rect 27804 10464 27856 10470
rect 27804 10406 27856 10412
rect 27816 9625 27844 10406
rect 27894 10160 27950 10169
rect 27894 10095 27950 10104
rect 27672 9540 27752 9568
rect 27802 9616 27858 9625
rect 27802 9551 27858 9560
rect 27620 9522 27672 9528
rect 27528 9444 27580 9450
rect 27528 9386 27580 9392
rect 27540 9353 27568 9386
rect 27526 9344 27582 9353
rect 27526 9279 27582 9288
rect 27908 9042 27936 10095
rect 27988 10056 28040 10062
rect 27988 9998 28040 10004
rect 28000 9178 28028 9998
rect 27988 9172 28040 9178
rect 27988 9114 28040 9120
rect 27436 9036 27488 9042
rect 27436 8978 27488 8984
rect 27896 9036 27948 9042
rect 27896 8978 27948 8984
rect 27804 8968 27856 8974
rect 27988 8968 28040 8974
rect 27804 8910 27856 8916
rect 27986 8936 27988 8945
rect 28040 8936 28042 8945
rect 27436 8900 27488 8906
rect 27436 8842 27488 8848
rect 27344 8016 27396 8022
rect 27344 7958 27396 7964
rect 27344 7472 27396 7478
rect 27448 7426 27476 8842
rect 27528 8492 27580 8498
rect 27528 8434 27580 8440
rect 27396 7420 27476 7426
rect 27344 7414 27476 7420
rect 27356 7398 27476 7414
rect 27540 7410 27568 8434
rect 27712 8424 27764 8430
rect 27712 8366 27764 8372
rect 27620 8288 27672 8294
rect 27620 8230 27672 8236
rect 27632 7478 27660 8230
rect 27620 7472 27672 7478
rect 27620 7414 27672 7420
rect 27448 7154 27476 7398
rect 27528 7404 27580 7410
rect 27528 7346 27580 7352
rect 27526 7168 27582 7177
rect 27448 7126 27526 7154
rect 27526 7103 27582 7112
rect 27540 6254 27568 7103
rect 27528 6248 27580 6254
rect 27528 6190 27580 6196
rect 27528 6112 27580 6118
rect 27528 6054 27580 6060
rect 27160 5228 27212 5234
rect 27160 5170 27212 5176
rect 27252 5228 27304 5234
rect 27252 5170 27304 5176
rect 27172 4729 27200 5170
rect 27540 5030 27568 6054
rect 27632 5574 27660 7414
rect 27724 7002 27752 8366
rect 27816 7546 27844 8910
rect 27986 8871 28042 8880
rect 27988 8832 28040 8838
rect 27988 8774 28040 8780
rect 27804 7540 27856 7546
rect 27804 7482 27856 7488
rect 27712 6996 27764 7002
rect 27712 6938 27764 6944
rect 27896 6996 27948 7002
rect 27896 6938 27948 6944
rect 27712 6860 27764 6866
rect 27712 6802 27764 6808
rect 27620 5568 27672 5574
rect 27620 5510 27672 5516
rect 27618 5128 27674 5137
rect 27618 5063 27674 5072
rect 27528 5024 27580 5030
rect 27528 4966 27580 4972
rect 27158 4720 27214 4729
rect 27158 4655 27214 4664
rect 27068 4548 27120 4554
rect 27068 4490 27120 4496
rect 27080 3777 27108 4490
rect 27066 3768 27122 3777
rect 27066 3703 27122 3712
rect 27172 3097 27200 4655
rect 27252 4004 27304 4010
rect 27304 3964 27384 3992
rect 27252 3946 27304 3952
rect 27250 3496 27306 3505
rect 27356 3466 27384 3964
rect 27540 3618 27568 4966
rect 27632 4554 27660 5063
rect 27724 4826 27752 6802
rect 27804 6724 27856 6730
rect 27804 6666 27856 6672
rect 27816 5817 27844 6666
rect 27802 5808 27858 5817
rect 27802 5743 27858 5752
rect 27712 4820 27764 4826
rect 27712 4762 27764 4768
rect 27620 4548 27672 4554
rect 27620 4490 27672 4496
rect 27804 4276 27856 4282
rect 27804 4218 27856 4224
rect 27710 3768 27766 3777
rect 27710 3703 27712 3712
rect 27764 3703 27766 3712
rect 27712 3674 27764 3680
rect 27448 3602 27568 3618
rect 27436 3596 27568 3602
rect 27488 3590 27568 3596
rect 27436 3538 27488 3544
rect 27250 3431 27252 3440
rect 27304 3431 27306 3440
rect 27344 3460 27396 3466
rect 27252 3402 27304 3408
rect 27344 3402 27396 3408
rect 27448 3346 27476 3538
rect 27356 3318 27476 3346
rect 27158 3088 27214 3097
rect 27356 3058 27384 3318
rect 27436 3188 27488 3194
rect 27436 3130 27488 3136
rect 27158 3023 27214 3032
rect 27344 3052 27396 3058
rect 27344 2994 27396 3000
rect 27160 2848 27212 2854
rect 27160 2790 27212 2796
rect 26976 1964 27028 1970
rect 26976 1906 27028 1912
rect 27172 800 27200 2790
rect 27448 800 27476 3130
rect 27526 3088 27582 3097
rect 27526 3023 27528 3032
rect 27580 3023 27582 3032
rect 27528 2994 27580 3000
rect 27816 2774 27844 4218
rect 27724 2746 27844 2774
rect 27724 800 27752 2746
rect 27908 2553 27936 6938
rect 28000 6798 28028 8774
rect 28092 6866 28120 13926
rect 28184 12646 28212 17303
rect 28276 16658 28304 18226
rect 28356 17264 28408 17270
rect 28356 17206 28408 17212
rect 28264 16652 28316 16658
rect 28264 16594 28316 16600
rect 28276 16454 28304 16594
rect 28264 16448 28316 16454
rect 28264 16390 28316 16396
rect 28264 16108 28316 16114
rect 28264 16050 28316 16056
rect 28276 15366 28304 16050
rect 28264 15360 28316 15366
rect 28264 15302 28316 15308
rect 28276 15162 28304 15302
rect 28264 15156 28316 15162
rect 28264 15098 28316 15104
rect 28264 13320 28316 13326
rect 28264 13262 28316 13268
rect 28276 12714 28304 13262
rect 28264 12708 28316 12714
rect 28264 12650 28316 12656
rect 28172 12640 28224 12646
rect 28172 12582 28224 12588
rect 28170 12472 28226 12481
rect 28368 12442 28396 17206
rect 28460 16658 28488 20742
rect 28552 17066 28580 21830
rect 28644 21554 28672 21898
rect 28632 21548 28684 21554
rect 28632 21490 28684 21496
rect 28816 21480 28868 21486
rect 28816 21422 28868 21428
rect 28724 21344 28776 21350
rect 28724 21286 28776 21292
rect 28736 21146 28764 21286
rect 28724 21140 28776 21146
rect 28724 21082 28776 21088
rect 28632 18692 28684 18698
rect 28632 18634 28684 18640
rect 28644 17882 28672 18634
rect 28632 17876 28684 17882
rect 28632 17818 28684 17824
rect 28736 17320 28764 21082
rect 28828 18426 28856 21422
rect 28908 20800 28960 20806
rect 28908 20742 28960 20748
rect 28816 18420 28868 18426
rect 28816 18362 28868 18368
rect 28828 18086 28856 18362
rect 28920 18358 28948 20742
rect 28908 18352 28960 18358
rect 28908 18294 28960 18300
rect 28816 18080 28868 18086
rect 28816 18022 28868 18028
rect 28906 17912 28962 17921
rect 28906 17847 28962 17856
rect 28644 17292 28764 17320
rect 28540 17060 28592 17066
rect 28540 17002 28592 17008
rect 28644 16794 28672 17292
rect 28920 17270 28948 17847
rect 28908 17264 28960 17270
rect 28908 17206 28960 17212
rect 29090 17232 29146 17241
rect 28724 17196 28776 17202
rect 28724 17138 28776 17144
rect 28816 17196 28868 17202
rect 29090 17167 29146 17176
rect 28816 17138 28868 17144
rect 28736 17105 28764 17138
rect 28722 17096 28778 17105
rect 28722 17031 28778 17040
rect 28632 16788 28684 16794
rect 28632 16730 28684 16736
rect 28448 16652 28500 16658
rect 28500 16612 28580 16640
rect 28448 16594 28500 16600
rect 28446 15736 28502 15745
rect 28446 15671 28502 15680
rect 28460 15638 28488 15671
rect 28448 15632 28500 15638
rect 28448 15574 28500 15580
rect 28446 15464 28502 15473
rect 28446 15399 28502 15408
rect 28170 12407 28226 12416
rect 28356 12436 28408 12442
rect 28184 11121 28212 12407
rect 28356 12378 28408 12384
rect 28368 12288 28396 12378
rect 28276 12260 28396 12288
rect 28170 11112 28226 11121
rect 28170 11047 28226 11056
rect 28172 10600 28224 10606
rect 28172 10542 28224 10548
rect 28184 10266 28212 10542
rect 28172 10260 28224 10266
rect 28172 10202 28224 10208
rect 28172 9716 28224 9722
rect 28172 9658 28224 9664
rect 28184 9110 28212 9658
rect 28172 9104 28224 9110
rect 28172 9046 28224 9052
rect 28170 8528 28226 8537
rect 28170 8463 28226 8472
rect 28184 7478 28212 8463
rect 28276 7886 28304 12260
rect 28460 12186 28488 15399
rect 28552 12986 28580 16612
rect 28724 16448 28776 16454
rect 28724 16390 28776 16396
rect 28736 15570 28764 16390
rect 28724 15564 28776 15570
rect 28724 15506 28776 15512
rect 28632 15020 28684 15026
rect 28632 14962 28684 14968
rect 28644 13802 28672 14962
rect 28828 14770 28856 17138
rect 29104 17066 29132 17167
rect 29092 17060 29144 17066
rect 29092 17002 29144 17008
rect 28908 16584 28960 16590
rect 28908 16526 28960 16532
rect 28920 16250 28948 16526
rect 29092 16448 29144 16454
rect 29092 16390 29144 16396
rect 28908 16244 28960 16250
rect 28908 16186 28960 16192
rect 28908 15564 28960 15570
rect 28908 15506 28960 15512
rect 28920 15450 28948 15506
rect 28920 15422 29040 15450
rect 29104 15434 29132 16390
rect 28908 15156 28960 15162
rect 28908 15098 28960 15104
rect 28920 14822 28948 15098
rect 28736 14742 28856 14770
rect 28908 14816 28960 14822
rect 28908 14758 28960 14764
rect 28632 13796 28684 13802
rect 28632 13738 28684 13744
rect 28632 13252 28684 13258
rect 28632 13194 28684 13200
rect 28540 12980 28592 12986
rect 28540 12922 28592 12928
rect 28644 12918 28672 13194
rect 28632 12912 28684 12918
rect 28632 12854 28684 12860
rect 28540 12640 28592 12646
rect 28540 12582 28592 12588
rect 28368 12158 28488 12186
rect 28368 12073 28396 12158
rect 28448 12096 28500 12102
rect 28354 12064 28410 12073
rect 28448 12038 28500 12044
rect 28354 11999 28410 12008
rect 28368 10538 28396 11999
rect 28460 10810 28488 12038
rect 28448 10804 28500 10810
rect 28448 10746 28500 10752
rect 28460 10674 28488 10746
rect 28448 10668 28500 10674
rect 28448 10610 28500 10616
rect 28356 10532 28408 10538
rect 28356 10474 28408 10480
rect 28552 9976 28580 12582
rect 28460 9948 28580 9976
rect 28460 9722 28488 9948
rect 28538 9888 28594 9897
rect 28538 9823 28594 9832
rect 28448 9716 28500 9722
rect 28448 9658 28500 9664
rect 28356 9648 28408 9654
rect 28356 9590 28408 9596
rect 28446 9616 28502 9625
rect 28368 8634 28396 9590
rect 28446 9551 28448 9560
rect 28500 9551 28502 9560
rect 28448 9522 28500 9528
rect 28448 8900 28500 8906
rect 28448 8842 28500 8848
rect 28356 8628 28408 8634
rect 28356 8570 28408 8576
rect 28264 7880 28316 7886
rect 28264 7822 28316 7828
rect 28172 7472 28224 7478
rect 28172 7414 28224 7420
rect 28276 7274 28304 7822
rect 28264 7268 28316 7274
rect 28264 7210 28316 7216
rect 28080 6860 28132 6866
rect 28080 6802 28132 6808
rect 27988 6792 28040 6798
rect 27988 6734 28040 6740
rect 28172 6792 28224 6798
rect 28172 6734 28224 6740
rect 28000 5386 28028 6734
rect 28184 6361 28212 6734
rect 28264 6452 28316 6458
rect 28264 6394 28316 6400
rect 28170 6352 28226 6361
rect 28170 6287 28226 6296
rect 28000 5358 28120 5386
rect 27988 5296 28040 5302
rect 27988 5238 28040 5244
rect 28000 4282 28028 5238
rect 28092 5166 28120 5358
rect 28080 5160 28132 5166
rect 28080 5102 28132 5108
rect 28080 5024 28132 5030
rect 28080 4966 28132 4972
rect 27988 4276 28040 4282
rect 27988 4218 28040 4224
rect 28092 4214 28120 4966
rect 28080 4208 28132 4214
rect 28080 4150 28132 4156
rect 28172 4208 28224 4214
rect 28172 4150 28224 4156
rect 28078 3632 28134 3641
rect 28078 3567 28134 3576
rect 28092 3398 28120 3567
rect 28080 3392 28132 3398
rect 28080 3334 28132 3340
rect 28092 3097 28120 3334
rect 28078 3088 28134 3097
rect 28078 3023 28134 3032
rect 28184 2922 28212 4150
rect 28276 3670 28304 6394
rect 28460 5302 28488 8842
rect 28552 8430 28580 9823
rect 28540 8424 28592 8430
rect 28540 8366 28592 8372
rect 28644 7410 28672 12854
rect 28736 10033 28764 14742
rect 29012 14634 29040 15422
rect 29092 15428 29144 15434
rect 29092 15370 29144 15376
rect 29092 14816 29144 14822
rect 29092 14758 29144 14764
rect 28920 14606 29040 14634
rect 28920 12238 28948 14606
rect 29104 14482 29132 14758
rect 29092 14476 29144 14482
rect 29092 14418 29144 14424
rect 28998 13968 29054 13977
rect 28998 13903 29054 13912
rect 29012 13802 29040 13903
rect 29000 13796 29052 13802
rect 29000 13738 29052 13744
rect 29092 13320 29144 13326
rect 29092 13262 29144 13268
rect 29104 12306 29132 13262
rect 29092 12300 29144 12306
rect 29092 12242 29144 12248
rect 28908 12232 28960 12238
rect 28908 12174 28960 12180
rect 29196 12170 29224 32370
rect 29276 28620 29328 28626
rect 29276 28562 29328 28568
rect 29288 17134 29316 28562
rect 29644 26308 29696 26314
rect 29644 26250 29696 26256
rect 29656 23322 29684 26250
rect 29644 23316 29696 23322
rect 29644 23258 29696 23264
rect 29460 18828 29512 18834
rect 29460 18770 29512 18776
rect 29368 17264 29420 17270
rect 29368 17206 29420 17212
rect 29276 17128 29328 17134
rect 29276 17070 29328 17076
rect 29276 16176 29328 16182
rect 29276 16118 29328 16124
rect 29288 15434 29316 16118
rect 29276 15428 29328 15434
rect 29276 15370 29328 15376
rect 29276 15088 29328 15094
rect 29276 15030 29328 15036
rect 29288 14618 29316 15030
rect 29276 14612 29328 14618
rect 29276 14554 29328 14560
rect 29276 14408 29328 14414
rect 29276 14350 29328 14356
rect 29288 14074 29316 14350
rect 29276 14068 29328 14074
rect 29276 14010 29328 14016
rect 29380 13954 29408 17206
rect 29472 16182 29500 18770
rect 29552 18284 29604 18290
rect 29552 18226 29604 18232
rect 29564 17921 29592 18226
rect 29550 17912 29606 17921
rect 29550 17847 29606 17856
rect 29656 17270 29684 23258
rect 29736 20936 29788 20942
rect 29736 20878 29788 20884
rect 29748 20262 29776 20878
rect 29736 20256 29788 20262
rect 29736 20198 29788 20204
rect 29748 19854 29776 20198
rect 29736 19848 29788 19854
rect 29736 19790 29788 19796
rect 29644 17264 29696 17270
rect 29644 17206 29696 17212
rect 29748 17082 29776 19790
rect 29840 18290 29868 50322
rect 31116 27600 31168 27606
rect 31116 27542 31168 27548
rect 30840 24200 30892 24206
rect 30840 24142 30892 24148
rect 30012 21616 30064 21622
rect 30012 21558 30064 21564
rect 30024 19446 30052 21558
rect 30748 21004 30800 21010
rect 30748 20946 30800 20952
rect 30380 20800 30432 20806
rect 30380 20742 30432 20748
rect 30012 19440 30064 19446
rect 30012 19382 30064 19388
rect 30392 19378 30420 20742
rect 30472 19848 30524 19854
rect 30472 19790 30524 19796
rect 30656 19848 30708 19854
rect 30656 19790 30708 19796
rect 30288 19372 30340 19378
rect 30288 19314 30340 19320
rect 30380 19372 30432 19378
rect 30380 19314 30432 19320
rect 30300 18834 30328 19314
rect 30288 18828 30340 18834
rect 30288 18770 30340 18776
rect 30012 18760 30064 18766
rect 30012 18702 30064 18708
rect 29828 18284 29880 18290
rect 29828 18226 29880 18232
rect 29920 18216 29972 18222
rect 29656 17054 29776 17082
rect 29840 18164 29920 18170
rect 29840 18158 29972 18164
rect 29840 18142 29960 18158
rect 29460 16176 29512 16182
rect 29460 16118 29512 16124
rect 29552 16040 29604 16046
rect 29552 15982 29604 15988
rect 29460 15972 29512 15978
rect 29460 15914 29512 15920
rect 29472 15706 29500 15914
rect 29460 15700 29512 15706
rect 29460 15642 29512 15648
rect 29288 13926 29408 13954
rect 29184 12164 29236 12170
rect 29184 12106 29236 12112
rect 29000 11348 29052 11354
rect 29000 11290 29052 11296
rect 29012 11234 29040 11290
rect 29196 11257 29224 12106
rect 28920 11206 29040 11234
rect 29182 11248 29238 11257
rect 28920 11150 28948 11206
rect 29182 11183 29238 11192
rect 28908 11144 28960 11150
rect 28908 11086 28960 11092
rect 29000 11144 29052 11150
rect 29000 11086 29052 11092
rect 29012 10713 29040 11086
rect 29092 10804 29144 10810
rect 29092 10746 29144 10752
rect 28998 10704 29054 10713
rect 28998 10639 29054 10648
rect 29104 10606 29132 10746
rect 29182 10704 29238 10713
rect 29182 10639 29238 10648
rect 29092 10600 29144 10606
rect 29092 10542 29144 10548
rect 29196 10470 29224 10639
rect 29184 10464 29236 10470
rect 29184 10406 29236 10412
rect 28906 10296 28962 10305
rect 28906 10231 28962 10240
rect 28816 10192 28868 10198
rect 28816 10134 28868 10140
rect 28828 10062 28856 10134
rect 28920 10062 28948 10231
rect 28816 10056 28868 10062
rect 28722 10024 28778 10033
rect 28816 9998 28868 10004
rect 28908 10056 28960 10062
rect 28908 9998 28960 10004
rect 28722 9959 28778 9968
rect 28736 9364 28764 9959
rect 28814 9616 28870 9625
rect 29288 9586 29316 13926
rect 29368 13864 29420 13870
rect 29368 13806 29420 13812
rect 28814 9551 28870 9560
rect 29276 9580 29328 9586
rect 28828 9518 28856 9551
rect 29380 9568 29408 13806
rect 29564 13190 29592 15982
rect 29656 14822 29684 17054
rect 29736 16108 29788 16114
rect 29736 16050 29788 16056
rect 29748 15706 29776 16050
rect 29736 15700 29788 15706
rect 29736 15642 29788 15648
rect 29736 15428 29788 15434
rect 29736 15370 29788 15376
rect 29644 14816 29696 14822
rect 29644 14758 29696 14764
rect 29644 14544 29696 14550
rect 29644 14486 29696 14492
rect 29656 13938 29684 14486
rect 29748 14414 29776 15370
rect 29840 15162 29868 18142
rect 30024 18086 30052 18702
rect 30378 18456 30434 18465
rect 30484 18426 30512 19790
rect 30564 19712 30616 19718
rect 30564 19654 30616 19660
rect 30576 18766 30604 19654
rect 30668 19514 30696 19790
rect 30656 19508 30708 19514
rect 30656 19450 30708 19456
rect 30564 18760 30616 18766
rect 30564 18702 30616 18708
rect 30656 18692 30708 18698
rect 30656 18634 30708 18640
rect 30668 18601 30696 18634
rect 30654 18592 30710 18601
rect 30654 18527 30710 18536
rect 30378 18391 30434 18400
rect 30472 18420 30524 18426
rect 30196 18216 30248 18222
rect 30196 18158 30248 18164
rect 29920 18080 29972 18086
rect 29920 18022 29972 18028
rect 30012 18080 30064 18086
rect 30012 18022 30064 18028
rect 29932 17542 29960 18022
rect 29920 17536 29972 17542
rect 29920 17478 29972 17484
rect 29828 15156 29880 15162
rect 29828 15098 29880 15104
rect 29826 15056 29882 15065
rect 29826 14991 29828 15000
rect 29880 14991 29882 15000
rect 29828 14962 29880 14968
rect 29736 14408 29788 14414
rect 29736 14350 29788 14356
rect 29644 13932 29696 13938
rect 29644 13874 29696 13880
rect 29552 13184 29604 13190
rect 29552 13126 29604 13132
rect 29748 12918 29776 14350
rect 29736 12912 29788 12918
rect 29736 12854 29788 12860
rect 29932 12764 29960 17478
rect 30012 17196 30064 17202
rect 30208 17184 30236 18158
rect 30392 17814 30420 18391
rect 30472 18362 30524 18368
rect 30656 17876 30708 17882
rect 30656 17818 30708 17824
rect 30380 17808 30432 17814
rect 30380 17750 30432 17756
rect 30472 17740 30524 17746
rect 30472 17682 30524 17688
rect 30484 17610 30512 17682
rect 30668 17610 30696 17818
rect 30472 17604 30524 17610
rect 30472 17546 30524 17552
rect 30656 17604 30708 17610
rect 30656 17546 30708 17552
rect 30064 17156 30236 17184
rect 30012 17138 30064 17144
rect 30024 16658 30052 17138
rect 30012 16652 30064 16658
rect 30012 16594 30064 16600
rect 30380 16516 30432 16522
rect 30380 16458 30432 16464
rect 30392 16250 30420 16458
rect 30380 16244 30432 16250
rect 30380 16186 30432 16192
rect 30484 16182 30512 17546
rect 30760 17270 30788 20946
rect 30852 17377 30880 24142
rect 31128 20806 31156 27542
rect 31312 23050 31340 60998
rect 32496 60104 32548 60110
rect 32496 60046 32548 60052
rect 32312 59968 32364 59974
rect 32312 59910 32364 59916
rect 31576 59424 31628 59430
rect 31576 59366 31628 59372
rect 31484 57248 31536 57254
rect 31484 57190 31536 57196
rect 31300 23044 31352 23050
rect 31300 22986 31352 22992
rect 31208 22092 31260 22098
rect 31208 22034 31260 22040
rect 31220 21010 31248 22034
rect 31208 21004 31260 21010
rect 31208 20946 31260 20952
rect 31024 20800 31076 20806
rect 31024 20742 31076 20748
rect 31116 20800 31168 20806
rect 31116 20742 31168 20748
rect 31300 20800 31352 20806
rect 31300 20742 31352 20748
rect 31036 19174 31064 20742
rect 31024 19168 31076 19174
rect 31024 19110 31076 19116
rect 30838 17368 30894 17377
rect 30838 17303 30894 17312
rect 30748 17264 30800 17270
rect 30748 17206 30800 17212
rect 30472 16176 30524 16182
rect 30472 16118 30524 16124
rect 30380 16108 30432 16114
rect 30380 16050 30432 16056
rect 30012 15904 30064 15910
rect 30012 15846 30064 15852
rect 30024 15434 30052 15846
rect 30012 15428 30064 15434
rect 30012 15370 30064 15376
rect 30104 15020 30156 15026
rect 30104 14962 30156 14968
rect 30012 14952 30064 14958
rect 30012 14894 30064 14900
rect 30024 13870 30052 14894
rect 30012 13864 30064 13870
rect 30012 13806 30064 13812
rect 29656 12736 29960 12764
rect 29458 10160 29514 10169
rect 29458 10095 29514 10104
rect 29472 9722 29500 10095
rect 29552 9920 29604 9926
rect 29552 9862 29604 9868
rect 29564 9761 29592 9862
rect 29550 9752 29606 9761
rect 29460 9716 29512 9722
rect 29550 9687 29552 9696
rect 29460 9658 29512 9664
rect 29604 9687 29606 9696
rect 29552 9658 29604 9664
rect 29380 9540 29500 9568
rect 29276 9522 29328 9528
rect 28816 9512 28868 9518
rect 28816 9454 28868 9460
rect 29092 9512 29144 9518
rect 29472 9500 29500 9540
rect 29472 9489 29592 9500
rect 29472 9480 29606 9489
rect 29472 9472 29550 9480
rect 29092 9454 29144 9460
rect 29000 9376 29052 9382
rect 28736 9336 28856 9364
rect 28724 8628 28776 8634
rect 28724 8570 28776 8576
rect 28736 7954 28764 8570
rect 28724 7948 28776 7954
rect 28724 7890 28776 7896
rect 28724 7812 28776 7818
rect 28724 7754 28776 7760
rect 28632 7404 28684 7410
rect 28632 7346 28684 7352
rect 28540 6860 28592 6866
rect 28540 6802 28592 6808
rect 28552 5710 28580 6802
rect 28644 6390 28672 7346
rect 28632 6384 28684 6390
rect 28632 6326 28684 6332
rect 28540 5704 28592 5710
rect 28540 5646 28592 5652
rect 28736 5642 28764 7754
rect 28828 5710 28856 9336
rect 29000 9318 29052 9324
rect 29012 8498 29040 9318
rect 29104 8906 29132 9454
rect 29550 9415 29606 9424
rect 29184 9036 29236 9042
rect 29184 8978 29236 8984
rect 29092 8900 29144 8906
rect 29092 8842 29144 8848
rect 29196 8820 29224 8978
rect 29196 8792 29316 8820
rect 29000 8492 29052 8498
rect 29000 8434 29052 8440
rect 29092 8288 29144 8294
rect 29092 8230 29144 8236
rect 29288 8242 29316 8792
rect 29552 8560 29604 8566
rect 29550 8528 29552 8537
rect 29604 8528 29606 8537
rect 29460 8492 29512 8498
rect 29550 8463 29606 8472
rect 29460 8434 29512 8440
rect 29104 7342 29132 8230
rect 29288 8214 29408 8242
rect 29276 7540 29328 7546
rect 29276 7482 29328 7488
rect 29092 7336 29144 7342
rect 29092 7278 29144 7284
rect 29092 6112 29144 6118
rect 29092 6054 29144 6060
rect 28908 5840 28960 5846
rect 28908 5782 28960 5788
rect 28816 5704 28868 5710
rect 28816 5646 28868 5652
rect 28724 5636 28776 5642
rect 28724 5578 28776 5584
rect 28448 5296 28500 5302
rect 28448 5238 28500 5244
rect 28814 5264 28870 5273
rect 28540 5228 28592 5234
rect 28814 5199 28870 5208
rect 28540 5170 28592 5176
rect 28356 4684 28408 4690
rect 28356 4626 28408 4632
rect 28264 3664 28316 3670
rect 28264 3606 28316 3612
rect 28368 2990 28396 4626
rect 28448 4140 28500 4146
rect 28448 4082 28500 4088
rect 28460 3398 28488 4082
rect 28552 3924 28580 5170
rect 28828 5098 28856 5199
rect 28632 5092 28684 5098
rect 28632 5034 28684 5040
rect 28816 5092 28868 5098
rect 28816 5034 28868 5040
rect 28644 4554 28672 5034
rect 28722 4720 28778 4729
rect 28722 4655 28778 4664
rect 28736 4622 28764 4655
rect 28724 4616 28776 4622
rect 28724 4558 28776 4564
rect 28632 4548 28684 4554
rect 28632 4490 28684 4496
rect 28816 4480 28868 4486
rect 28816 4422 28868 4428
rect 28724 3936 28776 3942
rect 28552 3896 28724 3924
rect 28724 3878 28776 3884
rect 28736 3534 28764 3878
rect 28724 3528 28776 3534
rect 28724 3470 28776 3476
rect 28448 3392 28500 3398
rect 28448 3334 28500 3340
rect 28356 2984 28408 2990
rect 28356 2926 28408 2932
rect 28172 2916 28224 2922
rect 28172 2858 28224 2864
rect 28828 2582 28856 4422
rect 28816 2576 28868 2582
rect 27894 2544 27950 2553
rect 28816 2518 28868 2524
rect 27894 2479 27950 2488
rect 27908 2446 27936 2479
rect 28920 2446 28948 5782
rect 29000 4004 29052 4010
rect 29000 3946 29052 3952
rect 29012 3058 29040 3946
rect 29104 3534 29132 6054
rect 29092 3528 29144 3534
rect 29092 3470 29144 3476
rect 29288 3466 29316 7482
rect 29380 3602 29408 8214
rect 29472 7886 29500 8434
rect 29460 7880 29512 7886
rect 29460 7822 29512 7828
rect 29656 6440 29684 12736
rect 29828 12368 29880 12374
rect 29828 12310 29880 12316
rect 29840 11286 29868 12310
rect 29920 12096 29972 12102
rect 29920 12038 29972 12044
rect 29932 11898 29960 12038
rect 29920 11892 29972 11898
rect 29920 11834 29972 11840
rect 29736 11280 29788 11286
rect 29736 11222 29788 11228
rect 29828 11280 29880 11286
rect 29828 11222 29880 11228
rect 29748 10470 29776 11222
rect 30010 10976 30066 10985
rect 30010 10911 30066 10920
rect 29828 10736 29880 10742
rect 29828 10678 29880 10684
rect 29736 10464 29788 10470
rect 29736 10406 29788 10412
rect 29840 9994 29868 10678
rect 29920 10668 29972 10674
rect 29920 10610 29972 10616
rect 29828 9988 29880 9994
rect 29828 9930 29880 9936
rect 29932 9674 29960 10610
rect 30024 10062 30052 10911
rect 30012 10056 30064 10062
rect 30012 9998 30064 10004
rect 30116 9994 30144 14962
rect 30196 14340 30248 14346
rect 30196 14282 30248 14288
rect 30208 12730 30236 14282
rect 30392 12850 30420 16050
rect 30472 15360 30524 15366
rect 30470 15328 30472 15337
rect 30524 15328 30526 15337
rect 30470 15263 30526 15272
rect 30472 15156 30524 15162
rect 30472 15098 30524 15104
rect 30484 15065 30512 15098
rect 30470 15056 30526 15065
rect 30470 14991 30526 15000
rect 30748 14544 30800 14550
rect 30668 14504 30748 14532
rect 30668 13802 30696 14504
rect 30748 14486 30800 14492
rect 30656 13796 30708 13802
rect 30656 13738 30708 13744
rect 30380 12844 30432 12850
rect 30380 12786 30432 12792
rect 30208 12702 30328 12730
rect 30300 11830 30328 12702
rect 30288 11824 30340 11830
rect 30288 11766 30340 11772
rect 30288 11212 30340 11218
rect 30288 11154 30340 11160
rect 30194 10840 30250 10849
rect 30300 10810 30328 11154
rect 30194 10775 30250 10784
rect 30288 10804 30340 10810
rect 30208 10062 30236 10775
rect 30288 10746 30340 10752
rect 30288 10464 30340 10470
rect 30288 10406 30340 10412
rect 30196 10056 30248 10062
rect 30196 9998 30248 10004
rect 30104 9988 30156 9994
rect 30104 9930 30156 9936
rect 30010 9752 30066 9761
rect 30010 9687 30066 9696
rect 29736 9648 29788 9654
rect 29734 9616 29736 9625
rect 29913 9646 29960 9674
rect 29788 9616 29790 9625
rect 29734 9551 29790 9560
rect 29913 9500 29941 9646
rect 29913 9472 29960 9500
rect 29828 9376 29880 9382
rect 29828 9318 29880 9324
rect 29736 9104 29788 9110
rect 29736 9046 29788 9052
rect 29748 8838 29776 9046
rect 29736 8832 29788 8838
rect 29736 8774 29788 8780
rect 29736 8424 29788 8430
rect 29736 8366 29788 8372
rect 29564 6412 29684 6440
rect 29368 3596 29420 3602
rect 29368 3538 29420 3544
rect 29276 3460 29328 3466
rect 29276 3402 29328 3408
rect 29090 3088 29146 3097
rect 29000 3052 29052 3058
rect 29090 3023 29146 3032
rect 29000 2994 29052 3000
rect 29104 2990 29132 3023
rect 29092 2984 29144 2990
rect 29092 2926 29144 2932
rect 29092 2848 29144 2854
rect 29092 2790 29144 2796
rect 27896 2440 27948 2446
rect 27896 2382 27948 2388
rect 28908 2440 28960 2446
rect 28908 2382 28960 2388
rect 28816 2372 28868 2378
rect 28816 2314 28868 2320
rect 27988 2100 28040 2106
rect 27988 2042 28040 2048
rect 28000 800 28028 2042
rect 28540 1556 28592 1562
rect 28540 1498 28592 1504
rect 28264 1420 28316 1426
rect 28264 1362 28316 1368
rect 28276 800 28304 1362
rect 28552 800 28580 1498
rect 28828 800 28856 2314
rect 29104 800 29132 2790
rect 29288 2774 29316 3402
rect 29564 3194 29592 6412
rect 29642 6352 29698 6361
rect 29642 6287 29698 6296
rect 29656 5914 29684 6287
rect 29748 5914 29776 8366
rect 29840 7954 29868 9318
rect 29828 7948 29880 7954
rect 29828 7890 29880 7896
rect 29840 6866 29868 7890
rect 29932 7546 29960 9472
rect 30024 8838 30052 9687
rect 30116 9042 30144 9930
rect 30300 9874 30328 10406
rect 30208 9846 30328 9874
rect 30208 9625 30236 9846
rect 30194 9616 30250 9625
rect 30194 9551 30250 9560
rect 30288 9580 30340 9586
rect 30288 9522 30340 9528
rect 30300 9330 30328 9522
rect 30208 9302 30328 9330
rect 30104 9036 30156 9042
rect 30104 8978 30156 8984
rect 30104 8900 30156 8906
rect 30104 8842 30156 8848
rect 30012 8832 30064 8838
rect 30012 8774 30064 8780
rect 30024 7886 30052 8774
rect 30116 8430 30144 8842
rect 30208 8498 30236 9302
rect 30288 9172 30340 9178
rect 30288 9114 30340 9120
rect 30196 8492 30248 8498
rect 30196 8434 30248 8440
rect 30104 8424 30156 8430
rect 30104 8366 30156 8372
rect 30196 8356 30248 8362
rect 30196 8298 30248 8304
rect 30012 7880 30064 7886
rect 30012 7822 30064 7828
rect 30208 7698 30236 8298
rect 30116 7670 30236 7698
rect 29920 7540 29972 7546
rect 29920 7482 29972 7488
rect 30012 7336 30064 7342
rect 30012 7278 30064 7284
rect 29918 7168 29974 7177
rect 29918 7103 29974 7112
rect 29828 6860 29880 6866
rect 29828 6802 29880 6808
rect 29644 5908 29696 5914
rect 29644 5850 29696 5856
rect 29736 5908 29788 5914
rect 29736 5850 29788 5856
rect 29734 5808 29790 5817
rect 29734 5743 29790 5752
rect 29748 5234 29776 5743
rect 29736 5228 29788 5234
rect 29736 5170 29788 5176
rect 29932 4468 29960 7103
rect 30024 5914 30052 7278
rect 30012 5908 30064 5914
rect 30012 5850 30064 5856
rect 30024 5030 30052 5850
rect 30116 5778 30144 7670
rect 30196 7540 30248 7546
rect 30196 7482 30248 7488
rect 30208 5778 30236 7482
rect 30300 6662 30328 9114
rect 30392 7392 30420 12786
rect 30472 12164 30524 12170
rect 30472 12106 30524 12112
rect 30484 11762 30512 12106
rect 30472 11756 30524 11762
rect 30472 11698 30524 11704
rect 30472 11348 30524 11354
rect 30472 11290 30524 11296
rect 30484 10062 30512 11290
rect 30668 11234 30696 13738
rect 30852 12434 30880 17303
rect 31024 15904 31076 15910
rect 31024 15846 31076 15852
rect 31036 14890 31064 15846
rect 31128 15434 31156 20742
rect 31208 18624 31260 18630
rect 31208 18566 31260 18572
rect 31220 18290 31248 18566
rect 31208 18284 31260 18290
rect 31208 18226 31260 18232
rect 31220 17678 31248 18226
rect 31312 18057 31340 20742
rect 31496 18834 31524 57190
rect 31484 18828 31536 18834
rect 31484 18770 31536 18776
rect 31392 18692 31444 18698
rect 31392 18634 31444 18640
rect 31298 18048 31354 18057
rect 31298 17983 31354 17992
rect 31404 17678 31432 18634
rect 31482 18048 31538 18057
rect 31482 17983 31538 17992
rect 31208 17672 31260 17678
rect 31208 17614 31260 17620
rect 31392 17672 31444 17678
rect 31392 17614 31444 17620
rect 31208 17128 31260 17134
rect 31208 17070 31260 17076
rect 31116 15428 31168 15434
rect 31116 15370 31168 15376
rect 31024 14884 31076 14890
rect 31024 14826 31076 14832
rect 31116 14612 31168 14618
rect 31116 14554 31168 14560
rect 31128 12850 31156 14554
rect 30932 12844 30984 12850
rect 30932 12786 30984 12792
rect 31116 12844 31168 12850
rect 31116 12786 31168 12792
rect 30944 12730 30972 12786
rect 30944 12702 31156 12730
rect 31024 12640 31076 12646
rect 31024 12582 31076 12588
rect 30576 11206 30696 11234
rect 30760 12406 30880 12434
rect 30760 11218 30788 12406
rect 30840 12096 30892 12102
rect 30840 12038 30892 12044
rect 30852 11830 30880 12038
rect 30840 11824 30892 11830
rect 30840 11766 30892 11772
rect 30932 11756 30984 11762
rect 30932 11698 30984 11704
rect 30748 11212 30800 11218
rect 30472 10056 30524 10062
rect 30472 9998 30524 10004
rect 30484 8362 30512 9998
rect 30472 8356 30524 8362
rect 30472 8298 30524 8304
rect 30472 8016 30524 8022
rect 30472 7958 30524 7964
rect 30484 7546 30512 7958
rect 30576 7721 30604 11206
rect 30748 11154 30800 11160
rect 30760 10198 30788 11154
rect 30656 10192 30708 10198
rect 30656 10134 30708 10140
rect 30748 10192 30800 10198
rect 30748 10134 30800 10140
rect 30668 10044 30696 10134
rect 30944 10044 30972 11698
rect 31036 10674 31064 12582
rect 31128 11150 31156 12702
rect 31220 12102 31248 17070
rect 31300 16040 31352 16046
rect 31300 15982 31352 15988
rect 31312 13938 31340 15982
rect 31300 13932 31352 13938
rect 31300 13874 31352 13880
rect 31312 12628 31340 13874
rect 31404 12889 31432 17614
rect 31496 13938 31524 17983
rect 31484 13932 31536 13938
rect 31484 13874 31536 13880
rect 31588 13530 31616 59366
rect 32324 55214 32352 59910
rect 32508 59770 32536 60046
rect 32496 59764 32548 59770
rect 32496 59706 32548 59712
rect 32496 56704 32548 56710
rect 32496 56646 32548 56652
rect 32324 55186 32444 55214
rect 32312 43648 32364 43654
rect 32312 43590 32364 43596
rect 32324 43314 32352 43590
rect 32312 43308 32364 43314
rect 32312 43250 32364 43256
rect 31760 35216 31812 35222
rect 31760 35158 31812 35164
rect 31772 35086 31800 35158
rect 31760 35080 31812 35086
rect 31760 35022 31812 35028
rect 32220 33516 32272 33522
rect 32220 33458 32272 33464
rect 32232 30666 32260 33458
rect 32220 30660 32272 30666
rect 32220 30602 32272 30608
rect 31668 19236 31720 19242
rect 31668 19178 31720 19184
rect 31680 18766 31708 19178
rect 31760 18828 31812 18834
rect 31760 18770 31812 18776
rect 31668 18760 31720 18766
rect 31668 18702 31720 18708
rect 31668 18216 31720 18222
rect 31668 18158 31720 18164
rect 31680 17898 31708 18158
rect 31772 18057 31800 18770
rect 32128 18284 32180 18290
rect 31864 18244 32128 18272
rect 31758 18048 31814 18057
rect 31758 17983 31814 17992
rect 31680 17870 31800 17898
rect 31772 17270 31800 17870
rect 31864 17338 31892 18244
rect 32128 18226 32180 18232
rect 32128 17604 32180 17610
rect 32128 17546 32180 17552
rect 31852 17332 31904 17338
rect 31852 17274 31904 17280
rect 31760 17264 31812 17270
rect 31760 17206 31812 17212
rect 32140 17066 32168 17546
rect 32128 17060 32180 17066
rect 32128 17002 32180 17008
rect 31666 16824 31722 16833
rect 31666 16759 31722 16768
rect 31680 16726 31708 16759
rect 31668 16720 31720 16726
rect 31668 16662 31720 16668
rect 31850 15872 31906 15881
rect 31850 15807 31906 15816
rect 31668 15700 31720 15706
rect 31668 15642 31720 15648
rect 31680 15502 31708 15642
rect 31668 15496 31720 15502
rect 31668 15438 31720 15444
rect 31760 14952 31812 14958
rect 31760 14894 31812 14900
rect 31772 14278 31800 14894
rect 31668 14272 31720 14278
rect 31668 14214 31720 14220
rect 31760 14272 31812 14278
rect 31760 14214 31812 14220
rect 31576 13524 31628 13530
rect 31576 13466 31628 13472
rect 31574 13424 31630 13433
rect 31574 13359 31576 13368
rect 31628 13359 31630 13368
rect 31576 13330 31628 13336
rect 31576 13252 31628 13258
rect 31576 13194 31628 13200
rect 31390 12880 31446 12889
rect 31390 12815 31392 12824
rect 31444 12815 31446 12824
rect 31392 12786 31444 12792
rect 31312 12600 31432 12628
rect 31300 12232 31352 12238
rect 31300 12174 31352 12180
rect 31208 12096 31260 12102
rect 31208 12038 31260 12044
rect 31220 11626 31248 12038
rect 31208 11620 31260 11626
rect 31208 11562 31260 11568
rect 31312 11558 31340 12174
rect 31404 12102 31432 12600
rect 31484 12300 31536 12306
rect 31484 12242 31536 12248
rect 31392 12096 31444 12102
rect 31392 12038 31444 12044
rect 31300 11552 31352 11558
rect 31300 11494 31352 11500
rect 31404 11370 31432 12038
rect 31496 11694 31524 12242
rect 31484 11688 31536 11694
rect 31484 11630 31536 11636
rect 31312 11342 31432 11370
rect 31116 11144 31168 11150
rect 31116 11086 31168 11092
rect 31312 11014 31340 11342
rect 31484 11144 31536 11150
rect 31390 11112 31446 11121
rect 31484 11086 31536 11092
rect 31390 11047 31446 11056
rect 31300 11008 31352 11014
rect 31300 10950 31352 10956
rect 31024 10668 31076 10674
rect 31024 10610 31076 10616
rect 30668 10016 30972 10044
rect 30654 9616 30710 9625
rect 30654 9551 30710 9560
rect 30668 9110 30696 9551
rect 30656 9104 30708 9110
rect 30656 9046 30708 9052
rect 30656 8492 30708 8498
rect 30656 8434 30708 8440
rect 30562 7712 30618 7721
rect 30562 7647 30618 7656
rect 30472 7540 30524 7546
rect 30472 7482 30524 7488
rect 30392 7364 30512 7392
rect 30380 7268 30432 7274
rect 30380 7210 30432 7216
rect 30392 7041 30420 7210
rect 30378 7032 30434 7041
rect 30378 6967 30434 6976
rect 30380 6724 30432 6730
rect 30380 6666 30432 6672
rect 30288 6656 30340 6662
rect 30288 6598 30340 6604
rect 30104 5772 30156 5778
rect 30104 5714 30156 5720
rect 30196 5772 30248 5778
rect 30196 5714 30248 5720
rect 30208 5352 30236 5714
rect 30116 5324 30236 5352
rect 30012 5024 30064 5030
rect 30012 4966 30064 4972
rect 30012 4480 30064 4486
rect 29932 4440 30012 4468
rect 30012 4422 30064 4428
rect 29736 4140 29788 4146
rect 29736 4082 29788 4088
rect 29644 4072 29696 4078
rect 29644 4014 29696 4020
rect 29552 3188 29604 3194
rect 29552 3130 29604 3136
rect 29196 2746 29316 2774
rect 29196 2446 29224 2746
rect 29368 2508 29420 2514
rect 29368 2450 29420 2456
rect 29184 2440 29236 2446
rect 29184 2382 29236 2388
rect 29380 800 29408 2450
rect 29656 800 29684 4014
rect 29748 3670 29776 4082
rect 30116 4010 30144 5324
rect 30194 5264 30250 5273
rect 30194 5199 30250 5208
rect 30208 5098 30236 5199
rect 30196 5092 30248 5098
rect 30196 5034 30248 5040
rect 30104 4004 30156 4010
rect 30104 3946 30156 3952
rect 29736 3664 29788 3670
rect 29736 3606 29788 3612
rect 30116 3602 30144 3946
rect 30392 3913 30420 6666
rect 30484 4214 30512 7364
rect 30564 7200 30616 7206
rect 30564 7142 30616 7148
rect 30576 6458 30604 7142
rect 30564 6452 30616 6458
rect 30564 6394 30616 6400
rect 30564 6316 30616 6322
rect 30564 6258 30616 6264
rect 30576 5234 30604 6258
rect 30564 5228 30616 5234
rect 30564 5170 30616 5176
rect 30564 4616 30616 4622
rect 30668 4604 30696 8434
rect 30616 4576 30696 4604
rect 30564 4558 30616 4564
rect 30472 4208 30524 4214
rect 30472 4150 30524 4156
rect 30378 3904 30434 3913
rect 30378 3839 30434 3848
rect 30104 3596 30156 3602
rect 30104 3538 30156 3544
rect 30196 3460 30248 3466
rect 30196 3402 30248 3408
rect 29920 2372 29972 2378
rect 29920 2314 29972 2320
rect 29932 800 29960 2314
rect 30208 800 30236 3402
rect 30760 3126 30788 10016
rect 31116 9988 31168 9994
rect 31116 9930 31168 9936
rect 31024 9580 31076 9586
rect 31024 9522 31076 9528
rect 31036 9382 31064 9522
rect 31024 9376 31076 9382
rect 31024 9318 31076 9324
rect 31024 8560 31076 8566
rect 31024 8502 31076 8508
rect 30930 8256 30986 8265
rect 30930 8191 30986 8200
rect 30944 8022 30972 8191
rect 30932 8016 30984 8022
rect 30932 7958 30984 7964
rect 31036 7886 31064 8502
rect 31024 7880 31076 7886
rect 31024 7822 31076 7828
rect 31128 7750 31156 9930
rect 31208 9920 31260 9926
rect 31208 9862 31260 9868
rect 31220 8362 31248 9862
rect 31300 9648 31352 9654
rect 31300 9590 31352 9596
rect 31312 8430 31340 9590
rect 31404 9110 31432 11047
rect 31496 11014 31524 11086
rect 31484 11008 31536 11014
rect 31484 10950 31536 10956
rect 31484 10668 31536 10674
rect 31484 10610 31536 10616
rect 31496 10266 31524 10610
rect 31588 10441 31616 13194
rect 31680 10690 31708 14214
rect 31760 14068 31812 14074
rect 31760 14010 31812 14016
rect 31772 11257 31800 14010
rect 31864 13938 31892 15807
rect 32140 15502 32168 17002
rect 32232 16522 32260 30602
rect 32416 26234 32444 55186
rect 32324 26206 32444 26234
rect 32220 16516 32272 16522
rect 32220 16458 32272 16464
rect 32128 15496 32180 15502
rect 32128 15438 32180 15444
rect 31944 15088 31996 15094
rect 31944 15030 31996 15036
rect 31956 13938 31984 15030
rect 32036 15020 32088 15026
rect 32036 14962 32088 14968
rect 32048 14618 32076 14962
rect 32036 14612 32088 14618
rect 32036 14554 32088 14560
rect 32034 14376 32090 14385
rect 32034 14311 32090 14320
rect 32048 14006 32076 14311
rect 32140 14074 32168 15438
rect 32128 14068 32180 14074
rect 32128 14010 32180 14016
rect 32036 14000 32088 14006
rect 32036 13942 32088 13948
rect 31852 13932 31904 13938
rect 31852 13874 31904 13880
rect 31944 13932 31996 13938
rect 31944 13874 31996 13880
rect 32232 13852 32260 16458
rect 32048 13824 32260 13852
rect 31944 12708 31996 12714
rect 31944 12650 31996 12656
rect 31852 12640 31904 12646
rect 31852 12582 31904 12588
rect 31864 12306 31892 12582
rect 31852 12300 31904 12306
rect 31852 12242 31904 12248
rect 31956 12238 31984 12650
rect 31944 12232 31996 12238
rect 31944 12174 31996 12180
rect 31852 11688 31904 11694
rect 31852 11630 31904 11636
rect 31758 11248 31814 11257
rect 31864 11218 31892 11630
rect 31944 11620 31996 11626
rect 31944 11562 31996 11568
rect 31758 11183 31814 11192
rect 31852 11212 31904 11218
rect 31852 11154 31904 11160
rect 31758 10704 31814 10713
rect 31680 10662 31758 10690
rect 31758 10639 31814 10648
rect 31760 10600 31812 10606
rect 31760 10542 31812 10548
rect 31574 10432 31630 10441
rect 31574 10367 31630 10376
rect 31484 10260 31536 10266
rect 31484 10202 31536 10208
rect 31772 9586 31800 10542
rect 31956 9722 31984 11562
rect 32048 10849 32076 13824
rect 32126 13288 32182 13297
rect 32126 13223 32128 13232
rect 32180 13223 32182 13232
rect 32128 13194 32180 13200
rect 32324 12442 32352 26206
rect 32404 24268 32456 24274
rect 32404 24210 32456 24216
rect 32416 23338 32444 24210
rect 32508 23526 32536 56646
rect 32600 46986 32628 60998
rect 33048 60512 33100 60518
rect 33048 60454 33100 60460
rect 33060 60110 33088 60454
rect 32680 60104 32732 60110
rect 32680 60046 32732 60052
rect 33048 60104 33100 60110
rect 33048 60046 33100 60052
rect 32692 59945 32720 60046
rect 32678 59936 32734 59945
rect 32678 59871 32734 59880
rect 32692 59770 32720 59871
rect 32680 59764 32732 59770
rect 32680 59706 32732 59712
rect 33048 59764 33100 59770
rect 33048 59706 33100 59712
rect 32956 59492 33008 59498
rect 32956 59434 33008 59440
rect 32968 56914 32996 59434
rect 32956 56908 33008 56914
rect 32956 56850 33008 56856
rect 33060 56846 33088 59706
rect 33048 56840 33100 56846
rect 33048 56782 33100 56788
rect 32588 46980 32640 46986
rect 32588 46922 32640 46928
rect 33048 43716 33100 43722
rect 33048 43658 33100 43664
rect 32772 43308 32824 43314
rect 32772 43250 32824 43256
rect 32784 43217 32812 43250
rect 32770 43208 32826 43217
rect 32770 43143 32826 43152
rect 32784 42770 32812 43143
rect 32956 43104 33008 43110
rect 32956 43046 33008 43052
rect 32772 42764 32824 42770
rect 32772 42706 32824 42712
rect 32772 42560 32824 42566
rect 32772 42502 32824 42508
rect 32496 23520 32548 23526
rect 32496 23462 32548 23468
rect 32416 23310 32536 23338
rect 32508 22094 32536 23310
rect 32508 22066 32720 22094
rect 32496 21140 32548 21146
rect 32496 21082 32548 21088
rect 32508 20806 32536 21082
rect 32496 20800 32548 20806
rect 32496 20742 32548 20748
rect 32496 20324 32548 20330
rect 32496 20266 32548 20272
rect 32508 19378 32536 20266
rect 32496 19372 32548 19378
rect 32496 19314 32548 19320
rect 32402 17776 32458 17785
rect 32402 17711 32404 17720
rect 32456 17711 32458 17720
rect 32404 17682 32456 17688
rect 32586 17640 32642 17649
rect 32586 17575 32642 17584
rect 32600 17270 32628 17575
rect 32588 17264 32640 17270
rect 32588 17206 32640 17212
rect 32404 17128 32456 17134
rect 32404 17070 32456 17076
rect 32416 16114 32444 17070
rect 32496 16516 32548 16522
rect 32496 16458 32548 16464
rect 32404 16108 32456 16114
rect 32404 16050 32456 16056
rect 32416 16017 32444 16050
rect 32402 16008 32458 16017
rect 32402 15943 32458 15952
rect 32404 13864 32456 13870
rect 32404 13806 32456 13812
rect 32312 12436 32364 12442
rect 32312 12378 32364 12384
rect 32310 12064 32366 12073
rect 32310 11999 32366 12008
rect 32324 11762 32352 11999
rect 32312 11756 32364 11762
rect 32312 11698 32364 11704
rect 32416 11626 32444 13806
rect 32508 13326 32536 16458
rect 32692 16114 32720 22066
rect 32588 16108 32640 16114
rect 32588 16050 32640 16056
rect 32680 16108 32732 16114
rect 32680 16050 32732 16056
rect 32600 15881 32628 16050
rect 32586 15872 32642 15881
rect 32586 15807 32642 15816
rect 32588 15156 32640 15162
rect 32588 15098 32640 15104
rect 32680 15156 32732 15162
rect 32680 15098 32732 15104
rect 32600 14822 32628 15098
rect 32588 14816 32640 14822
rect 32588 14758 32640 14764
rect 32692 14414 32720 15098
rect 32680 14408 32732 14414
rect 32680 14350 32732 14356
rect 32680 13932 32732 13938
rect 32680 13874 32732 13880
rect 32496 13320 32548 13326
rect 32496 13262 32548 13268
rect 32588 13252 32640 13258
rect 32588 13194 32640 13200
rect 32496 13184 32548 13190
rect 32496 13126 32548 13132
rect 32508 12306 32536 13126
rect 32600 12322 32628 13194
rect 32692 13161 32720 13874
rect 32678 13152 32734 13161
rect 32678 13087 32734 13096
rect 32680 12844 32732 12850
rect 32680 12786 32732 12792
rect 32692 12442 32720 12786
rect 32680 12436 32732 12442
rect 32680 12378 32732 12384
rect 32496 12300 32548 12306
rect 32600 12294 32720 12322
rect 32496 12242 32548 12248
rect 32588 12232 32640 12238
rect 32588 12174 32640 12180
rect 32404 11620 32456 11626
rect 32404 11562 32456 11568
rect 32128 11552 32180 11558
rect 32128 11494 32180 11500
rect 32220 11552 32272 11558
rect 32220 11494 32272 11500
rect 32140 11150 32168 11494
rect 32128 11144 32180 11150
rect 32128 11086 32180 11092
rect 32034 10840 32090 10849
rect 32034 10775 32090 10784
rect 32128 10804 32180 10810
rect 32128 10746 32180 10752
rect 32140 10713 32168 10746
rect 32126 10704 32182 10713
rect 32126 10639 32182 10648
rect 32232 10266 32260 11494
rect 32404 11280 32456 11286
rect 32404 11222 32456 11228
rect 32312 11144 32364 11150
rect 32312 11086 32364 11092
rect 32220 10260 32272 10266
rect 32220 10202 32272 10208
rect 32036 10124 32088 10130
rect 32036 10066 32088 10072
rect 31944 9716 31996 9722
rect 31944 9658 31996 9664
rect 31760 9580 31812 9586
rect 31760 9522 31812 9528
rect 31668 9444 31720 9450
rect 31668 9386 31720 9392
rect 31576 9376 31628 9382
rect 31576 9318 31628 9324
rect 31392 9104 31444 9110
rect 31392 9046 31444 9052
rect 31588 8974 31616 9318
rect 31484 8968 31536 8974
rect 31484 8910 31536 8916
rect 31576 8968 31628 8974
rect 31576 8910 31628 8916
rect 31392 8832 31444 8838
rect 31392 8774 31444 8780
rect 31300 8424 31352 8430
rect 31298 8392 31300 8401
rect 31352 8392 31354 8401
rect 31208 8356 31260 8362
rect 31298 8327 31354 8336
rect 31208 8298 31260 8304
rect 31220 7818 31248 8298
rect 31300 8288 31352 8294
rect 31300 8230 31352 8236
rect 31312 8022 31340 8230
rect 31300 8016 31352 8022
rect 31300 7958 31352 7964
rect 31208 7812 31260 7818
rect 31208 7754 31260 7760
rect 31116 7744 31168 7750
rect 31116 7686 31168 7692
rect 31206 7712 31262 7721
rect 31206 7647 31262 7656
rect 30838 7032 30894 7041
rect 30838 6967 30894 6976
rect 30852 6934 30880 6967
rect 30840 6928 30892 6934
rect 30840 6870 30892 6876
rect 31024 6860 31076 6866
rect 31024 6802 31076 6808
rect 30838 5400 30894 5409
rect 30838 5335 30894 5344
rect 30852 5302 30880 5335
rect 30840 5296 30892 5302
rect 30840 5238 30892 5244
rect 31036 5234 31064 6802
rect 31116 5364 31168 5370
rect 31116 5306 31168 5312
rect 31024 5228 31076 5234
rect 31024 5170 31076 5176
rect 31128 4554 31156 5306
rect 31116 4548 31168 4554
rect 31116 4490 31168 4496
rect 30932 4208 30984 4214
rect 30932 4150 30984 4156
rect 30840 3936 30892 3942
rect 30840 3878 30892 3884
rect 30748 3120 30800 3126
rect 30748 3062 30800 3068
rect 30852 3058 30880 3878
rect 30840 3052 30892 3058
rect 30840 2994 30892 3000
rect 30748 2984 30800 2990
rect 30748 2926 30800 2932
rect 30472 2372 30524 2378
rect 30472 2314 30524 2320
rect 30484 800 30512 2314
rect 30760 800 30788 2926
rect 30944 2446 30972 4150
rect 31220 4146 31248 7647
rect 31404 5370 31432 8774
rect 31496 7585 31524 8910
rect 31680 8838 31708 9386
rect 31850 9208 31906 9217
rect 31850 9143 31906 9152
rect 31668 8832 31720 8838
rect 31574 8800 31630 8809
rect 31668 8774 31720 8780
rect 31574 8735 31630 8744
rect 31588 8634 31616 8735
rect 31666 8664 31722 8673
rect 31576 8628 31628 8634
rect 31666 8599 31722 8608
rect 31576 8570 31628 8576
rect 31680 8401 31708 8599
rect 31760 8424 31812 8430
rect 31666 8392 31722 8401
rect 31760 8366 31812 8372
rect 31666 8327 31722 8336
rect 31668 8016 31720 8022
rect 31668 7958 31720 7964
rect 31482 7576 31538 7585
rect 31482 7511 31538 7520
rect 31576 7540 31628 7546
rect 31576 7482 31628 7488
rect 31588 6934 31616 7482
rect 31576 6928 31628 6934
rect 31576 6870 31628 6876
rect 31680 6866 31708 7958
rect 31668 6860 31720 6866
rect 31668 6802 31720 6808
rect 31484 6792 31536 6798
rect 31482 6760 31484 6769
rect 31576 6792 31628 6798
rect 31536 6760 31538 6769
rect 31576 6734 31628 6740
rect 31482 6695 31538 6704
rect 31588 5574 31616 6734
rect 31576 5568 31628 5574
rect 31576 5510 31628 5516
rect 31392 5364 31444 5370
rect 31392 5306 31444 5312
rect 31298 5264 31354 5273
rect 31298 5199 31300 5208
rect 31352 5199 31354 5208
rect 31300 5170 31352 5176
rect 31772 4826 31800 8366
rect 31864 8022 31892 9143
rect 31944 8900 31996 8906
rect 31944 8842 31996 8848
rect 31852 8016 31904 8022
rect 31852 7958 31904 7964
rect 31852 7744 31904 7750
rect 31852 7686 31904 7692
rect 31864 7002 31892 7686
rect 31852 6996 31904 7002
rect 31852 6938 31904 6944
rect 31956 5642 31984 8842
rect 31944 5636 31996 5642
rect 31944 5578 31996 5584
rect 31852 5568 31904 5574
rect 31852 5510 31904 5516
rect 31760 4820 31812 4826
rect 31760 4762 31812 4768
rect 31864 4758 31892 5510
rect 31852 4752 31904 4758
rect 31852 4694 31904 4700
rect 31942 4720 31998 4729
rect 32048 4690 32076 10066
rect 32128 10056 32180 10062
rect 32128 9998 32180 10004
rect 32218 10024 32274 10033
rect 32140 9722 32168 9998
rect 32218 9959 32274 9968
rect 32232 9926 32260 9959
rect 32220 9920 32272 9926
rect 32220 9862 32272 9868
rect 32128 9716 32180 9722
rect 32128 9658 32180 9664
rect 32232 9058 32260 9862
rect 32324 9081 32352 11086
rect 32416 10062 32444 11222
rect 32496 11212 32548 11218
rect 32496 11154 32548 11160
rect 32404 10056 32456 10062
rect 32404 9998 32456 10004
rect 32508 9178 32536 11154
rect 32600 10606 32628 12174
rect 32588 10600 32640 10606
rect 32588 10542 32640 10548
rect 32692 9722 32720 12294
rect 32784 11694 32812 42502
rect 32864 17604 32916 17610
rect 32864 17546 32916 17552
rect 32876 17134 32904 17546
rect 32864 17128 32916 17134
rect 32864 17070 32916 17076
rect 32876 14521 32904 17070
rect 32862 14512 32918 14521
rect 32862 14447 32918 14456
rect 32864 13184 32916 13190
rect 32864 13126 32916 13132
rect 32876 12782 32904 13126
rect 32968 12850 32996 43046
rect 33060 42702 33088 43658
rect 33152 42702 33180 61066
rect 33428 61062 33456 61678
rect 33520 61198 33548 63294
rect 33966 63294 34376 63322
rect 33966 63200 34022 63294
rect 33508 61192 33560 61198
rect 33508 61134 33560 61140
rect 34348 61112 34376 63294
rect 34702 63200 34758 64000
rect 35438 63322 35494 64000
rect 36174 63322 36230 64000
rect 36910 63322 36966 64000
rect 35438 63294 35848 63322
rect 35438 63200 35494 63294
rect 34716 61198 34744 63200
rect 34934 61500 35242 61509
rect 34934 61498 34940 61500
rect 34996 61498 35020 61500
rect 35076 61498 35100 61500
rect 35156 61498 35180 61500
rect 35236 61498 35242 61500
rect 34996 61446 34998 61498
rect 35178 61446 35180 61498
rect 34934 61444 34940 61446
rect 34996 61444 35020 61446
rect 35076 61444 35100 61446
rect 35156 61444 35180 61446
rect 35236 61444 35242 61446
rect 34934 61435 35242 61444
rect 35820 61282 35848 63294
rect 36174 63294 36400 63322
rect 36174 63200 36230 63294
rect 35820 61266 35940 61282
rect 35820 61260 35952 61266
rect 35820 61254 35900 61260
rect 35900 61202 35952 61208
rect 34704 61192 34756 61198
rect 34704 61134 34756 61140
rect 34520 61124 34572 61130
rect 34348 61084 34520 61112
rect 34520 61066 34572 61072
rect 35900 61124 35952 61130
rect 35900 61066 35952 61072
rect 33416 61056 33468 61062
rect 33416 60998 33468 61004
rect 35072 61056 35124 61062
rect 35072 60998 35124 61004
rect 35084 60518 35112 60998
rect 35072 60512 35124 60518
rect 35072 60454 35124 60460
rect 35716 60512 35768 60518
rect 35716 60454 35768 60460
rect 34934 60412 35242 60421
rect 34934 60410 34940 60412
rect 34996 60410 35020 60412
rect 35076 60410 35100 60412
rect 35156 60410 35180 60412
rect 35236 60410 35242 60412
rect 34996 60358 34998 60410
rect 35178 60358 35180 60410
rect 34934 60356 34940 60358
rect 34996 60356 35020 60358
rect 35076 60356 35100 60358
rect 35156 60356 35180 60358
rect 35236 60356 35242 60358
rect 34934 60347 35242 60356
rect 34520 60104 34572 60110
rect 34520 60046 34572 60052
rect 34532 57458 34560 60046
rect 34934 59324 35242 59333
rect 34934 59322 34940 59324
rect 34996 59322 35020 59324
rect 35076 59322 35100 59324
rect 35156 59322 35180 59324
rect 35236 59322 35242 59324
rect 34996 59270 34998 59322
rect 35178 59270 35180 59322
rect 34934 59268 34940 59270
rect 34996 59268 35020 59270
rect 35076 59268 35100 59270
rect 35156 59268 35180 59270
rect 35236 59268 35242 59270
rect 34934 59259 35242 59268
rect 34934 58236 35242 58245
rect 34934 58234 34940 58236
rect 34996 58234 35020 58236
rect 35076 58234 35100 58236
rect 35156 58234 35180 58236
rect 35236 58234 35242 58236
rect 34996 58182 34998 58234
rect 35178 58182 35180 58234
rect 34934 58180 34940 58182
rect 34996 58180 35020 58182
rect 35076 58180 35100 58182
rect 35156 58180 35180 58182
rect 35236 58180 35242 58182
rect 34934 58171 35242 58180
rect 35348 58132 35400 58138
rect 35348 58074 35400 58080
rect 34704 57860 34756 57866
rect 34704 57802 34756 57808
rect 34612 57520 34664 57526
rect 34612 57462 34664 57468
rect 34520 57452 34572 57458
rect 34520 57394 34572 57400
rect 34060 44532 34112 44538
rect 34060 44474 34112 44480
rect 34072 44402 34100 44474
rect 34060 44396 34112 44402
rect 34060 44338 34112 44344
rect 34152 44396 34204 44402
rect 34152 44338 34204 44344
rect 33692 43648 33744 43654
rect 33692 43590 33744 43596
rect 33704 43450 33732 43590
rect 33232 43444 33284 43450
rect 33232 43386 33284 43392
rect 33692 43444 33744 43450
rect 33692 43386 33744 43392
rect 33048 42696 33100 42702
rect 33048 42638 33100 42644
rect 33140 42696 33192 42702
rect 33140 42638 33192 42644
rect 33060 35834 33088 42638
rect 33244 36242 33272 43386
rect 33704 42702 33732 43386
rect 33692 42696 33744 42702
rect 33692 42638 33744 42644
rect 33876 42696 33928 42702
rect 33876 42638 33928 42644
rect 33888 42362 33916 42638
rect 33876 42356 33928 42362
rect 33876 42298 33928 42304
rect 33784 39296 33836 39302
rect 33784 39238 33836 39244
rect 33232 36236 33284 36242
rect 33232 36178 33284 36184
rect 33048 35828 33100 35834
rect 33048 35770 33100 35776
rect 33060 35494 33088 35770
rect 33048 35488 33100 35494
rect 33048 35430 33100 35436
rect 33140 29708 33192 29714
rect 33140 29650 33192 29656
rect 33152 26994 33180 29650
rect 33796 27606 33824 39238
rect 34164 33658 34192 44338
rect 34624 44266 34652 57462
rect 34612 44260 34664 44266
rect 34612 44202 34664 44208
rect 34244 43920 34296 43926
rect 34244 43862 34296 43868
rect 34256 42702 34284 43862
rect 34244 42696 34296 42702
rect 34244 42638 34296 42644
rect 34152 33652 34204 33658
rect 34152 33594 34204 33600
rect 34716 30802 34744 57802
rect 34934 57148 35242 57157
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57083 35242 57092
rect 34934 56060 35242 56069
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55995 35242 56004
rect 35360 55690 35388 58074
rect 35624 57928 35676 57934
rect 35624 57870 35676 57876
rect 35636 57390 35664 57870
rect 35728 57798 35756 60454
rect 35716 57792 35768 57798
rect 35716 57734 35768 57740
rect 35624 57384 35676 57390
rect 35624 57326 35676 57332
rect 35348 55684 35400 55690
rect 35348 55626 35400 55632
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 35360 45558 35388 55626
rect 35808 47592 35860 47598
rect 35808 47534 35860 47540
rect 35348 45552 35400 45558
rect 35348 45494 35400 45500
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 35360 43654 35388 45494
rect 35348 43648 35400 43654
rect 35348 43590 35400 43596
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 34796 42696 34848 42702
rect 34796 42638 34848 42644
rect 34704 30796 34756 30802
rect 34704 30738 34756 30744
rect 34060 28484 34112 28490
rect 34060 28426 34112 28432
rect 33784 27600 33836 27606
rect 33784 27542 33836 27548
rect 33140 26988 33192 26994
rect 33140 26930 33192 26936
rect 33140 23520 33192 23526
rect 33140 23462 33192 23468
rect 33152 22094 33180 23462
rect 33152 22066 33364 22094
rect 33140 19372 33192 19378
rect 33140 19314 33192 19320
rect 33048 18624 33100 18630
rect 33048 18566 33100 18572
rect 33060 17746 33088 18566
rect 33152 18465 33180 19314
rect 33138 18456 33194 18465
rect 33138 18391 33194 18400
rect 33048 17740 33100 17746
rect 33048 17682 33100 17688
rect 33048 17604 33100 17610
rect 33048 17546 33100 17552
rect 33060 17241 33088 17546
rect 33232 17536 33284 17542
rect 33232 17478 33284 17484
rect 33046 17232 33102 17241
rect 33046 17167 33102 17176
rect 33140 17128 33192 17134
rect 33140 17070 33192 17076
rect 33152 16794 33180 17070
rect 33140 16788 33192 16794
rect 33140 16730 33192 16736
rect 33048 16584 33100 16590
rect 33048 16526 33100 16532
rect 33060 16114 33088 16526
rect 33048 16108 33100 16114
rect 33048 16050 33100 16056
rect 33152 14940 33180 16730
rect 33244 16590 33272 17478
rect 33232 16584 33284 16590
rect 33232 16526 33284 16532
rect 33232 14952 33284 14958
rect 33152 14912 33232 14940
rect 33232 14894 33284 14900
rect 33048 14408 33100 14414
rect 33048 14350 33100 14356
rect 33060 14074 33088 14350
rect 33048 14068 33100 14074
rect 33048 14010 33100 14016
rect 33244 12918 33272 14894
rect 33232 12912 33284 12918
rect 33232 12854 33284 12860
rect 32956 12844 33008 12850
rect 32956 12786 33008 12792
rect 32864 12776 32916 12782
rect 33336 12730 33364 22066
rect 33692 20256 33744 20262
rect 33692 20198 33744 20204
rect 33704 19446 33732 20198
rect 33784 19508 33836 19514
rect 33784 19450 33836 19456
rect 33692 19440 33744 19446
rect 33692 19382 33744 19388
rect 33692 19236 33744 19242
rect 33692 19178 33744 19184
rect 33704 18902 33732 19178
rect 33692 18896 33744 18902
rect 33692 18838 33744 18844
rect 33692 18692 33744 18698
rect 33692 18634 33744 18640
rect 33704 17898 33732 18634
rect 33796 18086 33824 19450
rect 33876 18284 33928 18290
rect 33876 18226 33928 18232
rect 33784 18080 33836 18086
rect 33784 18022 33836 18028
rect 33782 17912 33838 17921
rect 33704 17870 33782 17898
rect 33782 17847 33838 17856
rect 33796 17746 33824 17847
rect 33784 17740 33836 17746
rect 33784 17682 33836 17688
rect 33888 17610 33916 18226
rect 33968 18148 34020 18154
rect 33968 18090 34020 18096
rect 33876 17604 33928 17610
rect 33876 17546 33928 17552
rect 33692 17536 33744 17542
rect 33692 17478 33744 17484
rect 33704 17338 33732 17478
rect 33692 17332 33744 17338
rect 33692 17274 33744 17280
rect 33980 17202 34008 18090
rect 33968 17196 34020 17202
rect 33968 17138 34020 17144
rect 33598 16824 33654 16833
rect 33598 16759 33600 16768
rect 33652 16759 33654 16768
rect 33600 16730 33652 16736
rect 33508 14884 33560 14890
rect 33508 14826 33560 14832
rect 33416 14476 33468 14482
rect 33416 14418 33468 14424
rect 33428 14006 33456 14418
rect 33520 14278 33548 14826
rect 33508 14272 33560 14278
rect 33508 14214 33560 14220
rect 33600 14272 33652 14278
rect 33600 14214 33652 14220
rect 33416 14000 33468 14006
rect 33416 13942 33468 13948
rect 32864 12718 32916 12724
rect 33152 12702 33364 12730
rect 33416 12776 33468 12782
rect 33416 12718 33468 12724
rect 32956 12436 33008 12442
rect 32956 12378 33008 12384
rect 32968 12322 32996 12378
rect 32876 12294 32996 12322
rect 32876 11830 32904 12294
rect 32956 12232 33008 12238
rect 32956 12174 33008 12180
rect 32864 11824 32916 11830
rect 32864 11766 32916 11772
rect 32772 11688 32824 11694
rect 32772 11630 32824 11636
rect 32772 11008 32824 11014
rect 32772 10950 32824 10956
rect 32680 9716 32732 9722
rect 32680 9658 32732 9664
rect 32680 9580 32732 9586
rect 32680 9522 32732 9528
rect 32588 9376 32640 9382
rect 32588 9318 32640 9324
rect 32496 9172 32548 9178
rect 32496 9114 32548 9120
rect 32600 9110 32628 9318
rect 32588 9104 32640 9110
rect 32140 9030 32260 9058
rect 32310 9072 32366 9081
rect 32140 6322 32168 9030
rect 32588 9046 32640 9052
rect 32310 9007 32366 9016
rect 32220 8968 32272 8974
rect 32220 8910 32272 8916
rect 32232 7886 32260 8910
rect 32220 7880 32272 7886
rect 32220 7822 32272 7828
rect 32232 7274 32260 7822
rect 32220 7268 32272 7274
rect 32220 7210 32272 7216
rect 32128 6316 32180 6322
rect 32128 6258 32180 6264
rect 32218 5672 32274 5681
rect 32218 5607 32274 5616
rect 31942 4655 31944 4664
rect 31996 4655 31998 4664
rect 32036 4684 32088 4690
rect 31944 4626 31996 4632
rect 32036 4626 32088 4632
rect 32232 4622 32260 5607
rect 32220 4616 32272 4622
rect 31482 4584 31538 4593
rect 32220 4558 32272 4564
rect 31482 4519 31538 4528
rect 31496 4146 31524 4519
rect 31576 4480 31628 4486
rect 32220 4480 32272 4486
rect 31576 4422 31628 4428
rect 32218 4448 32220 4457
rect 32272 4448 32274 4457
rect 31588 4282 31616 4422
rect 32218 4383 32274 4392
rect 31576 4276 31628 4282
rect 31576 4218 31628 4224
rect 31208 4140 31260 4146
rect 31208 4082 31260 4088
rect 31484 4140 31536 4146
rect 31484 4082 31536 4088
rect 31588 3534 31616 4218
rect 32036 3936 32088 3942
rect 32036 3878 32088 3884
rect 32048 3534 32076 3878
rect 32220 3596 32272 3602
rect 32220 3538 32272 3544
rect 31576 3528 31628 3534
rect 31576 3470 31628 3476
rect 32036 3528 32088 3534
rect 32036 3470 32088 3476
rect 32232 3126 32260 3538
rect 32220 3120 32272 3126
rect 32220 3062 32272 3068
rect 31576 2984 31628 2990
rect 31576 2926 31628 2932
rect 31300 2508 31352 2514
rect 31300 2450 31352 2456
rect 30932 2440 30984 2446
rect 30932 2382 30984 2388
rect 31024 2372 31076 2378
rect 31024 2314 31076 2320
rect 31036 800 31064 2314
rect 31312 800 31340 2450
rect 31588 800 31616 2926
rect 32324 2428 32352 9007
rect 32588 8832 32640 8838
rect 32588 8774 32640 8780
rect 32494 8256 32550 8265
rect 32494 8191 32550 8200
rect 32404 8084 32456 8090
rect 32404 8026 32456 8032
rect 32416 4536 32444 8026
rect 32508 8022 32536 8191
rect 32496 8016 32548 8022
rect 32496 7958 32548 7964
rect 32600 7410 32628 8774
rect 32588 7404 32640 7410
rect 32588 7346 32640 7352
rect 32692 6798 32720 9522
rect 32784 8537 32812 10950
rect 32968 10130 32996 12174
rect 33152 11762 33180 12702
rect 33232 12640 33284 12646
rect 33232 12582 33284 12588
rect 33140 11756 33192 11762
rect 33140 11698 33192 11704
rect 33140 11620 33192 11626
rect 33140 11562 33192 11568
rect 33152 11234 33180 11562
rect 33060 11206 33180 11234
rect 32956 10124 33008 10130
rect 32956 10066 33008 10072
rect 33060 9874 33088 11206
rect 32876 9846 33088 9874
rect 32770 8528 32826 8537
rect 32770 8463 32772 8472
rect 32824 8463 32826 8472
rect 32772 8434 32824 8440
rect 32772 7404 32824 7410
rect 32772 7346 32824 7352
rect 32680 6792 32732 6798
rect 32680 6734 32732 6740
rect 32586 6352 32642 6361
rect 32586 6287 32642 6296
rect 32600 5681 32628 6287
rect 32784 6186 32812 7346
rect 32772 6180 32824 6186
rect 32772 6122 32824 6128
rect 32876 5953 32904 9846
rect 32956 9716 33008 9722
rect 32956 9658 33008 9664
rect 32968 8809 32996 9658
rect 33140 9512 33192 9518
rect 33140 9454 33192 9460
rect 33152 9110 33180 9454
rect 33244 9217 33272 12582
rect 33428 12458 33456 12718
rect 33520 12646 33548 14214
rect 33508 12640 33560 12646
rect 33508 12582 33560 12588
rect 33336 12434 33456 12458
rect 33336 12406 33548 12434
rect 33414 10704 33470 10713
rect 33414 10639 33470 10648
rect 33324 10532 33376 10538
rect 33324 10474 33376 10480
rect 33336 10062 33364 10474
rect 33428 10062 33456 10639
rect 33324 10056 33376 10062
rect 33324 9998 33376 10004
rect 33416 10056 33468 10062
rect 33416 9998 33468 10004
rect 33324 9716 33376 9722
rect 33324 9658 33376 9664
rect 33230 9208 33286 9217
rect 33230 9143 33286 9152
rect 33140 9104 33192 9110
rect 33336 9092 33364 9658
rect 33414 9616 33470 9625
rect 33414 9551 33416 9560
rect 33468 9551 33470 9560
rect 33416 9522 33468 9528
rect 33140 9046 33192 9052
rect 33244 9064 33364 9092
rect 33152 8974 33180 9046
rect 33140 8968 33192 8974
rect 33140 8910 33192 8916
rect 33140 8832 33192 8838
rect 32954 8800 33010 8809
rect 32954 8735 33010 8744
rect 33060 8792 33140 8820
rect 33060 7750 33088 8792
rect 33140 8774 33192 8780
rect 33140 8492 33192 8498
rect 33140 8434 33192 8440
rect 33152 8022 33180 8434
rect 33140 8016 33192 8022
rect 33140 7958 33192 7964
rect 33140 7812 33192 7818
rect 33140 7754 33192 7760
rect 33048 7744 33100 7750
rect 33048 7686 33100 7692
rect 32956 6792 33008 6798
rect 32956 6734 33008 6740
rect 32862 5944 32918 5953
rect 32862 5879 32918 5888
rect 32968 5710 32996 6734
rect 33060 6662 33088 7686
rect 33152 7342 33180 7754
rect 33244 7410 33272 9064
rect 33520 8566 33548 12406
rect 33508 8560 33560 8566
rect 33508 8502 33560 8508
rect 33416 8356 33468 8362
rect 33416 8298 33468 8304
rect 33324 8016 33376 8022
rect 33324 7958 33376 7964
rect 33232 7404 33284 7410
rect 33232 7346 33284 7352
rect 33140 7336 33192 7342
rect 33140 7278 33192 7284
rect 33140 6860 33192 6866
rect 33140 6802 33192 6808
rect 33048 6656 33100 6662
rect 33048 6598 33100 6604
rect 33152 6254 33180 6802
rect 33232 6724 33284 6730
rect 33232 6666 33284 6672
rect 33140 6248 33192 6254
rect 33140 6190 33192 6196
rect 32956 5704 33008 5710
rect 32586 5672 32642 5681
rect 32956 5646 33008 5652
rect 32586 5607 32642 5616
rect 32586 5400 32642 5409
rect 32586 5335 32642 5344
rect 32600 5302 32628 5335
rect 32588 5296 32640 5302
rect 32588 5238 32640 5244
rect 33048 5092 33100 5098
rect 33048 5034 33100 5040
rect 32864 4684 32916 4690
rect 32864 4626 32916 4632
rect 32496 4548 32548 4554
rect 32416 4508 32496 4536
rect 32496 4490 32548 4496
rect 32876 4078 32904 4626
rect 32772 4072 32824 4078
rect 32770 4040 32772 4049
rect 32864 4072 32916 4078
rect 32824 4040 32826 4049
rect 32680 4004 32732 4010
rect 32864 4014 32916 4020
rect 32770 3975 32826 3984
rect 32680 3946 32732 3952
rect 32496 2848 32548 2854
rect 32496 2790 32548 2796
rect 32404 2440 32456 2446
rect 32324 2400 32404 2428
rect 32404 2382 32456 2388
rect 31852 2372 31904 2378
rect 31852 2314 31904 2320
rect 31864 800 31892 2314
rect 32128 2304 32180 2310
rect 32128 2246 32180 2252
rect 32140 800 32168 2246
rect 32508 1442 32536 2790
rect 32416 1414 32536 1442
rect 32416 800 32444 1414
rect 32692 800 32720 3946
rect 32784 2961 32812 3975
rect 32864 3528 32916 3534
rect 32864 3470 32916 3476
rect 32876 3398 32904 3470
rect 32864 3392 32916 3398
rect 32864 3334 32916 3340
rect 32956 3392 33008 3398
rect 32956 3334 33008 3340
rect 32770 2952 32826 2961
rect 32770 2887 32826 2896
rect 32968 800 32996 3334
rect 33060 3194 33088 5034
rect 33152 4622 33180 6190
rect 33244 5166 33272 6666
rect 33336 6186 33364 7958
rect 33324 6180 33376 6186
rect 33324 6122 33376 6128
rect 33232 5160 33284 5166
rect 33232 5102 33284 5108
rect 33140 4616 33192 4622
rect 33140 4558 33192 4564
rect 33152 4457 33180 4558
rect 33138 4448 33194 4457
rect 33138 4383 33194 4392
rect 33336 4282 33364 6122
rect 33428 4865 33456 8298
rect 33520 5545 33548 8502
rect 33612 7886 33640 14214
rect 33968 12844 34020 12850
rect 33968 12786 34020 12792
rect 33876 12164 33928 12170
rect 33876 12106 33928 12112
rect 33784 11144 33836 11150
rect 33784 11086 33836 11092
rect 33692 9988 33744 9994
rect 33692 9930 33744 9936
rect 33704 9722 33732 9930
rect 33692 9716 33744 9722
rect 33692 9658 33744 9664
rect 33692 9580 33744 9586
rect 33692 9522 33744 9528
rect 33704 9178 33732 9522
rect 33692 9172 33744 9178
rect 33692 9114 33744 9120
rect 33704 8906 33732 9114
rect 33692 8900 33744 8906
rect 33692 8842 33744 8848
rect 33704 8498 33732 8842
rect 33692 8492 33744 8498
rect 33692 8434 33744 8440
rect 33600 7880 33652 7886
rect 33600 7822 33652 7828
rect 33704 7177 33732 8434
rect 33690 7168 33746 7177
rect 33690 7103 33746 7112
rect 33692 6792 33744 6798
rect 33692 6734 33744 6740
rect 33704 6390 33732 6734
rect 33796 6458 33824 11086
rect 33888 11082 33916 12106
rect 33980 11762 34008 12786
rect 33968 11756 34020 11762
rect 33968 11698 34020 11704
rect 34072 11150 34100 28426
rect 34520 25832 34572 25838
rect 34520 25774 34572 25780
rect 34532 18630 34560 25774
rect 34704 21344 34756 21350
rect 34704 21286 34756 21292
rect 34612 20460 34664 20466
rect 34612 20402 34664 20408
rect 34624 19514 34652 20402
rect 34612 19508 34664 19514
rect 34612 19450 34664 19456
rect 34716 19394 34744 21286
rect 34624 19366 34744 19394
rect 34520 18624 34572 18630
rect 34520 18566 34572 18572
rect 34428 18080 34480 18086
rect 34428 18022 34480 18028
rect 34440 17678 34468 18022
rect 34428 17672 34480 17678
rect 34428 17614 34480 17620
rect 34520 17604 34572 17610
rect 34520 17546 34572 17552
rect 34336 17536 34388 17542
rect 34336 17478 34388 17484
rect 34348 16454 34376 17478
rect 34532 17377 34560 17546
rect 34518 17368 34574 17377
rect 34518 17303 34574 17312
rect 34336 16448 34388 16454
rect 34336 16390 34388 16396
rect 34152 15496 34204 15502
rect 34152 15438 34204 15444
rect 34164 12084 34192 15438
rect 34348 15434 34376 16390
rect 34336 15428 34388 15434
rect 34336 15370 34388 15376
rect 34336 14816 34388 14822
rect 34336 14758 34388 14764
rect 34348 14362 34376 14758
rect 34624 14482 34652 19366
rect 34704 19304 34756 19310
rect 34704 19246 34756 19252
rect 34716 18290 34744 19246
rect 34704 18284 34756 18290
rect 34704 18226 34756 18232
rect 34704 15020 34756 15026
rect 34704 14962 34756 14968
rect 34612 14476 34664 14482
rect 34612 14418 34664 14424
rect 34348 14334 34560 14362
rect 34532 14074 34560 14334
rect 34716 14260 34744 14962
rect 34808 14362 34836 42638
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 35820 33522 35848 47534
rect 35912 43722 35940 61066
rect 36084 61056 36136 61062
rect 36084 60998 36136 61004
rect 35992 57928 36044 57934
rect 35992 57870 36044 57876
rect 36004 57526 36032 57870
rect 35992 57520 36044 57526
rect 35992 57462 36044 57468
rect 35992 45416 36044 45422
rect 35992 45358 36044 45364
rect 35900 43716 35952 43722
rect 35900 43658 35952 43664
rect 36004 33522 36032 45358
rect 36096 33590 36124 60998
rect 36372 60790 36400 63294
rect 36910 63294 37228 63322
rect 36910 63200 36966 63294
rect 37200 61180 37228 63294
rect 37646 63200 37702 64000
rect 38382 63322 38438 64000
rect 39118 63322 39174 64000
rect 39854 63322 39910 64000
rect 38382 63294 38608 63322
rect 38382 63200 38438 63294
rect 37660 61198 37688 63200
rect 37280 61192 37332 61198
rect 37200 61152 37280 61180
rect 37280 61134 37332 61140
rect 37648 61192 37700 61198
rect 38580 61180 38608 63294
rect 39118 63294 39528 63322
rect 39118 63200 39174 63294
rect 39500 61198 39528 63294
rect 39854 63294 39988 63322
rect 39854 63200 39910 63294
rect 38660 61192 38712 61198
rect 38580 61152 38660 61180
rect 37648 61134 37700 61140
rect 38660 61134 38712 61140
rect 39488 61192 39540 61198
rect 39488 61134 39540 61140
rect 39960 61130 39988 63294
rect 40590 63200 40646 64000
rect 41326 63200 41382 64000
rect 42062 63200 42118 64000
rect 42798 63200 42854 64000
rect 43534 63200 43590 64000
rect 44270 63322 44326 64000
rect 45006 63322 45062 64000
rect 45742 63322 45798 64000
rect 46478 63322 46534 64000
rect 44270 63294 44588 63322
rect 44270 63200 44326 63294
rect 40224 61600 40276 61606
rect 40224 61542 40276 61548
rect 40236 61402 40264 61542
rect 40224 61396 40276 61402
rect 40224 61338 40276 61344
rect 40604 61198 40632 63200
rect 40592 61192 40644 61198
rect 40592 61134 40644 61140
rect 38016 61124 38068 61130
rect 38016 61066 38068 61072
rect 39948 61124 40000 61130
rect 39948 61066 40000 61072
rect 36360 60784 36412 60790
rect 36360 60726 36412 60732
rect 38028 58546 38056 61066
rect 39120 61056 39172 61062
rect 39120 60998 39172 61004
rect 40316 61056 40368 61062
rect 40316 60998 40368 61004
rect 37924 58540 37976 58546
rect 37924 58482 37976 58488
rect 38016 58540 38068 58546
rect 38016 58482 38068 58488
rect 36912 58472 36964 58478
rect 36912 58414 36964 58420
rect 36268 57928 36320 57934
rect 36268 57870 36320 57876
rect 36280 56846 36308 57870
rect 36268 56840 36320 56846
rect 36268 56782 36320 56788
rect 36280 36854 36308 56782
rect 36360 46368 36412 46374
rect 36360 46310 36412 46316
rect 36372 45490 36400 46310
rect 36360 45484 36412 45490
rect 36360 45426 36412 45432
rect 36636 45484 36688 45490
rect 36636 45426 36688 45432
rect 36648 40458 36676 45426
rect 36924 45354 36952 58414
rect 37188 58404 37240 58410
rect 37188 58346 37240 58352
rect 37200 45422 37228 58346
rect 37936 58342 37964 58482
rect 37556 58336 37608 58342
rect 37556 58278 37608 58284
rect 37924 58336 37976 58342
rect 37924 58278 37976 58284
rect 37464 45484 37516 45490
rect 37464 45426 37516 45432
rect 37188 45416 37240 45422
rect 37188 45358 37240 45364
rect 36912 45348 36964 45354
rect 36912 45290 36964 45296
rect 36820 44804 36872 44810
rect 36820 44746 36872 44752
rect 36636 40452 36688 40458
rect 36636 40394 36688 40400
rect 36268 36848 36320 36854
rect 36268 36790 36320 36796
rect 36084 33584 36136 33590
rect 36084 33526 36136 33532
rect 35808 33516 35860 33522
rect 35808 33458 35860 33464
rect 35992 33516 36044 33522
rect 35992 33458 36044 33464
rect 36004 33386 36032 33458
rect 35992 33380 36044 33386
rect 35992 33322 36044 33328
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 35532 29708 35584 29714
rect 35532 29650 35584 29656
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34888 20936 34940 20942
rect 34888 20878 34940 20884
rect 34900 20534 34928 20878
rect 34888 20528 34940 20534
rect 34888 20470 34940 20476
rect 35348 20392 35400 20398
rect 35348 20334 35400 20340
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 35360 20058 35388 20334
rect 35348 20052 35400 20058
rect 35348 19994 35400 20000
rect 35070 19952 35126 19961
rect 35070 19887 35126 19896
rect 35084 19514 35112 19887
rect 35072 19508 35124 19514
rect 35072 19450 35124 19456
rect 35084 19310 35112 19450
rect 35072 19304 35124 19310
rect 35072 19246 35124 19252
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35440 18624 35492 18630
rect 35440 18566 35492 18572
rect 35348 18216 35400 18222
rect 35348 18158 35400 18164
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35164 17740 35216 17746
rect 35164 17682 35216 17688
rect 35176 17649 35204 17682
rect 35256 17672 35308 17678
rect 35162 17640 35218 17649
rect 35256 17614 35308 17620
rect 35162 17575 35218 17584
rect 35268 17270 35296 17614
rect 35256 17264 35308 17270
rect 35256 17206 35308 17212
rect 35360 16998 35388 18158
rect 35348 16992 35400 16998
rect 35348 16934 35400 16940
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35360 16794 35388 16934
rect 35348 16788 35400 16794
rect 35348 16730 35400 16736
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35256 14612 35308 14618
rect 35256 14554 35308 14560
rect 35072 14476 35124 14482
rect 35072 14418 35124 14424
rect 35164 14476 35216 14482
rect 35164 14418 35216 14424
rect 34808 14334 35020 14362
rect 34888 14272 34940 14278
rect 34716 14232 34888 14260
rect 34888 14214 34940 14220
rect 34992 14090 35020 14334
rect 35084 14278 35112 14418
rect 35072 14272 35124 14278
rect 35072 14214 35124 14220
rect 34520 14068 34572 14074
rect 34520 14010 34572 14016
rect 34808 14062 35020 14090
rect 34612 13864 34664 13870
rect 34612 13806 34664 13812
rect 34520 13728 34572 13734
rect 34520 13670 34572 13676
rect 34532 12850 34560 13670
rect 34520 12844 34572 12850
rect 34520 12786 34572 12792
rect 34242 12744 34298 12753
rect 34624 12730 34652 13806
rect 34704 13728 34756 13734
rect 34704 13670 34756 13676
rect 34716 13190 34744 13670
rect 34704 13184 34756 13190
rect 34704 13126 34756 13132
rect 34704 12844 34756 12850
rect 34704 12786 34756 12792
rect 34242 12679 34298 12688
rect 34532 12702 34652 12730
rect 34256 12238 34284 12679
rect 34532 12646 34560 12702
rect 34520 12640 34572 12646
rect 34520 12582 34572 12588
rect 34244 12232 34296 12238
rect 34244 12174 34296 12180
rect 34164 12056 34284 12084
rect 34152 11824 34204 11830
rect 34152 11766 34204 11772
rect 34060 11144 34112 11150
rect 34060 11086 34112 11092
rect 33876 11076 33928 11082
rect 33876 11018 33928 11024
rect 33888 10198 33916 11018
rect 34060 11008 34112 11014
rect 34060 10950 34112 10956
rect 33876 10192 33928 10198
rect 33928 10152 34008 10180
rect 33876 10134 33928 10140
rect 33980 9654 34008 10152
rect 33968 9648 34020 9654
rect 33968 9590 34020 9596
rect 33876 9512 33928 9518
rect 33876 9454 33928 9460
rect 33888 8537 33916 9454
rect 33874 8528 33930 8537
rect 33874 8463 33876 8472
rect 33928 8463 33930 8472
rect 33876 8434 33928 8440
rect 33968 8288 34020 8294
rect 33968 8230 34020 8236
rect 33980 8090 34008 8230
rect 33968 8084 34020 8090
rect 33968 8026 34020 8032
rect 33876 7268 33928 7274
rect 33876 7210 33928 7216
rect 33784 6452 33836 6458
rect 33784 6394 33836 6400
rect 33692 6384 33744 6390
rect 33692 6326 33744 6332
rect 33888 6322 33916 7210
rect 33876 6316 33928 6322
rect 33796 6276 33876 6304
rect 33796 5710 33824 6276
rect 33876 6258 33928 6264
rect 34072 5794 34100 10950
rect 34164 9994 34192 11766
rect 34256 10130 34284 12056
rect 34428 11144 34480 11150
rect 34428 11086 34480 11092
rect 34336 11008 34388 11014
rect 34336 10950 34388 10956
rect 34348 10742 34376 10950
rect 34336 10736 34388 10742
rect 34336 10678 34388 10684
rect 34440 10441 34468 11086
rect 34426 10432 34482 10441
rect 34426 10367 34482 10376
rect 34428 10260 34480 10266
rect 34428 10202 34480 10208
rect 34244 10124 34296 10130
rect 34244 10066 34296 10072
rect 34152 9988 34204 9994
rect 34152 9930 34204 9936
rect 34152 9172 34204 9178
rect 34440 9160 34468 10202
rect 34532 9450 34560 12582
rect 34520 9444 34572 9450
rect 34520 9386 34572 9392
rect 34152 9114 34204 9120
rect 34348 9132 34468 9160
rect 34164 7886 34192 9114
rect 34244 8968 34296 8974
rect 34348 8945 34376 9132
rect 34428 9036 34480 9042
rect 34428 8978 34480 8984
rect 34244 8910 34296 8916
rect 34334 8936 34390 8945
rect 34256 8634 34284 8910
rect 34334 8871 34390 8880
rect 34244 8628 34296 8634
rect 34244 8570 34296 8576
rect 34440 8498 34468 8978
rect 34428 8492 34480 8498
rect 34428 8434 34480 8440
rect 34428 8288 34480 8294
rect 34428 8230 34480 8236
rect 34152 7880 34204 7886
rect 34152 7822 34204 7828
rect 34152 7744 34204 7750
rect 34152 7686 34204 7692
rect 33888 5766 34100 5794
rect 33784 5704 33836 5710
rect 33784 5646 33836 5652
rect 33506 5536 33562 5545
rect 33506 5471 33562 5480
rect 33796 5302 33824 5646
rect 33784 5296 33836 5302
rect 33784 5238 33836 5244
rect 33414 4856 33470 4865
rect 33414 4791 33470 4800
rect 33416 4480 33468 4486
rect 33416 4422 33468 4428
rect 33508 4480 33560 4486
rect 33508 4422 33560 4428
rect 33324 4276 33376 4282
rect 33324 4218 33376 4224
rect 33428 4214 33456 4422
rect 33416 4208 33468 4214
rect 33416 4150 33468 4156
rect 33416 3936 33468 3942
rect 33416 3878 33468 3884
rect 33232 3596 33284 3602
rect 33232 3538 33284 3544
rect 33048 3188 33100 3194
rect 33048 3130 33100 3136
rect 33244 800 33272 3538
rect 33428 3534 33456 3878
rect 33324 3528 33376 3534
rect 33324 3470 33376 3476
rect 33416 3528 33468 3534
rect 33416 3470 33468 3476
rect 33336 3398 33364 3470
rect 33324 3392 33376 3398
rect 33324 3334 33376 3340
rect 33520 2990 33548 4422
rect 33692 4276 33744 4282
rect 33692 4218 33744 4224
rect 33600 3936 33652 3942
rect 33600 3878 33652 3884
rect 33508 2984 33560 2990
rect 33508 2926 33560 2932
rect 33612 2020 33640 3878
rect 33704 3738 33732 4218
rect 33692 3732 33744 3738
rect 33692 3674 33744 3680
rect 33888 3398 33916 5766
rect 34060 5636 34112 5642
rect 34060 5578 34112 5584
rect 34072 4078 34100 5578
rect 34164 5409 34192 7686
rect 34336 7404 34388 7410
rect 34336 7346 34388 7352
rect 34348 7002 34376 7346
rect 34336 6996 34388 7002
rect 34336 6938 34388 6944
rect 34440 6866 34468 8230
rect 34612 8016 34664 8022
rect 34612 7958 34664 7964
rect 34428 6860 34480 6866
rect 34428 6802 34480 6808
rect 34624 6322 34652 7958
rect 34716 7818 34744 12786
rect 34808 10606 34836 14062
rect 35176 13870 35204 14418
rect 35268 14385 35296 14554
rect 35254 14376 35310 14385
rect 35254 14311 35310 14320
rect 35164 13864 35216 13870
rect 35164 13806 35216 13812
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 35348 12232 35400 12238
rect 35346 12200 35348 12209
rect 35400 12200 35402 12209
rect 35346 12135 35402 12144
rect 35348 11756 35400 11762
rect 35348 11698 35400 11704
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 35360 11354 35388 11698
rect 35348 11348 35400 11354
rect 35348 11290 35400 11296
rect 35254 10840 35310 10849
rect 34980 10804 35032 10810
rect 35254 10775 35310 10784
rect 34980 10746 35032 10752
rect 34796 10600 34848 10606
rect 34796 10542 34848 10548
rect 34992 10470 35020 10746
rect 35268 10674 35296 10775
rect 35256 10668 35308 10674
rect 35256 10610 35308 10616
rect 34980 10464 35032 10470
rect 34980 10406 35032 10412
rect 35348 10464 35400 10470
rect 35348 10406 35400 10412
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 35360 10130 35388 10406
rect 34796 10124 34848 10130
rect 34796 10066 34848 10072
rect 35348 10124 35400 10130
rect 35348 10066 35400 10072
rect 34704 7812 34756 7818
rect 34704 7754 34756 7760
rect 34704 7404 34756 7410
rect 34704 7346 34756 7352
rect 34612 6316 34664 6322
rect 34612 6258 34664 6264
rect 34716 6202 34744 7346
rect 34624 6174 34744 6202
rect 34244 5568 34296 5574
rect 34244 5510 34296 5516
rect 34150 5400 34206 5409
rect 34150 5335 34206 5344
rect 34152 5024 34204 5030
rect 34152 4966 34204 4972
rect 34164 4282 34192 4966
rect 34152 4276 34204 4282
rect 34152 4218 34204 4224
rect 34060 4072 34112 4078
rect 34060 4014 34112 4020
rect 33968 3528 34020 3534
rect 33968 3470 34020 3476
rect 33876 3392 33928 3398
rect 33876 3334 33928 3340
rect 33876 2984 33928 2990
rect 33520 1992 33640 2020
rect 33796 2944 33876 2972
rect 33520 800 33548 1992
rect 33796 800 33824 2944
rect 33876 2926 33928 2932
rect 33980 2774 34008 3470
rect 34060 3392 34112 3398
rect 34060 3334 34112 3340
rect 33888 2746 34008 2774
rect 33888 2378 33916 2746
rect 33876 2372 33928 2378
rect 33876 2314 33928 2320
rect 34072 800 34100 3334
rect 34256 2582 34284 5510
rect 34428 5024 34480 5030
rect 34428 4966 34480 4972
rect 34440 4146 34468 4966
rect 34624 4729 34652 6174
rect 34808 5710 34836 10066
rect 35164 9988 35216 9994
rect 35164 9930 35216 9936
rect 35348 9988 35400 9994
rect 35348 9930 35400 9936
rect 35176 9450 35204 9930
rect 35164 9444 35216 9450
rect 35164 9386 35216 9392
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 35360 8634 35388 9930
rect 35348 8628 35400 8634
rect 35348 8570 35400 8576
rect 35452 8378 35480 18566
rect 35544 12306 35572 29650
rect 36636 26920 36688 26926
rect 36636 26862 36688 26868
rect 36648 22094 36676 26862
rect 36556 22066 36676 22094
rect 35992 21956 36044 21962
rect 35992 21898 36044 21904
rect 35808 21888 35860 21894
rect 35808 21830 35860 21836
rect 35820 21486 35848 21830
rect 35900 21548 35952 21554
rect 35900 21490 35952 21496
rect 35808 21480 35860 21486
rect 35808 21422 35860 21428
rect 35624 21344 35676 21350
rect 35624 21286 35676 21292
rect 35716 21344 35768 21350
rect 35716 21286 35768 21292
rect 35636 19854 35664 21286
rect 35624 19848 35676 19854
rect 35624 19790 35676 19796
rect 35728 19802 35756 21286
rect 35808 20392 35860 20398
rect 35808 20334 35860 20340
rect 35820 19990 35848 20334
rect 35912 20262 35940 21490
rect 36004 21010 36032 21898
rect 35992 21004 36044 21010
rect 35992 20946 36044 20952
rect 36084 20460 36136 20466
rect 36084 20402 36136 20408
rect 35900 20256 35952 20262
rect 35900 20198 35952 20204
rect 35808 19984 35860 19990
rect 35808 19926 35860 19932
rect 35728 19774 35848 19802
rect 35912 19786 35940 20198
rect 35716 19168 35768 19174
rect 35716 19110 35768 19116
rect 35728 18902 35756 19110
rect 35716 18896 35768 18902
rect 35716 18838 35768 18844
rect 35624 18216 35676 18222
rect 35624 18158 35676 18164
rect 35636 14482 35664 18158
rect 35624 14476 35676 14482
rect 35624 14418 35676 14424
rect 35624 14068 35676 14074
rect 35624 14010 35676 14016
rect 35532 12300 35584 12306
rect 35532 12242 35584 12248
rect 35532 10668 35584 10674
rect 35532 10610 35584 10616
rect 35544 10266 35572 10610
rect 35532 10260 35584 10266
rect 35532 10202 35584 10208
rect 35530 10160 35586 10169
rect 35530 10095 35586 10104
rect 35544 9353 35572 10095
rect 35530 9344 35586 9353
rect 35530 9279 35586 9288
rect 35452 8350 35572 8378
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 35164 7880 35216 7886
rect 35164 7822 35216 7828
rect 35176 7478 35204 7822
rect 35438 7576 35494 7585
rect 35438 7511 35440 7520
rect 35492 7511 35494 7520
rect 35440 7482 35492 7488
rect 35164 7472 35216 7478
rect 35164 7414 35216 7420
rect 35348 7472 35400 7478
rect 35348 7414 35400 7420
rect 35360 7342 35388 7414
rect 35348 7336 35400 7342
rect 35348 7278 35400 7284
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 35360 6866 35388 7278
rect 35348 6860 35400 6866
rect 35348 6802 35400 6808
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 35360 5778 35388 6802
rect 35452 6322 35480 7482
rect 35440 6316 35492 6322
rect 35440 6258 35492 6264
rect 35440 6112 35492 6118
rect 35440 6054 35492 6060
rect 35348 5772 35400 5778
rect 35348 5714 35400 5720
rect 35452 5710 35480 6054
rect 34796 5704 34848 5710
rect 34796 5646 34848 5652
rect 35440 5704 35492 5710
rect 35440 5646 35492 5652
rect 34808 5302 34836 5646
rect 34796 5296 34848 5302
rect 34796 5238 34848 5244
rect 35348 5228 35400 5234
rect 35348 5170 35400 5176
rect 34796 5160 34848 5166
rect 34796 5102 34848 5108
rect 34704 5024 34756 5030
rect 34704 4966 34756 4972
rect 34610 4720 34666 4729
rect 34610 4655 34666 4664
rect 34520 4548 34572 4554
rect 34520 4490 34572 4496
rect 34428 4140 34480 4146
rect 34428 4082 34480 4088
rect 34336 3460 34388 3466
rect 34336 3402 34388 3408
rect 34348 2990 34376 3402
rect 34532 3058 34560 4490
rect 34716 3534 34744 4966
rect 34704 3528 34756 3534
rect 34704 3470 34756 3476
rect 34612 3460 34664 3466
rect 34612 3402 34664 3408
rect 34520 3052 34572 3058
rect 34520 2994 34572 3000
rect 34336 2984 34388 2990
rect 34336 2926 34388 2932
rect 34520 2848 34572 2854
rect 34520 2790 34572 2796
rect 34336 2644 34388 2650
rect 34336 2586 34388 2592
rect 34244 2576 34296 2582
rect 34244 2518 34296 2524
rect 34348 800 34376 2586
rect 34532 2514 34560 2790
rect 34520 2508 34572 2514
rect 34520 2450 34572 2456
rect 34624 800 34652 3402
rect 34808 1442 34836 5102
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 35360 4826 35388 5170
rect 35440 5160 35492 5166
rect 35440 5102 35492 5108
rect 35348 4820 35400 4826
rect 35348 4762 35400 4768
rect 35452 4026 35480 5102
rect 35360 3998 35480 4026
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34888 2440 34940 2446
rect 34888 2382 34940 2388
rect 34900 1970 34928 2382
rect 34888 1964 34940 1970
rect 34888 1906 34940 1912
rect 35360 1442 35388 3998
rect 35440 3936 35492 3942
rect 35440 3878 35492 3884
rect 35452 3398 35480 3878
rect 35440 3392 35492 3398
rect 35440 3334 35492 3340
rect 35544 2310 35572 8350
rect 35636 8022 35664 14010
rect 35728 13938 35756 18838
rect 35820 16674 35848 19774
rect 35900 19780 35952 19786
rect 35900 19722 35952 19728
rect 35912 18766 35940 19722
rect 36096 19514 36124 20402
rect 36360 19712 36412 19718
rect 36360 19654 36412 19660
rect 36372 19514 36400 19654
rect 36084 19508 36136 19514
rect 36084 19450 36136 19456
rect 36360 19508 36412 19514
rect 36360 19450 36412 19456
rect 36452 19508 36504 19514
rect 36452 19450 36504 19456
rect 36464 19258 36492 19450
rect 36372 19230 36492 19258
rect 36372 18902 36400 19230
rect 36452 19168 36504 19174
rect 36452 19110 36504 19116
rect 36464 18970 36492 19110
rect 36452 18964 36504 18970
rect 36452 18906 36504 18912
rect 36360 18896 36412 18902
rect 36360 18838 36412 18844
rect 35900 18760 35952 18766
rect 35900 18702 35952 18708
rect 36556 17513 36584 22066
rect 36636 21480 36688 21486
rect 36636 21422 36688 21428
rect 36648 20874 36676 21422
rect 36636 20868 36688 20874
rect 36636 20810 36688 20816
rect 36648 19310 36676 20810
rect 36636 19304 36688 19310
rect 36636 19246 36688 19252
rect 36648 18086 36676 19246
rect 36728 18692 36780 18698
rect 36728 18634 36780 18640
rect 36636 18080 36688 18086
rect 36636 18022 36688 18028
rect 36542 17504 36598 17513
rect 36542 17439 36598 17448
rect 35992 17264 36044 17270
rect 35992 17206 36044 17212
rect 35820 16646 35940 16674
rect 35912 15994 35940 16646
rect 35820 15966 35940 15994
rect 35716 13932 35768 13938
rect 35716 13874 35768 13880
rect 35820 13818 35848 15966
rect 36004 15910 36032 17206
rect 36084 16652 36136 16658
rect 36084 16594 36136 16600
rect 35992 15904 36044 15910
rect 35992 15846 36044 15852
rect 35900 14816 35952 14822
rect 35900 14758 35952 14764
rect 35912 14278 35940 14758
rect 35992 14544 36044 14550
rect 35992 14486 36044 14492
rect 35900 14272 35952 14278
rect 35900 14214 35952 14220
rect 35728 13790 35848 13818
rect 35728 11150 35756 13790
rect 35808 13456 35860 13462
rect 35808 13398 35860 13404
rect 35820 12850 35848 13398
rect 36004 13258 36032 14486
rect 35992 13252 36044 13258
rect 35992 13194 36044 13200
rect 36004 12918 36032 13194
rect 35992 12912 36044 12918
rect 35992 12854 36044 12860
rect 35808 12844 35860 12850
rect 35808 12786 35860 12792
rect 36096 12434 36124 16594
rect 36360 16584 36412 16590
rect 36360 16526 36412 16532
rect 36372 15502 36400 16526
rect 36556 16522 36584 17439
rect 36740 16658 36768 18634
rect 36728 16652 36780 16658
rect 36728 16594 36780 16600
rect 36544 16516 36596 16522
rect 36544 16458 36596 16464
rect 36452 16448 36504 16454
rect 36452 16390 36504 16396
rect 36728 16448 36780 16454
rect 36728 16390 36780 16396
rect 36464 15502 36492 16390
rect 36360 15496 36412 15502
rect 36360 15438 36412 15444
rect 36452 15496 36504 15502
rect 36452 15438 36504 15444
rect 36372 15094 36400 15438
rect 36740 15366 36768 16390
rect 36728 15360 36780 15366
rect 36728 15302 36780 15308
rect 36360 15088 36412 15094
rect 36360 15030 36412 15036
rect 36268 13320 36320 13326
rect 36266 13288 36268 13297
rect 36360 13320 36412 13326
rect 36320 13288 36322 13297
rect 36360 13262 36412 13268
rect 36266 13223 36322 13232
rect 36268 12844 36320 12850
rect 36268 12786 36320 12792
rect 36280 12594 36308 12786
rect 36372 12714 36400 13262
rect 36636 13184 36688 13190
rect 36636 13126 36688 13132
rect 36450 12880 36506 12889
rect 36450 12815 36452 12824
rect 36504 12815 36506 12824
rect 36452 12786 36504 12792
rect 36360 12708 36412 12714
rect 36360 12650 36412 12656
rect 36280 12566 36400 12594
rect 36004 12406 36124 12434
rect 35808 12232 35860 12238
rect 35808 12174 35860 12180
rect 35900 12232 35952 12238
rect 35900 12174 35952 12180
rect 35820 12073 35848 12174
rect 35806 12064 35862 12073
rect 35806 11999 35862 12008
rect 35912 11830 35940 12174
rect 35900 11824 35952 11830
rect 35900 11766 35952 11772
rect 35808 11552 35860 11558
rect 35808 11494 35860 11500
rect 35820 11218 35848 11494
rect 36004 11218 36032 12406
rect 36082 12200 36138 12209
rect 36082 12135 36138 12144
rect 36096 11286 36124 12135
rect 36084 11280 36136 11286
rect 36084 11222 36136 11228
rect 35808 11212 35860 11218
rect 35808 11154 35860 11160
rect 35992 11212 36044 11218
rect 35992 11154 36044 11160
rect 35716 11144 35768 11150
rect 36004 11098 36032 11154
rect 35716 11086 35768 11092
rect 35820 11070 36032 11098
rect 36372 11082 36400 12566
rect 36360 11076 36412 11082
rect 35820 10996 35848 11070
rect 36360 11018 36412 11024
rect 35728 10968 35848 10996
rect 36084 11008 36136 11014
rect 35728 8022 35756 10968
rect 36084 10950 36136 10956
rect 36096 10713 36124 10950
rect 36082 10704 36138 10713
rect 36082 10639 36138 10648
rect 36174 10024 36230 10033
rect 36174 9959 36230 9968
rect 36188 9926 36216 9959
rect 36176 9920 36228 9926
rect 36176 9862 36228 9868
rect 35992 9580 36044 9586
rect 35992 9522 36044 9528
rect 35900 9376 35952 9382
rect 35900 9318 35952 9324
rect 35912 8974 35940 9318
rect 36004 9178 36032 9522
rect 35992 9172 36044 9178
rect 35992 9114 36044 9120
rect 35900 8968 35952 8974
rect 35900 8910 35952 8916
rect 35912 8498 35940 8910
rect 35992 8832 36044 8838
rect 35992 8774 36044 8780
rect 35900 8492 35952 8498
rect 35900 8434 35952 8440
rect 35808 8424 35860 8430
rect 35808 8366 35860 8372
rect 35820 8090 35848 8366
rect 35808 8084 35860 8090
rect 35808 8026 35860 8032
rect 35624 8016 35676 8022
rect 35624 7958 35676 7964
rect 35716 8016 35768 8022
rect 35716 7958 35768 7964
rect 35728 7410 35756 7958
rect 36004 7478 36032 8774
rect 35992 7472 36044 7478
rect 35992 7414 36044 7420
rect 35716 7404 35768 7410
rect 35716 7346 35768 7352
rect 35992 7200 36044 7206
rect 35992 7142 36044 7148
rect 35806 6760 35862 6769
rect 35624 6724 35676 6730
rect 35806 6695 35808 6704
rect 35624 6666 35676 6672
rect 35860 6695 35862 6704
rect 35808 6666 35860 6672
rect 35636 5370 35664 6666
rect 35900 6656 35952 6662
rect 35900 6598 35952 6604
rect 35912 6322 35940 6598
rect 35900 6316 35952 6322
rect 35900 6258 35952 6264
rect 35808 6248 35860 6254
rect 35808 6190 35860 6196
rect 35820 5846 35848 6190
rect 35900 6112 35952 6118
rect 35900 6054 35952 6060
rect 35808 5840 35860 5846
rect 35808 5782 35860 5788
rect 35624 5364 35676 5370
rect 35624 5306 35676 5312
rect 35912 5234 35940 6054
rect 35900 5228 35952 5234
rect 35900 5170 35952 5176
rect 35624 4616 35676 4622
rect 35624 4558 35676 4564
rect 35636 4010 35664 4558
rect 35716 4072 35768 4078
rect 36004 4049 36032 7142
rect 35716 4014 35768 4020
rect 35990 4040 36046 4049
rect 35624 4004 35676 4010
rect 35624 3946 35676 3952
rect 35636 3126 35664 3946
rect 35728 3466 35756 4014
rect 35990 3975 36046 3984
rect 36084 3596 36136 3602
rect 36084 3538 36136 3544
rect 35716 3460 35768 3466
rect 35716 3402 35768 3408
rect 35624 3120 35676 3126
rect 35624 3062 35676 3068
rect 36096 2990 36124 3538
rect 36188 3534 36216 9862
rect 36268 9376 36320 9382
rect 36268 9318 36320 9324
rect 36280 9042 36308 9318
rect 36464 9110 36492 12786
rect 36648 12306 36676 13126
rect 36636 12300 36688 12306
rect 36636 12242 36688 12248
rect 36740 11937 36768 15302
rect 36832 13938 36860 44746
rect 37280 42696 37332 42702
rect 37278 42664 37280 42673
rect 37332 42664 37334 42673
rect 37476 42634 37504 45426
rect 37278 42599 37334 42608
rect 37464 42628 37516 42634
rect 37464 42570 37516 42576
rect 37004 38888 37056 38894
rect 37004 38830 37056 38836
rect 37016 22094 37044 38830
rect 37476 37942 37504 42570
rect 37464 37936 37516 37942
rect 37464 37878 37516 37884
rect 37280 36712 37332 36718
rect 37280 36654 37332 36660
rect 37292 35834 37320 36654
rect 37280 35828 37332 35834
rect 37280 35770 37332 35776
rect 37568 32910 37596 58278
rect 37936 57390 37964 58278
rect 37924 57384 37976 57390
rect 37924 57326 37976 57332
rect 37924 46980 37976 46986
rect 37924 46922 37976 46928
rect 37648 33312 37700 33318
rect 37648 33254 37700 33260
rect 37556 32904 37608 32910
rect 37556 32846 37608 32852
rect 37280 28076 37332 28082
rect 37280 28018 37332 28024
rect 37292 22166 37320 28018
rect 37280 22160 37332 22166
rect 37280 22102 37332 22108
rect 36924 22066 37044 22094
rect 36820 13932 36872 13938
rect 36820 13874 36872 13880
rect 36924 12434 36952 22066
rect 37280 21004 37332 21010
rect 37280 20946 37332 20952
rect 37292 20398 37320 20946
rect 37280 20392 37332 20398
rect 37280 20334 37332 20340
rect 37292 19310 37320 20334
rect 37280 19304 37332 19310
rect 37280 19246 37332 19252
rect 37004 18964 37056 18970
rect 37004 18906 37056 18912
rect 37016 18601 37044 18906
rect 37188 18624 37240 18630
rect 37002 18592 37058 18601
rect 37188 18566 37240 18572
rect 37002 18527 37058 18536
rect 37200 16250 37228 18566
rect 37188 16244 37240 16250
rect 37188 16186 37240 16192
rect 37004 16040 37056 16046
rect 37004 15982 37056 15988
rect 36832 12406 36952 12434
rect 36726 11928 36782 11937
rect 36726 11863 36782 11872
rect 36544 11348 36596 11354
rect 36544 11290 36596 11296
rect 36556 10577 36584 11290
rect 36542 10568 36598 10577
rect 36542 10503 36598 10512
rect 36636 10124 36688 10130
rect 36636 10066 36688 10072
rect 36544 9580 36596 9586
rect 36544 9522 36596 9528
rect 36452 9104 36504 9110
rect 36450 9072 36452 9081
rect 36504 9072 36506 9081
rect 36268 9036 36320 9042
rect 36450 9007 36506 9016
rect 36268 8978 36320 8984
rect 36464 6662 36492 9007
rect 36556 7993 36584 9522
rect 36648 8809 36676 10066
rect 36634 8800 36690 8809
rect 36634 8735 36690 8744
rect 36542 7984 36598 7993
rect 36542 7919 36598 7928
rect 36556 7750 36584 7919
rect 36544 7744 36596 7750
rect 36544 7686 36596 7692
rect 36556 7410 36584 7686
rect 36544 7404 36596 7410
rect 36544 7346 36596 7352
rect 36648 7290 36676 8735
rect 36728 8492 36780 8498
rect 36728 8434 36780 8440
rect 36740 7546 36768 8434
rect 36728 7540 36780 7546
rect 36728 7482 36780 7488
rect 36832 7426 36860 12406
rect 36912 10260 36964 10266
rect 36912 10202 36964 10208
rect 36924 10062 36952 10202
rect 36912 10056 36964 10062
rect 36912 9998 36964 10004
rect 36912 8288 36964 8294
rect 36912 8230 36964 8236
rect 36924 7886 36952 8230
rect 36912 7880 36964 7886
rect 36912 7822 36964 7828
rect 36556 7262 36676 7290
rect 36740 7398 36860 7426
rect 36912 7404 36964 7410
rect 36452 6656 36504 6662
rect 36452 6598 36504 6604
rect 36268 6180 36320 6186
rect 36268 6122 36320 6128
rect 36280 4146 36308 6122
rect 36360 5568 36412 5574
rect 36360 5510 36412 5516
rect 36372 5409 36400 5510
rect 36358 5400 36414 5409
rect 36358 5335 36414 5344
rect 36372 4486 36400 5335
rect 36452 5296 36504 5302
rect 36452 5238 36504 5244
rect 36360 4480 36412 4486
rect 36360 4422 36412 4428
rect 36268 4140 36320 4146
rect 36268 4082 36320 4088
rect 36266 4040 36322 4049
rect 36266 3975 36322 3984
rect 36176 3528 36228 3534
rect 36176 3470 36228 3476
rect 36280 3058 36308 3975
rect 36358 3360 36414 3369
rect 36358 3295 36414 3304
rect 36268 3052 36320 3058
rect 36268 2994 36320 3000
rect 36084 2984 36136 2990
rect 36084 2926 36136 2932
rect 36372 2774 36400 3295
rect 36464 3058 36492 5238
rect 36556 4758 36584 7262
rect 36740 7154 36768 7398
rect 36912 7346 36964 7352
rect 36924 7206 36952 7346
rect 36648 7126 36768 7154
rect 36912 7200 36964 7206
rect 36912 7142 36964 7148
rect 36544 4752 36596 4758
rect 36544 4694 36596 4700
rect 36544 3392 36596 3398
rect 36544 3334 36596 3340
rect 36556 3126 36584 3334
rect 36544 3120 36596 3126
rect 36544 3062 36596 3068
rect 36452 3052 36504 3058
rect 36452 2994 36504 3000
rect 36542 2952 36598 2961
rect 36542 2887 36598 2896
rect 36280 2746 36400 2774
rect 35532 2304 35584 2310
rect 35532 2246 35584 2252
rect 35716 1556 35768 1562
rect 35716 1498 35768 1504
rect 34808 1414 34928 1442
rect 34900 800 34928 1414
rect 35176 1414 35388 1442
rect 35176 800 35204 1414
rect 35440 1216 35492 1222
rect 35440 1158 35492 1164
rect 35452 800 35480 1158
rect 35728 800 35756 1498
rect 35992 1420 36044 1426
rect 35992 1362 36044 1368
rect 36004 800 36032 1362
rect 36280 800 36308 2746
rect 36556 800 36584 2887
rect 36648 2378 36676 7126
rect 36728 6792 36780 6798
rect 36728 6734 36780 6740
rect 36740 6662 36768 6734
rect 36728 6656 36780 6662
rect 36728 6598 36780 6604
rect 36924 6186 36952 7142
rect 36912 6180 36964 6186
rect 36912 6122 36964 6128
rect 36820 4752 36872 4758
rect 36820 4694 36872 4700
rect 36728 4072 36780 4078
rect 36728 4014 36780 4020
rect 36636 2372 36688 2378
rect 36636 2314 36688 2320
rect 36740 1562 36768 4014
rect 36832 3602 36860 4694
rect 36820 3596 36872 3602
rect 36820 3538 36872 3544
rect 36820 2916 36872 2922
rect 36872 2876 36952 2904
rect 36820 2858 36872 2864
rect 36924 2514 36952 2876
rect 36912 2508 36964 2514
rect 36912 2450 36964 2456
rect 37016 2038 37044 15982
rect 37200 15910 37228 16186
rect 37188 15904 37240 15910
rect 37188 15846 37240 15852
rect 37292 13297 37320 19246
rect 37372 14408 37424 14414
rect 37372 14350 37424 14356
rect 37384 14074 37412 14350
rect 37372 14068 37424 14074
rect 37372 14010 37424 14016
rect 37372 13932 37424 13938
rect 37372 13874 37424 13880
rect 37278 13288 37334 13297
rect 37278 13223 37334 13232
rect 37292 13190 37320 13223
rect 37096 13184 37148 13190
rect 37096 13126 37148 13132
rect 37280 13184 37332 13190
rect 37280 13126 37332 13132
rect 37108 12782 37136 13126
rect 37188 12980 37240 12986
rect 37188 12922 37240 12928
rect 37096 12776 37148 12782
rect 37096 12718 37148 12724
rect 37108 12646 37136 12718
rect 37096 12640 37148 12646
rect 37096 12582 37148 12588
rect 37200 11898 37228 12922
rect 37188 11892 37240 11898
rect 37188 11834 37240 11840
rect 37096 11076 37148 11082
rect 37096 11018 37148 11024
rect 37108 8974 37136 11018
rect 37384 10062 37412 13874
rect 37462 13152 37518 13161
rect 37462 13087 37518 13096
rect 37476 10062 37504 13087
rect 37372 10056 37424 10062
rect 37372 9998 37424 10004
rect 37464 10056 37516 10062
rect 37464 9998 37516 10004
rect 37464 9920 37516 9926
rect 37464 9862 37516 9868
rect 37476 9586 37504 9862
rect 37464 9580 37516 9586
rect 37464 9522 37516 9528
rect 37556 9376 37608 9382
rect 37556 9318 37608 9324
rect 37188 9036 37240 9042
rect 37188 8978 37240 8984
rect 37096 8968 37148 8974
rect 37094 8936 37096 8945
rect 37148 8936 37150 8945
rect 37094 8871 37150 8880
rect 37096 8424 37148 8430
rect 37096 8366 37148 8372
rect 37108 3194 37136 8366
rect 37200 6866 37228 8978
rect 37464 8900 37516 8906
rect 37464 8842 37516 8848
rect 37280 8832 37332 8838
rect 37280 8774 37332 8780
rect 37292 8498 37320 8774
rect 37476 8673 37504 8842
rect 37462 8664 37518 8673
rect 37462 8599 37518 8608
rect 37568 8498 37596 9318
rect 37660 8566 37688 33254
rect 37832 20256 37884 20262
rect 37832 20198 37884 20204
rect 37844 19786 37872 20198
rect 37832 19780 37884 19786
rect 37832 19722 37884 19728
rect 37832 13320 37884 13326
rect 37832 13262 37884 13268
rect 37844 12850 37872 13262
rect 37832 12844 37884 12850
rect 37832 12786 37884 12792
rect 37936 12102 37964 46922
rect 38016 45484 38068 45490
rect 38016 45426 38068 45432
rect 38028 45393 38056 45426
rect 38014 45384 38070 45393
rect 38014 45319 38070 45328
rect 39132 34746 39160 60998
rect 39396 54528 39448 54534
rect 39396 54470 39448 54476
rect 39120 34740 39172 34746
rect 39120 34682 39172 34688
rect 38384 21616 38436 21622
rect 38384 21558 38436 21564
rect 38200 21548 38252 21554
rect 38200 21490 38252 21496
rect 38212 20942 38240 21490
rect 38396 21418 38424 21558
rect 38844 21480 38896 21486
rect 38844 21422 38896 21428
rect 38384 21412 38436 21418
rect 38384 21354 38436 21360
rect 38476 21344 38528 21350
rect 38476 21286 38528 21292
rect 38488 20942 38516 21286
rect 38200 20936 38252 20942
rect 38200 20878 38252 20884
rect 38476 20936 38528 20942
rect 38476 20878 38528 20884
rect 38212 20262 38240 20878
rect 38856 20874 38884 21422
rect 38844 20868 38896 20874
rect 38844 20810 38896 20816
rect 38660 20800 38712 20806
rect 38660 20742 38712 20748
rect 38672 20398 38700 20742
rect 38752 20460 38804 20466
rect 38752 20402 38804 20408
rect 38660 20392 38712 20398
rect 38660 20334 38712 20340
rect 38200 20256 38252 20262
rect 38200 20198 38252 20204
rect 38292 19916 38344 19922
rect 38292 19858 38344 19864
rect 38304 19786 38332 19858
rect 38764 19854 38792 20402
rect 38752 19848 38804 19854
rect 38752 19790 38804 19796
rect 38292 19780 38344 19786
rect 38292 19722 38344 19728
rect 38304 18834 38332 19722
rect 38660 19712 38712 19718
rect 38660 19654 38712 19660
rect 38292 18828 38344 18834
rect 38292 18770 38344 18776
rect 38384 18692 38436 18698
rect 38384 18634 38436 18640
rect 38396 18222 38424 18634
rect 38384 18216 38436 18222
rect 38384 18158 38436 18164
rect 38290 17096 38346 17105
rect 38290 17031 38346 17040
rect 38200 16992 38252 16998
rect 38200 16934 38252 16940
rect 38212 16590 38240 16934
rect 38200 16584 38252 16590
rect 38200 16526 38252 16532
rect 38304 13530 38332 17031
rect 38396 16969 38424 18158
rect 38566 17504 38622 17513
rect 38566 17439 38622 17448
rect 38580 17270 38608 17439
rect 38672 17377 38700 19654
rect 38764 18290 38792 19790
rect 38844 18760 38896 18766
rect 38844 18702 38896 18708
rect 38752 18284 38804 18290
rect 38752 18226 38804 18232
rect 38764 17490 38792 18226
rect 38856 17882 38884 18702
rect 39212 18692 39264 18698
rect 39212 18634 39264 18640
rect 39028 18624 39080 18630
rect 39028 18566 39080 18572
rect 39040 18290 39068 18566
rect 39028 18284 39080 18290
rect 39028 18226 39080 18232
rect 39028 18080 39080 18086
rect 39028 18022 39080 18028
rect 38844 17876 38896 17882
rect 38844 17818 38896 17824
rect 39040 17728 39068 18022
rect 39120 17740 39172 17746
rect 39040 17700 39120 17728
rect 38936 17672 38988 17678
rect 38936 17614 38988 17620
rect 38948 17490 38976 17614
rect 38764 17462 38976 17490
rect 38658 17368 38714 17377
rect 38658 17303 38714 17312
rect 38752 17332 38804 17338
rect 38752 17274 38804 17280
rect 38568 17264 38620 17270
rect 38764 17241 38792 17274
rect 38568 17206 38620 17212
rect 38750 17232 38806 17241
rect 38750 17167 38806 17176
rect 38752 17128 38804 17134
rect 38474 17096 38530 17105
rect 38474 17031 38476 17040
rect 38528 17031 38530 17040
rect 38672 17088 38752 17116
rect 38476 17002 38528 17008
rect 38382 16960 38438 16969
rect 38382 16895 38438 16904
rect 38672 16454 38700 17088
rect 38752 17070 38804 17076
rect 38844 17128 38896 17134
rect 38844 17070 38896 17076
rect 38856 16969 38884 17070
rect 38842 16960 38898 16969
rect 38842 16895 38898 16904
rect 38948 16726 38976 17462
rect 38936 16720 38988 16726
rect 38936 16662 38988 16668
rect 38752 16652 38804 16658
rect 38752 16594 38804 16600
rect 38384 16448 38436 16454
rect 38384 16390 38436 16396
rect 38660 16448 38712 16454
rect 38660 16390 38712 16396
rect 38200 13524 38252 13530
rect 38200 13466 38252 13472
rect 38292 13524 38344 13530
rect 38292 13466 38344 13472
rect 38212 12918 38240 13466
rect 38016 12912 38068 12918
rect 38016 12854 38068 12860
rect 38200 12912 38252 12918
rect 38200 12854 38252 12860
rect 38028 12170 38056 12854
rect 38396 12764 38424 16390
rect 38764 16182 38792 16594
rect 38842 16280 38898 16289
rect 38842 16215 38898 16224
rect 38856 16182 38884 16215
rect 38752 16176 38804 16182
rect 38752 16118 38804 16124
rect 38844 16176 38896 16182
rect 38844 16118 38896 16124
rect 38844 16040 38896 16046
rect 38844 15982 38896 15988
rect 38752 14952 38804 14958
rect 38672 14912 38752 14940
rect 38476 14816 38528 14822
rect 38476 14758 38528 14764
rect 38568 14816 38620 14822
rect 38568 14758 38620 14764
rect 38488 13938 38516 14758
rect 38476 13932 38528 13938
rect 38476 13874 38528 13880
rect 38580 13433 38608 14758
rect 38672 13870 38700 14912
rect 38752 14894 38804 14900
rect 38660 13864 38712 13870
rect 38660 13806 38712 13812
rect 38566 13424 38622 13433
rect 38566 13359 38622 13368
rect 38672 13326 38700 13806
rect 38660 13320 38712 13326
rect 38660 13262 38712 13268
rect 38476 13252 38528 13258
rect 38476 13194 38528 13200
rect 38212 12736 38424 12764
rect 38016 12164 38068 12170
rect 38016 12106 38068 12112
rect 37924 12096 37976 12102
rect 37924 12038 37976 12044
rect 38028 11626 38056 12106
rect 38106 12064 38162 12073
rect 38106 11999 38162 12008
rect 38016 11620 38068 11626
rect 38016 11562 38068 11568
rect 37830 11112 37886 11121
rect 37830 11047 37886 11056
rect 37740 10600 37792 10606
rect 37740 10542 37792 10548
rect 37752 10198 37780 10542
rect 37740 10192 37792 10198
rect 37740 10134 37792 10140
rect 37752 9994 37780 10134
rect 37740 9988 37792 9994
rect 37740 9930 37792 9936
rect 37844 9586 37872 11047
rect 38016 10600 38068 10606
rect 38016 10542 38068 10548
rect 37832 9580 37884 9586
rect 37832 9522 37884 9528
rect 38028 9466 38056 10542
rect 38120 10470 38148 11999
rect 38108 10464 38160 10470
rect 38108 10406 38160 10412
rect 38120 9586 38148 10406
rect 38108 9580 38160 9586
rect 38108 9522 38160 9528
rect 37752 9438 38056 9466
rect 37752 8974 37780 9438
rect 37740 8968 37792 8974
rect 37740 8910 37792 8916
rect 38016 8900 38068 8906
rect 38016 8842 38068 8848
rect 37648 8560 37700 8566
rect 37648 8502 37700 8508
rect 37280 8492 37332 8498
rect 37280 8434 37332 8440
rect 37556 8492 37608 8498
rect 37556 8434 37608 8440
rect 37292 8106 37320 8434
rect 38028 8430 38056 8842
rect 38016 8424 38068 8430
rect 37462 8392 37518 8401
rect 38016 8366 38068 8372
rect 37462 8327 37518 8336
rect 37292 8078 37412 8106
rect 37280 8016 37332 8022
rect 37280 7958 37332 7964
rect 37292 7274 37320 7958
rect 37280 7268 37332 7274
rect 37280 7210 37332 7216
rect 37188 6860 37240 6866
rect 37188 6802 37240 6808
rect 37280 6316 37332 6322
rect 37280 6258 37332 6264
rect 37188 5228 37240 5234
rect 37188 5170 37240 5176
rect 37200 4554 37228 5170
rect 37188 4548 37240 4554
rect 37188 4490 37240 4496
rect 37200 4146 37228 4490
rect 37188 4140 37240 4146
rect 37188 4082 37240 4088
rect 37188 3732 37240 3738
rect 37188 3674 37240 3680
rect 37096 3188 37148 3194
rect 37096 3130 37148 3136
rect 37200 2774 37228 3674
rect 37292 2961 37320 6258
rect 37384 5710 37412 8078
rect 37372 5704 37424 5710
rect 37372 5646 37424 5652
rect 37384 5234 37412 5646
rect 37372 5228 37424 5234
rect 37372 5170 37424 5176
rect 37372 4684 37424 4690
rect 37372 4626 37424 4632
rect 37384 4214 37412 4626
rect 37476 4486 37504 8327
rect 38212 8294 38240 12736
rect 38384 11144 38436 11150
rect 38304 11104 38384 11132
rect 38304 9874 38332 11104
rect 38384 11086 38436 11092
rect 38384 10056 38436 10062
rect 38488 10044 38516 13194
rect 38672 11082 38700 13262
rect 38752 11756 38804 11762
rect 38752 11698 38804 11704
rect 38660 11076 38712 11082
rect 38660 11018 38712 11024
rect 38672 10606 38700 11018
rect 38764 10606 38792 11698
rect 38660 10600 38712 10606
rect 38660 10542 38712 10548
rect 38752 10600 38804 10606
rect 38752 10542 38804 10548
rect 38750 10296 38806 10305
rect 38750 10231 38752 10240
rect 38804 10231 38806 10240
rect 38752 10202 38804 10208
rect 38614 10192 38666 10198
rect 38666 10160 38714 10169
rect 38614 10134 38658 10140
rect 38626 10118 38658 10134
rect 38658 10095 38714 10104
rect 38436 10016 38516 10044
rect 38568 10056 38620 10062
rect 38384 9998 38436 10004
rect 38620 10016 38700 10044
rect 38856 10033 38884 15982
rect 38936 15156 38988 15162
rect 38936 15098 38988 15104
rect 38948 14074 38976 15098
rect 38936 14068 38988 14074
rect 38936 14010 38988 14016
rect 38948 13462 38976 14010
rect 38936 13456 38988 13462
rect 38936 13398 38988 13404
rect 39040 12753 39068 17700
rect 39120 17682 39172 17688
rect 39120 17536 39172 17542
rect 39120 17478 39172 17484
rect 39132 16998 39160 17478
rect 39120 16992 39172 16998
rect 39120 16934 39172 16940
rect 39120 14340 39172 14346
rect 39120 14282 39172 14288
rect 39132 14074 39160 14282
rect 39120 14068 39172 14074
rect 39120 14010 39172 14016
rect 39224 12832 39252 18634
rect 39304 17060 39356 17066
rect 39304 17002 39356 17008
rect 39316 13258 39344 17002
rect 39304 13252 39356 13258
rect 39304 13194 39356 13200
rect 39132 12804 39252 12832
rect 39026 12744 39082 12753
rect 39026 12679 39082 12688
rect 38936 11756 38988 11762
rect 38936 11698 38988 11704
rect 38948 11218 38976 11698
rect 38936 11212 38988 11218
rect 38936 11154 38988 11160
rect 38568 9998 38620 10004
rect 38568 9920 38620 9926
rect 38304 9846 38516 9874
rect 38672 9897 38700 10016
rect 38842 10024 38898 10033
rect 38842 9959 38898 9968
rect 38568 9862 38620 9868
rect 38658 9888 38714 9897
rect 38384 9716 38436 9722
rect 38384 9658 38436 9664
rect 38396 9217 38424 9658
rect 38382 9208 38438 9217
rect 38382 9143 38438 9152
rect 38488 8974 38516 9846
rect 38580 9586 38608 9862
rect 38658 9823 38714 9832
rect 38750 9752 38806 9761
rect 38856 9738 38884 9959
rect 38750 9687 38806 9696
rect 38847 9710 38884 9738
rect 38764 9625 38792 9687
rect 38750 9616 38806 9625
rect 38568 9580 38620 9586
rect 38568 9522 38620 9528
rect 38660 9580 38712 9586
rect 38847 9602 38875 9710
rect 38847 9586 38884 9602
rect 38750 9551 38806 9560
rect 38844 9580 38896 9586
rect 38660 9522 38712 9528
rect 38844 9522 38896 9528
rect 38566 9072 38622 9081
rect 38566 9007 38568 9016
rect 38620 9007 38622 9016
rect 38568 8978 38620 8984
rect 38476 8968 38528 8974
rect 38476 8910 38528 8916
rect 38384 8832 38436 8838
rect 38384 8774 38436 8780
rect 38290 8664 38346 8673
rect 38290 8599 38346 8608
rect 37936 8266 38240 8294
rect 37740 8084 37792 8090
rect 37740 8026 37792 8032
rect 37752 7750 37780 8026
rect 37740 7744 37792 7750
rect 37740 7686 37792 7692
rect 37648 5840 37700 5846
rect 37648 5782 37700 5788
rect 37556 5568 37608 5574
rect 37556 5510 37608 5516
rect 37464 4480 37516 4486
rect 37464 4422 37516 4428
rect 37372 4208 37424 4214
rect 37372 4150 37424 4156
rect 37370 3904 37426 3913
rect 37370 3839 37426 3848
rect 37384 3534 37412 3839
rect 37568 3534 37596 5510
rect 37660 5234 37688 5782
rect 37740 5704 37792 5710
rect 37740 5646 37792 5652
rect 37648 5228 37700 5234
rect 37648 5170 37700 5176
rect 37648 4208 37700 4214
rect 37648 4150 37700 4156
rect 37372 3528 37424 3534
rect 37372 3470 37424 3476
rect 37556 3528 37608 3534
rect 37556 3470 37608 3476
rect 37370 3088 37426 3097
rect 37370 3023 37426 3032
rect 37278 2952 37334 2961
rect 37278 2887 37334 2896
rect 37108 2746 37228 2774
rect 37004 2032 37056 2038
rect 37004 1974 37056 1980
rect 36912 1896 36964 1902
rect 36912 1838 36964 1844
rect 36924 1698 36952 1838
rect 36912 1692 36964 1698
rect 36912 1634 36964 1640
rect 36728 1556 36780 1562
rect 36728 1498 36780 1504
rect 36820 1352 36872 1358
rect 36820 1294 36872 1300
rect 36832 800 36860 1294
rect 37108 800 37136 2746
rect 37384 800 37412 3023
rect 37464 2916 37516 2922
rect 37464 2858 37516 2864
rect 37476 1426 37504 2858
rect 37464 1420 37516 1426
rect 37464 1362 37516 1368
rect 37660 800 37688 4150
rect 37752 3194 37780 5646
rect 37832 5024 37884 5030
rect 37832 4966 37884 4972
rect 37844 4622 37872 4966
rect 37936 4690 37964 8266
rect 38106 6216 38162 6225
rect 38106 6151 38162 6160
rect 38016 5636 38068 5642
rect 38016 5578 38068 5584
rect 37924 4684 37976 4690
rect 37924 4626 37976 4632
rect 37832 4616 37884 4622
rect 37832 4558 37884 4564
rect 37832 3936 37884 3942
rect 37832 3878 37884 3884
rect 37740 3188 37792 3194
rect 37740 3130 37792 3136
rect 37844 1358 37872 3878
rect 38028 2774 38056 5578
rect 38120 2990 38148 6151
rect 38200 4548 38252 4554
rect 38200 4490 38252 4496
rect 38108 2984 38160 2990
rect 38108 2926 38160 2932
rect 37936 2746 38056 2774
rect 37936 2446 37964 2746
rect 37924 2440 37976 2446
rect 37924 2382 37976 2388
rect 37924 1692 37976 1698
rect 37924 1634 37976 1640
rect 37832 1352 37884 1358
rect 37832 1294 37884 1300
rect 37936 800 37964 1634
rect 38212 800 38240 4490
rect 38304 3670 38332 8599
rect 38396 7954 38424 8774
rect 38488 8537 38516 8910
rect 38474 8528 38530 8537
rect 38474 8463 38530 8472
rect 38672 8129 38700 9522
rect 38844 9444 38896 9450
rect 38844 9386 38896 9392
rect 38856 8922 38884 9386
rect 38936 9172 38988 9178
rect 38936 9114 38988 9120
rect 38764 8894 38884 8922
rect 38658 8120 38714 8129
rect 38658 8055 38714 8064
rect 38658 7984 38714 7993
rect 38384 7948 38436 7954
rect 38658 7919 38660 7928
rect 38384 7890 38436 7896
rect 38712 7919 38714 7928
rect 38660 7890 38712 7896
rect 38660 7812 38712 7818
rect 38660 7754 38712 7760
rect 38568 7540 38620 7546
rect 38568 7482 38620 7488
rect 38580 7342 38608 7482
rect 38568 7336 38620 7342
rect 38568 7278 38620 7284
rect 38382 6488 38438 6497
rect 38382 6423 38438 6432
rect 38396 5846 38424 6423
rect 38384 5840 38436 5846
rect 38384 5782 38436 5788
rect 38580 5778 38608 7278
rect 38672 6866 38700 7754
rect 38660 6860 38712 6866
rect 38660 6802 38712 6808
rect 38568 5772 38620 5778
rect 38568 5714 38620 5720
rect 38476 5092 38528 5098
rect 38476 5034 38528 5040
rect 38292 3664 38344 3670
rect 38344 3624 38424 3652
rect 38292 3606 38344 3612
rect 38292 3460 38344 3466
rect 38292 3402 38344 3408
rect 38304 3097 38332 3402
rect 38396 3194 38424 3624
rect 38384 3188 38436 3194
rect 38384 3130 38436 3136
rect 38290 3088 38346 3097
rect 38290 3023 38346 3032
rect 38488 800 38516 5034
rect 38764 4554 38792 8894
rect 38844 8288 38896 8294
rect 38844 8230 38896 8236
rect 38856 8022 38884 8230
rect 38948 8022 38976 9114
rect 38844 8016 38896 8022
rect 38844 7958 38896 7964
rect 38936 8016 38988 8022
rect 38936 7958 38988 7964
rect 38835 7846 38887 7852
rect 38835 7788 38887 7794
rect 38856 5642 38884 7788
rect 38844 5636 38896 5642
rect 38844 5578 38896 5584
rect 38936 5568 38988 5574
rect 38936 5510 38988 5516
rect 38948 5234 38976 5510
rect 38936 5228 38988 5234
rect 38936 5170 38988 5176
rect 38844 5024 38896 5030
rect 38844 4966 38896 4972
rect 38752 4548 38804 4554
rect 38752 4490 38804 4496
rect 38856 4146 38884 4966
rect 39040 4690 39068 12679
rect 39132 11830 39160 12804
rect 39210 12608 39266 12617
rect 39210 12543 39266 12552
rect 39120 11824 39172 11830
rect 39120 11766 39172 11772
rect 39120 10600 39172 10606
rect 39120 10542 39172 10548
rect 39132 9761 39160 10542
rect 39118 9752 39174 9761
rect 39118 9687 39174 9696
rect 39224 9654 39252 12543
rect 39408 10962 39436 54470
rect 39488 50380 39540 50386
rect 39488 50322 39540 50328
rect 39500 17066 39528 50322
rect 40132 47660 40184 47666
rect 40132 47602 40184 47608
rect 39580 38412 39632 38418
rect 39580 38354 39632 38360
rect 39488 17060 39540 17066
rect 39488 17002 39540 17008
rect 39488 16720 39540 16726
rect 39488 16662 39540 16668
rect 39500 16250 39528 16662
rect 39488 16244 39540 16250
rect 39488 16186 39540 16192
rect 39488 14884 39540 14890
rect 39488 14826 39540 14832
rect 39500 14618 39528 14826
rect 39488 14612 39540 14618
rect 39488 14554 39540 14560
rect 39500 14006 39528 14554
rect 39488 14000 39540 14006
rect 39488 13942 39540 13948
rect 39408 10934 39528 10962
rect 39396 10804 39448 10810
rect 39396 10746 39448 10752
rect 39408 9994 39436 10746
rect 39396 9988 39448 9994
rect 39396 9930 39448 9936
rect 39212 9648 39264 9654
rect 39212 9590 39264 9596
rect 39304 9444 39356 9450
rect 39304 9386 39356 9392
rect 39316 9042 39344 9386
rect 39304 9036 39356 9042
rect 39304 8978 39356 8984
rect 39394 8936 39450 8945
rect 39394 8871 39450 8880
rect 39212 8492 39264 8498
rect 39212 8434 39264 8440
rect 39120 8424 39172 8430
rect 39120 8366 39172 8372
rect 39028 4684 39080 4690
rect 39028 4626 39080 4632
rect 38844 4140 38896 4146
rect 38844 4082 38896 4088
rect 38568 3392 38620 3398
rect 38566 3360 38568 3369
rect 38620 3360 38622 3369
rect 38566 3295 38622 3304
rect 38844 3188 38896 3194
rect 38844 3130 38896 3136
rect 38568 2984 38620 2990
rect 38568 2926 38620 2932
rect 38580 1222 38608 2926
rect 38568 1216 38620 1222
rect 38856 1170 38884 3130
rect 38936 3052 38988 3058
rect 39040 3040 39068 4626
rect 39132 3602 39160 8366
rect 39224 8090 39252 8434
rect 39212 8084 39264 8090
rect 39212 8026 39264 8032
rect 39210 7984 39266 7993
rect 39408 7954 39436 8871
rect 39210 7919 39266 7928
rect 39396 7948 39448 7954
rect 39224 7886 39252 7919
rect 39396 7890 39448 7896
rect 39212 7880 39264 7886
rect 39212 7822 39264 7828
rect 39304 6112 39356 6118
rect 39304 6054 39356 6060
rect 39212 5024 39264 5030
rect 39212 4966 39264 4972
rect 39224 4486 39252 4966
rect 39212 4480 39264 4486
rect 39212 4422 39264 4428
rect 39120 3596 39172 3602
rect 39120 3538 39172 3544
rect 39316 3058 39344 6054
rect 39500 4690 39528 10934
rect 39592 6905 39620 38354
rect 39672 23044 39724 23050
rect 39672 22986 39724 22992
rect 39684 22094 39712 22986
rect 39684 22066 39896 22094
rect 39672 20324 39724 20330
rect 39672 20266 39724 20272
rect 39684 19990 39712 20266
rect 39764 20256 39816 20262
rect 39764 20198 39816 20204
rect 39672 19984 39724 19990
rect 39672 19926 39724 19932
rect 39776 19718 39804 20198
rect 39764 19712 39816 19718
rect 39764 19654 39816 19660
rect 39672 17536 39724 17542
rect 39670 17504 39672 17513
rect 39724 17504 39726 17513
rect 39670 17439 39726 17448
rect 39684 16794 39712 17439
rect 39762 17096 39818 17105
rect 39762 17031 39764 17040
rect 39816 17031 39818 17040
rect 39764 17002 39816 17008
rect 39672 16788 39724 16794
rect 39672 16730 39724 16736
rect 39764 16108 39816 16114
rect 39764 16050 39816 16056
rect 39672 7948 39724 7954
rect 39672 7890 39724 7896
rect 39684 7750 39712 7890
rect 39672 7744 39724 7750
rect 39672 7686 39724 7692
rect 39578 6896 39634 6905
rect 39578 6831 39634 6840
rect 39672 5228 39724 5234
rect 39672 5170 39724 5176
rect 39488 4684 39540 4690
rect 39488 4626 39540 4632
rect 39684 3738 39712 5170
rect 39672 3732 39724 3738
rect 39672 3674 39724 3680
rect 38988 3012 39068 3040
rect 39304 3052 39356 3058
rect 38936 2994 38988 3000
rect 39304 2994 39356 3000
rect 39580 3052 39632 3058
rect 39580 2994 39632 3000
rect 39304 2372 39356 2378
rect 39304 2314 39356 2320
rect 38568 1158 38620 1164
rect 38764 1142 38884 1170
rect 38764 800 38792 1142
rect 39028 1080 39080 1086
rect 39028 1022 39080 1028
rect 39040 800 39068 1022
rect 39316 800 39344 2314
rect 39592 800 39620 2994
rect 39776 1970 39804 16050
rect 39868 11558 39896 22066
rect 39948 20596 40000 20602
rect 39948 20538 40000 20544
rect 39960 19378 39988 20538
rect 39948 19372 40000 19378
rect 39948 19314 40000 19320
rect 40038 18864 40094 18873
rect 40038 18799 40040 18808
rect 40092 18799 40094 18808
rect 40040 18770 40092 18776
rect 40040 18080 40092 18086
rect 40040 18022 40092 18028
rect 40052 16998 40080 18022
rect 40040 16992 40092 16998
rect 40040 16934 40092 16940
rect 40144 16182 40172 47602
rect 40328 35086 40356 60998
rect 41340 60874 41368 63200
rect 41880 61600 41932 61606
rect 41880 61542 41932 61548
rect 41512 61260 41564 61266
rect 41512 61202 41564 61208
rect 41340 60846 41460 60874
rect 41432 60790 41460 60846
rect 41420 60784 41472 60790
rect 41420 60726 41472 60732
rect 40776 60648 40828 60654
rect 40776 60590 40828 60596
rect 40592 60104 40644 60110
rect 40592 60046 40644 60052
rect 40604 59498 40632 60046
rect 40788 60042 40816 60590
rect 40868 60512 40920 60518
rect 40868 60454 40920 60460
rect 40880 60110 40908 60454
rect 41144 60240 41196 60246
rect 41144 60182 41196 60188
rect 40868 60104 40920 60110
rect 40868 60046 40920 60052
rect 40960 60104 41012 60110
rect 40960 60046 41012 60052
rect 40776 60036 40828 60042
rect 40776 59978 40828 59984
rect 40592 59492 40644 59498
rect 40592 59434 40644 59440
rect 40972 58478 41000 60046
rect 40960 58472 41012 58478
rect 40960 58414 41012 58420
rect 40972 56302 41000 58414
rect 40960 56296 41012 56302
rect 40960 56238 41012 56244
rect 40868 55888 40920 55894
rect 40868 55830 40920 55836
rect 40500 55344 40552 55350
rect 40500 55286 40552 55292
rect 40512 53514 40540 55286
rect 40880 55282 40908 55830
rect 40972 55282 41000 56238
rect 40868 55276 40920 55282
rect 40868 55218 40920 55224
rect 40960 55276 41012 55282
rect 40960 55218 41012 55224
rect 40868 53712 40920 53718
rect 40868 53654 40920 53660
rect 40500 53508 40552 53514
rect 40500 53450 40552 53456
rect 40880 51074 40908 53654
rect 41156 51474 41184 60182
rect 41524 60178 41552 61202
rect 41696 61056 41748 61062
rect 41696 60998 41748 61004
rect 41512 60172 41564 60178
rect 41512 60114 41564 60120
rect 41236 59016 41288 59022
rect 41236 58958 41288 58964
rect 41248 56438 41276 58958
rect 41512 58540 41564 58546
rect 41512 58482 41564 58488
rect 41328 58336 41380 58342
rect 41328 58278 41380 58284
rect 41340 56846 41368 58278
rect 41524 58138 41552 58482
rect 41512 58132 41564 58138
rect 41512 58074 41564 58080
rect 41328 56840 41380 56846
rect 41328 56782 41380 56788
rect 41236 56432 41288 56438
rect 41236 56374 41288 56380
rect 41248 55418 41276 56374
rect 41328 56160 41380 56166
rect 41328 56102 41380 56108
rect 41236 55412 41288 55418
rect 41236 55354 41288 55360
rect 41236 55276 41288 55282
rect 41236 55218 41288 55224
rect 41248 53582 41276 55218
rect 41340 55214 41368 56102
rect 41340 55186 41644 55214
rect 41236 53576 41288 53582
rect 41236 53518 41288 53524
rect 41144 51468 41196 51474
rect 41144 51410 41196 51416
rect 40880 51046 41092 51074
rect 40592 35692 40644 35698
rect 40592 35634 40644 35640
rect 40408 35624 40460 35630
rect 40408 35566 40460 35572
rect 40420 35442 40448 35566
rect 40604 35562 40632 35634
rect 40592 35556 40644 35562
rect 40592 35498 40644 35504
rect 40420 35414 40724 35442
rect 40696 35290 40724 35414
rect 40684 35284 40736 35290
rect 40684 35226 40736 35232
rect 40500 35148 40552 35154
rect 40500 35090 40552 35096
rect 40316 35080 40368 35086
rect 40316 35022 40368 35028
rect 40408 35080 40460 35086
rect 40408 35022 40460 35028
rect 40420 34474 40448 35022
rect 40408 34468 40460 34474
rect 40408 34410 40460 34416
rect 40420 33658 40448 34410
rect 40408 33652 40460 33658
rect 40408 33594 40460 33600
rect 40408 33448 40460 33454
rect 40408 33390 40460 33396
rect 40316 25764 40368 25770
rect 40316 25706 40368 25712
rect 40224 20256 40276 20262
rect 40224 20198 40276 20204
rect 40236 19786 40264 20198
rect 40224 19780 40276 19786
rect 40224 19722 40276 19728
rect 40328 17270 40356 25706
rect 40316 17264 40368 17270
rect 40316 17206 40368 17212
rect 40132 16176 40184 16182
rect 40132 16118 40184 16124
rect 40038 15600 40094 15609
rect 40038 15535 40094 15544
rect 39948 14408 40000 14414
rect 39948 14350 40000 14356
rect 39856 11552 39908 11558
rect 39856 11494 39908 11500
rect 39856 11280 39908 11286
rect 39856 11222 39908 11228
rect 39868 4078 39896 11222
rect 39960 11150 39988 14350
rect 40052 12238 40080 15535
rect 40132 15428 40184 15434
rect 40132 15370 40184 15376
rect 40144 12434 40172 15370
rect 40316 15020 40368 15026
rect 40316 14962 40368 14968
rect 40328 14618 40356 14962
rect 40224 14612 40276 14618
rect 40224 14554 40276 14560
rect 40316 14612 40368 14618
rect 40316 14554 40368 14560
rect 40236 14498 40264 14554
rect 40236 14470 40356 14498
rect 40144 12406 40264 12434
rect 40040 12232 40092 12238
rect 40040 12174 40092 12180
rect 40132 12232 40184 12238
rect 40132 12174 40184 12180
rect 40052 11393 40080 12174
rect 40144 11801 40172 12174
rect 40130 11792 40186 11801
rect 40130 11727 40186 11736
rect 40236 11676 40264 12406
rect 40144 11648 40264 11676
rect 40038 11384 40094 11393
rect 40038 11319 40094 11328
rect 39948 11144 40000 11150
rect 39948 11086 40000 11092
rect 39960 8566 39988 11086
rect 40040 9104 40092 9110
rect 40040 9046 40092 9052
rect 39948 8560 40000 8566
rect 39948 8502 40000 8508
rect 40052 7886 40080 9046
rect 40040 7880 40092 7886
rect 40040 7822 40092 7828
rect 40144 7342 40172 11648
rect 40328 9926 40356 14470
rect 40316 9920 40368 9926
rect 40316 9862 40368 9868
rect 40316 9376 40368 9382
rect 40316 9318 40368 9324
rect 40224 8968 40276 8974
rect 40222 8936 40224 8945
rect 40276 8936 40278 8945
rect 40222 8871 40278 8880
rect 40132 7336 40184 7342
rect 40132 7278 40184 7284
rect 40040 5636 40092 5642
rect 40040 5578 40092 5584
rect 39948 5568 40000 5574
rect 39948 5510 40000 5516
rect 39856 4072 39908 4078
rect 39856 4014 39908 4020
rect 39960 4010 39988 5510
rect 39948 4004 40000 4010
rect 39948 3946 40000 3952
rect 39960 3913 39988 3946
rect 39946 3904 40002 3913
rect 39946 3839 40002 3848
rect 40052 2774 40080 5578
rect 40224 5296 40276 5302
rect 40224 5238 40276 5244
rect 40236 5098 40264 5238
rect 40224 5092 40276 5098
rect 40224 5034 40276 5040
rect 40328 4758 40356 9318
rect 40316 4752 40368 4758
rect 40316 4694 40368 4700
rect 40132 4548 40184 4554
rect 40132 4490 40184 4496
rect 40144 4146 40172 4490
rect 40316 4480 40368 4486
rect 40236 4440 40316 4468
rect 40132 4140 40184 4146
rect 40132 4082 40184 4088
rect 40130 4040 40186 4049
rect 40130 3975 40186 3984
rect 40144 3602 40172 3975
rect 40132 3596 40184 3602
rect 40132 3538 40184 3544
rect 40236 3126 40264 4440
rect 40316 4422 40368 4428
rect 40420 3126 40448 33390
rect 40512 5846 40540 35090
rect 41064 22094 41092 51046
rect 41616 26234 41644 55186
rect 41708 35630 41736 60998
rect 41788 59084 41840 59090
rect 41788 59026 41840 59032
rect 41800 58478 41828 59026
rect 41892 59022 41920 61542
rect 42076 61198 42104 63200
rect 42708 61736 42760 61742
rect 42708 61678 42760 61684
rect 42616 61396 42668 61402
rect 42616 61338 42668 61344
rect 42064 61192 42116 61198
rect 42064 61134 42116 61140
rect 42156 60104 42208 60110
rect 42156 60046 42208 60052
rect 42340 60104 42392 60110
rect 42340 60046 42392 60052
rect 41972 59968 42024 59974
rect 41972 59910 42024 59916
rect 41984 59401 42012 59910
rect 42168 59634 42196 60046
rect 42352 59770 42380 60046
rect 42340 59764 42392 59770
rect 42340 59706 42392 59712
rect 42352 59634 42380 59706
rect 42156 59628 42208 59634
rect 42156 59570 42208 59576
rect 42340 59628 42392 59634
rect 42340 59570 42392 59576
rect 41970 59392 42026 59401
rect 41970 59327 42026 59336
rect 41880 59016 41932 59022
rect 41880 58958 41932 58964
rect 42340 58880 42392 58886
rect 42340 58822 42392 58828
rect 41788 58472 41840 58478
rect 41788 58414 41840 58420
rect 42064 55276 42116 55282
rect 42064 55218 42116 55224
rect 41788 50448 41840 50454
rect 41788 50390 41840 50396
rect 41696 35624 41748 35630
rect 41696 35566 41748 35572
rect 41696 27124 41748 27130
rect 41696 27066 41748 27072
rect 40880 22066 41092 22094
rect 41524 26206 41644 26234
rect 40776 19372 40828 19378
rect 40776 19314 40828 19320
rect 40592 18624 40644 18630
rect 40592 18566 40644 18572
rect 40604 17678 40632 18566
rect 40592 17672 40644 17678
rect 40592 17614 40644 17620
rect 40684 17264 40736 17270
rect 40684 17206 40736 17212
rect 40592 16108 40644 16114
rect 40592 16050 40644 16056
rect 40604 15366 40632 16050
rect 40592 15360 40644 15366
rect 40592 15302 40644 15308
rect 40604 12238 40632 15302
rect 40592 12232 40644 12238
rect 40592 12174 40644 12180
rect 40604 11830 40632 12174
rect 40592 11824 40644 11830
rect 40592 11766 40644 11772
rect 40604 9586 40632 11766
rect 40592 9580 40644 9586
rect 40592 9522 40644 9528
rect 40500 5840 40552 5846
rect 40500 5782 40552 5788
rect 40696 5370 40724 17206
rect 40788 12442 40816 19314
rect 40880 16590 40908 22066
rect 41144 20936 41196 20942
rect 41144 20878 41196 20884
rect 41156 20398 41184 20878
rect 41420 20800 41472 20806
rect 41420 20742 41472 20748
rect 41432 20466 41460 20742
rect 41420 20460 41472 20466
rect 41420 20402 41472 20408
rect 41144 20392 41196 20398
rect 41144 20334 41196 20340
rect 41156 18873 41184 20334
rect 41524 19122 41552 26206
rect 41708 22094 41736 27066
rect 41616 22066 41736 22094
rect 41616 20890 41644 22066
rect 41696 21480 41748 21486
rect 41696 21422 41748 21428
rect 41708 21010 41736 21422
rect 41696 21004 41748 21010
rect 41696 20946 41748 20952
rect 41616 20862 41736 20890
rect 41604 20256 41656 20262
rect 41604 20198 41656 20204
rect 41616 19786 41644 20198
rect 41604 19780 41656 19786
rect 41604 19722 41656 19728
rect 41524 19094 41644 19122
rect 41142 18864 41198 18873
rect 41142 18799 41198 18808
rect 40960 18624 41012 18630
rect 40958 18592 40960 18601
rect 41012 18592 41014 18601
rect 40958 18527 41014 18536
rect 40972 18426 41000 18527
rect 40960 18420 41012 18426
rect 40960 18362 41012 18368
rect 40960 18080 41012 18086
rect 40960 18022 41012 18028
rect 40972 17270 41000 18022
rect 40960 17264 41012 17270
rect 40960 17206 41012 17212
rect 41052 17264 41104 17270
rect 41052 17206 41104 17212
rect 41064 16674 41092 17206
rect 40972 16646 41092 16674
rect 40868 16584 40920 16590
rect 40868 16526 40920 16532
rect 40868 16448 40920 16454
rect 40868 16390 40920 16396
rect 40880 12986 40908 16390
rect 40972 15910 41000 16646
rect 41052 16584 41104 16590
rect 41052 16526 41104 16532
rect 41064 16250 41092 16526
rect 41052 16244 41104 16250
rect 41052 16186 41104 16192
rect 40960 15904 41012 15910
rect 40958 15872 40960 15881
rect 41012 15872 41014 15881
rect 40958 15807 41014 15816
rect 41050 15600 41106 15609
rect 41050 15535 41106 15544
rect 41064 15502 41092 15535
rect 41052 15496 41104 15502
rect 41052 15438 41104 15444
rect 41156 14958 41184 18799
rect 41328 17264 41380 17270
rect 41326 17232 41328 17241
rect 41380 17232 41382 17241
rect 41326 17167 41382 17176
rect 41236 16516 41288 16522
rect 41236 16458 41288 16464
rect 41328 16516 41380 16522
rect 41328 16458 41380 16464
rect 41420 16516 41472 16522
rect 41420 16458 41472 16464
rect 41248 15502 41276 16458
rect 41340 15706 41368 16458
rect 41328 15700 41380 15706
rect 41328 15642 41380 15648
rect 41432 15570 41460 16458
rect 41616 16046 41644 19094
rect 41708 18170 41736 20862
rect 41800 18358 41828 50390
rect 41972 22432 42024 22438
rect 41972 22374 42024 22380
rect 41984 20806 42012 22374
rect 41972 20800 42024 20806
rect 41972 20742 42024 20748
rect 41880 19168 41932 19174
rect 41878 19136 41880 19145
rect 41932 19136 41934 19145
rect 41878 19071 41934 19080
rect 41880 18624 41932 18630
rect 41880 18566 41932 18572
rect 41788 18352 41840 18358
rect 41788 18294 41840 18300
rect 41708 18142 41828 18170
rect 41696 16108 41748 16114
rect 41696 16050 41748 16056
rect 41604 16040 41656 16046
rect 41604 15982 41656 15988
rect 41708 15706 41736 16050
rect 41696 15700 41748 15706
rect 41696 15642 41748 15648
rect 41420 15564 41472 15570
rect 41420 15506 41472 15512
rect 41236 15496 41288 15502
rect 41236 15438 41288 15444
rect 41144 14952 41196 14958
rect 41144 14894 41196 14900
rect 41052 14816 41104 14822
rect 41052 14758 41104 14764
rect 41064 14482 41092 14758
rect 41052 14476 41104 14482
rect 41052 14418 41104 14424
rect 40868 12980 40920 12986
rect 40868 12922 40920 12928
rect 41144 12776 41196 12782
rect 41144 12718 41196 12724
rect 40776 12436 40828 12442
rect 40776 12378 40828 12384
rect 41156 11540 41184 12718
rect 41248 12374 41276 15438
rect 41800 15434 41828 18142
rect 41892 17542 41920 18566
rect 41880 17536 41932 17542
rect 41880 17478 41932 17484
rect 41788 15428 41840 15434
rect 41788 15370 41840 15376
rect 41604 14816 41656 14822
rect 41604 14758 41656 14764
rect 41616 14006 41644 14758
rect 41788 14272 41840 14278
rect 41788 14214 41840 14220
rect 41604 14000 41656 14006
rect 41604 13942 41656 13948
rect 41512 13932 41564 13938
rect 41512 13874 41564 13880
rect 41696 13932 41748 13938
rect 41696 13874 41748 13880
rect 41420 13320 41472 13326
rect 41420 13262 41472 13268
rect 41236 12368 41288 12374
rect 41236 12310 41288 12316
rect 41248 12238 41276 12310
rect 41236 12232 41288 12238
rect 41236 12174 41288 12180
rect 41432 12170 41460 13262
rect 41420 12164 41472 12170
rect 41420 12106 41472 12112
rect 41432 11694 41460 12106
rect 41524 11694 41552 13874
rect 41604 13388 41656 13394
rect 41604 13330 41656 13336
rect 41236 11688 41288 11694
rect 41420 11688 41472 11694
rect 41288 11648 41368 11676
rect 41236 11630 41288 11636
rect 41156 11512 41276 11540
rect 41144 11076 41196 11082
rect 41144 11018 41196 11024
rect 40960 11008 41012 11014
rect 40960 10950 41012 10956
rect 40972 10146 41000 10950
rect 41156 10810 41184 11018
rect 41144 10804 41196 10810
rect 41144 10746 41196 10752
rect 40972 10118 41184 10146
rect 41248 10130 41276 11512
rect 41340 11354 41368 11648
rect 41420 11630 41472 11636
rect 41512 11688 41564 11694
rect 41512 11630 41564 11636
rect 41328 11348 41380 11354
rect 41328 11290 41380 11296
rect 41418 11248 41474 11257
rect 41418 11183 41474 11192
rect 41052 10056 41104 10062
rect 41052 9998 41104 10004
rect 40776 9920 40828 9926
rect 40776 9862 40828 9868
rect 40788 9586 40816 9862
rect 40776 9580 40828 9586
rect 40776 9522 40828 9528
rect 40868 8968 40920 8974
rect 40868 8910 40920 8916
rect 40880 8362 40908 8910
rect 40960 8832 41012 8838
rect 40960 8774 41012 8780
rect 40972 8634 41000 8774
rect 40960 8628 41012 8634
rect 40960 8570 41012 8576
rect 40868 8356 40920 8362
rect 40868 8298 40920 8304
rect 40684 5364 40736 5370
rect 40684 5306 40736 5312
rect 40500 5228 40552 5234
rect 40500 5170 40552 5176
rect 40224 3120 40276 3126
rect 40224 3062 40276 3068
rect 40408 3120 40460 3126
rect 40408 3062 40460 3068
rect 40512 2774 40540 5170
rect 40682 5128 40738 5137
rect 40682 5063 40738 5072
rect 40696 5030 40724 5063
rect 40684 5024 40736 5030
rect 40684 4966 40736 4972
rect 40776 4820 40828 4826
rect 40776 4762 40828 4768
rect 40788 4554 40816 4762
rect 40960 4616 41012 4622
rect 40960 4558 41012 4564
rect 40776 4548 40828 4554
rect 40776 4490 40828 4496
rect 40592 4140 40644 4146
rect 40592 4082 40644 4088
rect 40604 3398 40632 4082
rect 40788 3670 40816 4490
rect 40776 3664 40828 3670
rect 40776 3606 40828 3612
rect 40868 3596 40920 3602
rect 40868 3538 40920 3544
rect 40592 3392 40644 3398
rect 40592 3334 40644 3340
rect 40684 3188 40736 3194
rect 40684 3130 40736 3136
rect 39868 2746 40080 2774
rect 40420 2746 40540 2774
rect 39764 1964 39816 1970
rect 39764 1906 39816 1912
rect 39868 800 39896 2746
rect 40224 2440 40276 2446
rect 40224 2382 40276 2388
rect 40236 1170 40264 2382
rect 40144 1142 40264 1170
rect 40144 800 40172 1142
rect 40420 800 40448 2746
rect 40696 800 40724 3130
rect 40880 2650 40908 3538
rect 40972 3534 41000 4558
rect 40960 3528 41012 3534
rect 40960 3470 41012 3476
rect 40960 2916 41012 2922
rect 40960 2858 41012 2864
rect 40868 2644 40920 2650
rect 40868 2586 40920 2592
rect 40972 800 41000 2858
rect 41064 2106 41092 9998
rect 41156 5114 41184 10118
rect 41236 10124 41288 10130
rect 41236 10066 41288 10072
rect 41248 8906 41276 10066
rect 41328 9172 41380 9178
rect 41328 9114 41380 9120
rect 41340 8906 41368 9114
rect 41236 8900 41288 8906
rect 41236 8842 41288 8848
rect 41328 8900 41380 8906
rect 41328 8842 41380 8848
rect 41432 5846 41460 11183
rect 41616 11098 41644 13330
rect 41708 13190 41736 13874
rect 41696 13184 41748 13190
rect 41696 13126 41748 13132
rect 41800 12850 41828 14214
rect 41788 12844 41840 12850
rect 41788 12786 41840 12792
rect 41694 11792 41750 11801
rect 41694 11727 41750 11736
rect 41524 11070 41644 11098
rect 41420 5840 41472 5846
rect 41420 5782 41472 5788
rect 41420 5636 41472 5642
rect 41420 5578 41472 5584
rect 41156 5086 41276 5114
rect 41144 5024 41196 5030
rect 41144 4966 41196 4972
rect 41156 3534 41184 4966
rect 41144 3528 41196 3534
rect 41144 3470 41196 3476
rect 41248 3346 41276 5086
rect 41156 3318 41276 3346
rect 41156 3058 41184 3318
rect 41432 3210 41460 5578
rect 41524 4146 41552 11070
rect 41604 5228 41656 5234
rect 41604 5170 41656 5176
rect 41512 4140 41564 4146
rect 41512 4082 41564 4088
rect 41248 3182 41460 3210
rect 41144 3052 41196 3058
rect 41144 2994 41196 3000
rect 41052 2100 41104 2106
rect 41052 2042 41104 2048
rect 41248 800 41276 3182
rect 41512 3052 41564 3058
rect 41512 2994 41564 3000
rect 41524 800 41552 2994
rect 41616 2854 41644 5170
rect 41708 5030 41736 11727
rect 41800 9110 41828 12786
rect 41892 9353 41920 17478
rect 41984 10674 42012 20742
rect 42076 16590 42104 55218
rect 42156 19780 42208 19786
rect 42156 19722 42208 19728
rect 42168 19174 42196 19722
rect 42246 19272 42302 19281
rect 42246 19207 42248 19216
rect 42300 19207 42302 19216
rect 42248 19178 42300 19184
rect 42156 19168 42208 19174
rect 42156 19110 42208 19116
rect 42248 18828 42300 18834
rect 42248 18770 42300 18776
rect 42260 18222 42288 18770
rect 42156 18216 42208 18222
rect 42156 18158 42208 18164
rect 42248 18216 42300 18222
rect 42248 18158 42300 18164
rect 42064 16584 42116 16590
rect 42064 16526 42116 16532
rect 42064 16244 42116 16250
rect 42064 16186 42116 16192
rect 42076 15978 42104 16186
rect 42168 16182 42196 18158
rect 42156 16176 42208 16182
rect 42156 16118 42208 16124
rect 42064 15972 42116 15978
rect 42064 15914 42116 15920
rect 42064 13728 42116 13734
rect 42064 13670 42116 13676
rect 42076 12850 42104 13670
rect 42064 12844 42116 12850
rect 42064 12786 42116 12792
rect 42154 12472 42210 12481
rect 42352 12442 42380 58822
rect 42628 58546 42656 61338
rect 42720 59650 42748 61678
rect 42812 61198 42840 63200
rect 42800 61192 42852 61198
rect 43548 61180 43576 63200
rect 44560 61198 44588 63294
rect 45006 63294 45508 63322
rect 45006 63200 45062 63294
rect 45480 61282 45508 63294
rect 45742 63294 46152 63322
rect 45742 63200 45798 63294
rect 45480 61254 45600 61282
rect 45572 61198 45600 61254
rect 46124 61198 46152 63294
rect 46478 63294 46704 63322
rect 46478 63200 46534 63294
rect 43628 61192 43680 61198
rect 43548 61152 43628 61180
rect 42800 61134 42852 61140
rect 43628 61134 43680 61140
rect 44548 61192 44600 61198
rect 44548 61134 44600 61140
rect 45560 61192 45612 61198
rect 45560 61134 45612 61140
rect 46112 61192 46164 61198
rect 46112 61134 46164 61140
rect 42892 61124 42944 61130
rect 42892 61066 42944 61072
rect 42720 59622 42840 59650
rect 42812 59566 42840 59622
rect 42708 59560 42760 59566
rect 42708 59502 42760 59508
rect 42800 59560 42852 59566
rect 42800 59502 42852 59508
rect 42616 58540 42668 58546
rect 42616 58482 42668 58488
rect 42720 57361 42748 59502
rect 42706 57352 42762 57361
rect 42706 57287 42762 57296
rect 42904 36922 42932 61066
rect 44456 61056 44508 61062
rect 44456 60998 44508 61004
rect 45376 61056 45428 61062
rect 45376 60998 45428 61004
rect 46112 61056 46164 61062
rect 46112 60998 46164 61004
rect 44468 60858 44496 60998
rect 44456 60852 44508 60858
rect 44456 60794 44508 60800
rect 44180 60512 44232 60518
rect 44180 60454 44232 60460
rect 43536 60036 43588 60042
rect 43536 59978 43588 59984
rect 43548 59566 43576 59978
rect 43536 59560 43588 59566
rect 43536 59502 43588 59508
rect 43996 56840 44048 56846
rect 43996 56782 44048 56788
rect 42892 36916 42944 36922
rect 42892 36858 42944 36864
rect 43260 34468 43312 34474
rect 43260 34410 43312 34416
rect 42432 22160 42484 22166
rect 42432 22102 42484 22108
rect 42444 18358 42472 22102
rect 43272 22094 43300 34410
rect 43628 23520 43680 23526
rect 43628 23462 43680 23468
rect 43640 22094 43668 23462
rect 43272 22066 43392 22094
rect 43640 22066 43760 22094
rect 42892 20936 42944 20942
rect 42892 20878 42944 20884
rect 42984 20936 43036 20942
rect 42984 20878 43036 20884
rect 42524 20868 42576 20874
rect 42524 20810 42576 20816
rect 42536 20534 42564 20810
rect 42524 20528 42576 20534
rect 42524 20470 42576 20476
rect 42536 19990 42564 20470
rect 42708 20392 42760 20398
rect 42708 20334 42760 20340
rect 42524 19984 42576 19990
rect 42524 19926 42576 19932
rect 42720 19854 42748 20334
rect 42708 19848 42760 19854
rect 42708 19790 42760 19796
rect 42800 19712 42852 19718
rect 42800 19654 42852 19660
rect 42812 19378 42840 19654
rect 42800 19372 42852 19378
rect 42800 19314 42852 19320
rect 42904 18902 42932 20878
rect 42616 18896 42668 18902
rect 42616 18838 42668 18844
rect 42892 18896 42944 18902
rect 42892 18838 42944 18844
rect 42628 18426 42656 18838
rect 42996 18748 43024 20878
rect 43076 20800 43128 20806
rect 43076 20742 43128 20748
rect 43088 20534 43116 20742
rect 43076 20528 43128 20534
rect 43076 20470 43128 20476
rect 43076 19712 43128 19718
rect 43076 19654 43128 19660
rect 42904 18744 43024 18748
rect 42892 18738 43024 18744
rect 42944 18720 43024 18738
rect 42892 18680 42944 18686
rect 43088 18442 43116 19654
rect 43168 19372 43220 19378
rect 43168 19314 43220 19320
rect 43180 18698 43208 19314
rect 43260 19168 43312 19174
rect 43260 19110 43312 19116
rect 43272 18902 43300 19110
rect 43260 18896 43312 18902
rect 43260 18838 43312 18844
rect 43168 18692 43220 18698
rect 43168 18634 43220 18640
rect 42616 18420 42668 18426
rect 42616 18362 42668 18368
rect 42996 18414 43116 18442
rect 42432 18352 42484 18358
rect 42800 18352 42852 18358
rect 42432 18294 42484 18300
rect 42798 18320 42800 18329
rect 42852 18320 42854 18329
rect 42444 16130 42472 18294
rect 42708 18284 42760 18290
rect 42798 18255 42854 18264
rect 42892 18284 42944 18290
rect 42708 18226 42760 18232
rect 42892 18226 42944 18232
rect 42720 16658 42748 18226
rect 42904 16726 42932 18226
rect 42892 16720 42944 16726
rect 42892 16662 42944 16668
rect 42708 16652 42760 16658
rect 42708 16594 42760 16600
rect 42890 16552 42946 16561
rect 42890 16487 42946 16496
rect 42904 16182 42932 16487
rect 42892 16176 42944 16182
rect 42444 16102 42656 16130
rect 42892 16118 42944 16124
rect 42444 15502 42472 16102
rect 42524 16040 42576 16046
rect 42524 15982 42576 15988
rect 42628 15994 42656 16102
rect 42892 16040 42944 16046
rect 42628 15988 42892 15994
rect 42628 15982 42944 15988
rect 42536 15706 42564 15982
rect 42628 15966 42932 15982
rect 42524 15700 42576 15706
rect 42524 15642 42576 15648
rect 42432 15496 42484 15502
rect 42432 15438 42484 15444
rect 42522 14512 42578 14521
rect 42522 14447 42578 14456
rect 42154 12407 42210 12416
rect 42340 12436 42392 12442
rect 42064 12232 42116 12238
rect 42064 12174 42116 12180
rect 42076 11762 42104 12174
rect 42064 11756 42116 11762
rect 42064 11698 42116 11704
rect 42064 11552 42116 11558
rect 42064 11494 42116 11500
rect 42076 11286 42104 11494
rect 42064 11280 42116 11286
rect 42064 11222 42116 11228
rect 42064 11008 42116 11014
rect 42064 10950 42116 10956
rect 42076 10742 42104 10950
rect 42064 10736 42116 10742
rect 42064 10678 42116 10684
rect 41972 10668 42024 10674
rect 41972 10610 42024 10616
rect 41878 9344 41934 9353
rect 41878 9279 41934 9288
rect 41788 9104 41840 9110
rect 41788 9046 41840 9052
rect 41970 5808 42026 5817
rect 41970 5743 42026 5752
rect 41880 5228 41932 5234
rect 41880 5170 41932 5176
rect 41696 5024 41748 5030
rect 41696 4966 41748 4972
rect 41604 2848 41656 2854
rect 41604 2790 41656 2796
rect 41892 2774 41920 5170
rect 41984 3670 42012 5743
rect 42064 4208 42116 4214
rect 42064 4150 42116 4156
rect 41972 3664 42024 3670
rect 41972 3606 42024 3612
rect 41800 2746 41920 2774
rect 41800 800 41828 2746
rect 42076 800 42104 4150
rect 42168 3058 42196 12407
rect 42340 12378 42392 12384
rect 42248 12164 42300 12170
rect 42248 12106 42300 12112
rect 42260 11218 42288 12106
rect 42430 11384 42486 11393
rect 42430 11319 42486 11328
rect 42248 11212 42300 11218
rect 42248 11154 42300 11160
rect 42444 11150 42472 11319
rect 42432 11144 42484 11150
rect 42432 11086 42484 11092
rect 42432 9580 42484 9586
rect 42432 9522 42484 9528
rect 42444 3738 42472 9522
rect 42536 8430 42564 14447
rect 42800 14068 42852 14074
rect 42800 14010 42852 14016
rect 42812 13938 42840 14010
rect 42800 13932 42852 13938
rect 42800 13874 42852 13880
rect 42616 13320 42668 13326
rect 42616 13262 42668 13268
rect 42628 13190 42656 13262
rect 42616 13184 42668 13190
rect 42616 13126 42668 13132
rect 42800 12980 42852 12986
rect 42800 12922 42852 12928
rect 42708 11688 42760 11694
rect 42708 11630 42760 11636
rect 42720 11558 42748 11630
rect 42708 11552 42760 11558
rect 42708 11494 42760 11500
rect 42616 11144 42668 11150
rect 42616 11086 42668 11092
rect 42524 8424 42576 8430
rect 42524 8366 42576 8372
rect 42536 7886 42564 8366
rect 42524 7880 42576 7886
rect 42524 7822 42576 7828
rect 42524 4548 42576 4554
rect 42524 4490 42576 4496
rect 42536 3942 42564 4490
rect 42628 4162 42656 11086
rect 42812 5370 42840 12922
rect 42892 11824 42944 11830
rect 42892 11766 42944 11772
rect 42904 11150 42932 11766
rect 42892 11144 42944 11150
rect 42892 11086 42944 11092
rect 42892 10736 42944 10742
rect 42892 10678 42944 10684
rect 42904 10169 42932 10678
rect 42890 10160 42946 10169
rect 42890 10095 42946 10104
rect 42904 5386 42932 10095
rect 42996 8498 43024 18414
rect 43364 18290 43392 22066
rect 43444 20868 43496 20874
rect 43444 20810 43496 20816
rect 43456 20262 43484 20810
rect 43536 20528 43588 20534
rect 43536 20470 43588 20476
rect 43444 20256 43496 20262
rect 43444 20198 43496 20204
rect 43076 18284 43128 18290
rect 43076 18226 43128 18232
rect 43352 18284 43404 18290
rect 43352 18226 43404 18232
rect 43088 17610 43116 18226
rect 43168 18216 43220 18222
rect 43168 18158 43220 18164
rect 43180 17954 43208 18158
rect 43180 17926 43300 17954
rect 43076 17604 43128 17610
rect 43076 17546 43128 17552
rect 43168 16516 43220 16522
rect 43168 16458 43220 16464
rect 43180 16250 43208 16458
rect 43168 16244 43220 16250
rect 43168 16186 43220 16192
rect 43272 16046 43300 17926
rect 43260 16040 43312 16046
rect 43260 15982 43312 15988
rect 43548 15026 43576 20470
rect 43732 19718 43760 22066
rect 43904 20596 43956 20602
rect 43904 20538 43956 20544
rect 43812 20256 43864 20262
rect 43812 20198 43864 20204
rect 43720 19712 43772 19718
rect 43720 19654 43772 19660
rect 43732 19446 43760 19654
rect 43720 19440 43772 19446
rect 43720 19382 43772 19388
rect 43824 19292 43852 20198
rect 43916 19446 43944 20538
rect 43904 19440 43956 19446
rect 43904 19382 43956 19388
rect 43824 19264 43944 19292
rect 43916 19174 43944 19264
rect 43904 19168 43956 19174
rect 43626 19136 43682 19145
rect 43904 19110 43956 19116
rect 43626 19071 43682 19080
rect 43640 18766 43668 19071
rect 43628 18760 43680 18766
rect 43628 18702 43680 18708
rect 43720 18692 43772 18698
rect 43720 18634 43772 18640
rect 43536 15020 43588 15026
rect 43536 14962 43588 14968
rect 43168 14952 43220 14958
rect 43168 14894 43220 14900
rect 43076 14408 43128 14414
rect 43076 14350 43128 14356
rect 43088 13938 43116 14350
rect 43076 13932 43128 13938
rect 43076 13874 43128 13880
rect 43180 13326 43208 14894
rect 43260 14408 43312 14414
rect 43260 14350 43312 14356
rect 43272 13530 43300 14350
rect 43352 13864 43404 13870
rect 43548 13818 43576 14962
rect 43352 13806 43404 13812
rect 43260 13524 43312 13530
rect 43260 13466 43312 13472
rect 43168 13320 43220 13326
rect 43168 13262 43220 13268
rect 43180 12782 43208 13262
rect 43364 12986 43392 13806
rect 43456 13790 43576 13818
rect 43352 12980 43404 12986
rect 43352 12922 43404 12928
rect 43168 12776 43220 12782
rect 43168 12718 43220 12724
rect 43456 12714 43484 13790
rect 43536 13728 43588 13734
rect 43588 13676 43668 13682
rect 43536 13670 43668 13676
rect 43548 13654 43668 13670
rect 43536 12912 43588 12918
rect 43536 12854 43588 12860
rect 43444 12708 43496 12714
rect 43444 12650 43496 12656
rect 43352 12164 43404 12170
rect 43352 12106 43404 12112
rect 43260 12096 43312 12102
rect 43260 12038 43312 12044
rect 43272 11762 43300 12038
rect 43076 11756 43128 11762
rect 43076 11698 43128 11704
rect 43260 11756 43312 11762
rect 43260 11698 43312 11704
rect 43088 11286 43116 11698
rect 43168 11552 43220 11558
rect 43168 11494 43220 11500
rect 43076 11280 43128 11286
rect 43076 11222 43128 11228
rect 43180 10962 43208 11494
rect 43088 10934 43208 10962
rect 42984 8492 43036 8498
rect 42984 8434 43036 8440
rect 42800 5364 42852 5370
rect 42904 5358 43024 5386
rect 42800 5306 42852 5312
rect 42892 5228 42944 5234
rect 42892 5170 42944 5176
rect 42628 4134 42748 4162
rect 42614 4040 42670 4049
rect 42614 3975 42670 3984
rect 42524 3936 42576 3942
rect 42524 3878 42576 3884
rect 42432 3732 42484 3738
rect 42432 3674 42484 3680
rect 42536 3534 42564 3878
rect 42524 3528 42576 3534
rect 42524 3470 42576 3476
rect 42628 3058 42656 3975
rect 42720 3913 42748 4134
rect 42706 3904 42762 3913
rect 42706 3839 42762 3848
rect 42708 3664 42760 3670
rect 42708 3606 42760 3612
rect 42156 3052 42208 3058
rect 42156 2994 42208 3000
rect 42616 3052 42668 3058
rect 42616 2994 42668 3000
rect 42340 2848 42392 2854
rect 42340 2790 42392 2796
rect 42248 2304 42300 2310
rect 42248 2246 42300 2252
rect 42260 2038 42288 2246
rect 42248 2032 42300 2038
rect 42248 1974 42300 1980
rect 42352 800 42380 2790
rect 42614 2680 42670 2689
rect 42614 2615 42670 2624
rect 42628 2446 42656 2615
rect 42616 2440 42668 2446
rect 42616 2382 42668 2388
rect 42720 1748 42748 3606
rect 42800 2644 42852 2650
rect 42800 2586 42852 2592
rect 42812 2446 42840 2586
rect 42800 2440 42852 2446
rect 42800 2382 42852 2388
rect 42628 1720 42748 1748
rect 42628 800 42656 1720
rect 42904 800 42932 5170
rect 42996 4690 43024 5358
rect 42984 4684 43036 4690
rect 42984 4626 43036 4632
rect 42984 3052 43036 3058
rect 42984 2994 43036 3000
rect 42996 2514 43024 2994
rect 42984 2508 43036 2514
rect 42984 2450 43036 2456
rect 43088 1766 43116 10934
rect 43168 8288 43220 8294
rect 43168 8230 43220 8236
rect 43180 8022 43208 8230
rect 43168 8016 43220 8022
rect 43168 7958 43220 7964
rect 43168 7336 43220 7342
rect 43168 7278 43220 7284
rect 43180 5370 43208 7278
rect 43168 5364 43220 5370
rect 43168 5306 43220 5312
rect 43364 4758 43392 12106
rect 43444 8900 43496 8906
rect 43444 8842 43496 8848
rect 43456 8294 43484 8842
rect 43444 8288 43496 8294
rect 43444 8230 43496 8236
rect 43456 7886 43484 8230
rect 43444 7880 43496 7886
rect 43444 7822 43496 7828
rect 43352 4752 43404 4758
rect 43352 4694 43404 4700
rect 43364 4593 43392 4694
rect 43350 4584 43406 4593
rect 43350 4519 43406 4528
rect 43364 4146 43392 4519
rect 43352 4140 43404 4146
rect 43180 4100 43352 4128
rect 43180 3058 43208 4100
rect 43352 4082 43404 4088
rect 43444 4072 43496 4078
rect 43350 4040 43406 4049
rect 43444 4014 43496 4020
rect 43350 3975 43406 3984
rect 43364 3602 43392 3975
rect 43456 3777 43484 4014
rect 43548 4010 43576 12854
rect 43640 4826 43668 13654
rect 43732 13190 43760 18634
rect 43916 17134 43944 19110
rect 43904 17128 43956 17134
rect 43904 17070 43956 17076
rect 43720 13184 43772 13190
rect 43720 13126 43772 13132
rect 43720 12164 43772 12170
rect 43720 12106 43772 12112
rect 43732 11694 43760 12106
rect 43720 11688 43772 11694
rect 43720 11630 43772 11636
rect 43720 8900 43772 8906
rect 43720 8842 43772 8848
rect 43732 8090 43760 8842
rect 43916 8430 43944 17070
rect 44008 11830 44036 56782
rect 44192 55350 44220 60454
rect 44180 55344 44232 55350
rect 44180 55286 44232 55292
rect 45388 53174 45416 60998
rect 46124 53514 46152 60998
rect 46676 60790 46704 63294
rect 47214 63200 47270 64000
rect 47950 63322 48006 64000
rect 47950 63294 48268 63322
rect 47950 63200 48006 63294
rect 46848 61668 46900 61674
rect 46848 61610 46900 61616
rect 46860 61402 46888 61610
rect 46848 61396 46900 61402
rect 46848 61338 46900 61344
rect 47228 61198 47256 63200
rect 47216 61192 47268 61198
rect 48240 61180 48268 63294
rect 48686 63200 48742 64000
rect 49422 63322 49478 64000
rect 49422 63294 49648 63322
rect 49422 63200 49478 63294
rect 48700 61198 48728 63200
rect 49424 61804 49476 61810
rect 49424 61746 49476 61752
rect 49436 61402 49464 61746
rect 49424 61396 49476 61402
rect 49424 61338 49476 61344
rect 48320 61192 48372 61198
rect 48240 61152 48320 61180
rect 47216 61134 47268 61140
rect 48320 61134 48372 61140
rect 48688 61192 48740 61198
rect 49620 61180 49648 63294
rect 50158 63200 50214 64000
rect 50894 63322 50950 64000
rect 50894 63294 51028 63322
rect 50894 63200 50950 63294
rect 49700 61192 49752 61198
rect 49620 61152 49700 61180
rect 48688 61134 48740 61140
rect 49700 61134 49752 61140
rect 46848 61056 46900 61062
rect 46848 60998 46900 61004
rect 50068 61056 50120 61062
rect 50068 60998 50120 61004
rect 46664 60784 46716 60790
rect 46664 60726 46716 60732
rect 46860 56370 46888 60998
rect 49608 56772 49660 56778
rect 49608 56714 49660 56720
rect 46848 56364 46900 56370
rect 46848 56306 46900 56312
rect 49620 56166 49648 56714
rect 49608 56160 49660 56166
rect 49608 56102 49660 56108
rect 50080 55214 50108 60998
rect 50172 60790 50200 63200
rect 51000 61180 51028 63294
rect 51630 63200 51686 64000
rect 52366 63200 52422 64000
rect 53102 63322 53158 64000
rect 53838 63322 53894 64000
rect 54574 63322 54630 64000
rect 55310 63322 55366 64000
rect 53102 63294 53236 63322
rect 53102 63200 53158 63294
rect 51448 61600 51500 61606
rect 51448 61542 51500 61548
rect 51460 61402 51488 61542
rect 51448 61396 51500 61402
rect 51448 61338 51500 61344
rect 51644 61198 51672 63200
rect 51080 61192 51132 61198
rect 51000 61152 51080 61180
rect 51080 61134 51132 61140
rect 51632 61192 51684 61198
rect 51632 61134 51684 61140
rect 50294 60956 50602 60965
rect 50294 60954 50300 60956
rect 50356 60954 50380 60956
rect 50436 60954 50460 60956
rect 50516 60954 50540 60956
rect 50596 60954 50602 60956
rect 50356 60902 50358 60954
rect 50538 60902 50540 60954
rect 50294 60900 50300 60902
rect 50356 60900 50380 60902
rect 50436 60900 50460 60902
rect 50516 60900 50540 60902
rect 50596 60900 50602 60902
rect 50294 60891 50602 60900
rect 52380 60874 52408 63200
rect 53208 61198 53236 63294
rect 53838 63294 54156 63322
rect 53838 63200 53894 63294
rect 53380 61260 53432 61266
rect 53380 61202 53432 61208
rect 53196 61192 53248 61198
rect 53392 61169 53420 61202
rect 54128 61198 54156 63294
rect 54574 63294 54708 63322
rect 54574 63200 54630 63294
rect 54116 61192 54168 61198
rect 53196 61134 53248 61140
rect 53378 61160 53434 61169
rect 54116 61134 54168 61140
rect 53378 61095 53434 61104
rect 53196 61056 53248 61062
rect 53196 60998 53248 61004
rect 54300 61056 54352 61062
rect 54300 60998 54352 61004
rect 52380 60846 52500 60874
rect 52472 60790 52500 60846
rect 50160 60784 50212 60790
rect 50160 60726 50212 60732
rect 52460 60784 52512 60790
rect 52460 60726 52512 60732
rect 50436 60512 50488 60518
rect 50436 60454 50488 60460
rect 53104 60512 53156 60518
rect 53104 60454 53156 60460
rect 50448 60246 50476 60454
rect 50436 60240 50488 60246
rect 50436 60182 50488 60188
rect 50294 59868 50602 59877
rect 50294 59866 50300 59868
rect 50356 59866 50380 59868
rect 50436 59866 50460 59868
rect 50516 59866 50540 59868
rect 50596 59866 50602 59868
rect 50356 59814 50358 59866
rect 50538 59814 50540 59866
rect 50294 59812 50300 59814
rect 50356 59812 50380 59814
rect 50436 59812 50460 59814
rect 50516 59812 50540 59814
rect 50596 59812 50602 59814
rect 50294 59803 50602 59812
rect 53116 59634 53144 60454
rect 53104 59628 53156 59634
rect 53104 59570 53156 59576
rect 50294 58780 50602 58789
rect 50294 58778 50300 58780
rect 50356 58778 50380 58780
rect 50436 58778 50460 58780
rect 50516 58778 50540 58780
rect 50596 58778 50602 58780
rect 50356 58726 50358 58778
rect 50538 58726 50540 58778
rect 50294 58724 50300 58726
rect 50356 58724 50380 58726
rect 50436 58724 50460 58726
rect 50516 58724 50540 58726
rect 50596 58724 50602 58726
rect 50294 58715 50602 58724
rect 52460 58336 52512 58342
rect 52460 58278 52512 58284
rect 52472 57934 52500 58278
rect 52460 57928 52512 57934
rect 52460 57870 52512 57876
rect 50294 57692 50602 57701
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57627 50602 57636
rect 51724 56772 51776 56778
rect 51724 56714 51776 56720
rect 50294 56604 50602 56613
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56539 50602 56548
rect 50294 55516 50602 55525
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55451 50602 55460
rect 50080 55186 50200 55214
rect 46112 53508 46164 53514
rect 46112 53450 46164 53456
rect 45376 53168 45428 53174
rect 45376 53110 45428 53116
rect 45744 44396 45796 44402
rect 45744 44338 45796 44344
rect 45100 40452 45152 40458
rect 45100 40394 45152 40400
rect 44180 37800 44232 37806
rect 44180 37742 44232 37748
rect 44192 31142 44220 37742
rect 44180 31136 44232 31142
rect 44180 31078 44232 31084
rect 44824 29504 44876 29510
rect 44824 29446 44876 29452
rect 44456 25288 44508 25294
rect 44456 25230 44508 25236
rect 44088 23112 44140 23118
rect 44088 23054 44140 23060
rect 44100 20602 44128 23054
rect 44364 20936 44416 20942
rect 44364 20878 44416 20884
rect 44088 20596 44140 20602
rect 44088 20538 44140 20544
rect 44100 18834 44128 20538
rect 44376 20466 44404 20878
rect 44364 20460 44416 20466
rect 44364 20402 44416 20408
rect 44468 19990 44496 25230
rect 44836 22982 44864 29446
rect 44824 22976 44876 22982
rect 44824 22918 44876 22924
rect 44456 19984 44508 19990
rect 44456 19926 44508 19932
rect 44468 19310 44496 19926
rect 44456 19304 44508 19310
rect 44456 19246 44508 19252
rect 44088 18828 44140 18834
rect 44088 18770 44140 18776
rect 44180 18284 44232 18290
rect 44180 18226 44232 18232
rect 44192 16998 44220 18226
rect 44180 16992 44232 16998
rect 44180 16934 44232 16940
rect 44732 16652 44784 16658
rect 44732 16594 44784 16600
rect 44180 16108 44232 16114
rect 44180 16050 44232 16056
rect 44192 15502 44220 16050
rect 44180 15496 44232 15502
rect 44180 15438 44232 15444
rect 44088 14068 44140 14074
rect 44088 14010 44140 14016
rect 43996 11824 44048 11830
rect 43996 11766 44048 11772
rect 44100 10062 44128 14010
rect 44192 11898 44220 15438
rect 44364 14952 44416 14958
rect 44364 14894 44416 14900
rect 44376 14618 44404 14894
rect 44364 14612 44416 14618
rect 44364 14554 44416 14560
rect 44548 14612 44600 14618
rect 44548 14554 44600 14560
rect 44560 13258 44588 14554
rect 44548 13252 44600 13258
rect 44548 13194 44600 13200
rect 44456 13184 44508 13190
rect 44456 13126 44508 13132
rect 44180 11892 44232 11898
rect 44180 11834 44232 11840
rect 44192 10674 44220 11834
rect 44272 11824 44324 11830
rect 44272 11766 44324 11772
rect 44180 10668 44232 10674
rect 44180 10610 44232 10616
rect 44088 10056 44140 10062
rect 44088 9998 44140 10004
rect 43996 9512 44048 9518
rect 43996 9454 44048 9460
rect 43904 8424 43956 8430
rect 43904 8366 43956 8372
rect 43720 8084 43772 8090
rect 43720 8026 43772 8032
rect 44008 7886 44036 9454
rect 44100 9042 44128 9998
rect 44284 9654 44312 11766
rect 44468 11150 44496 13126
rect 44640 12368 44692 12374
rect 44640 12310 44692 12316
rect 44456 11144 44508 11150
rect 44456 11086 44508 11092
rect 44546 10296 44602 10305
rect 44546 10231 44602 10240
rect 44560 10198 44588 10231
rect 44548 10192 44600 10198
rect 44548 10134 44600 10140
rect 44272 9648 44324 9654
rect 44272 9590 44324 9596
rect 44180 9580 44232 9586
rect 44180 9522 44232 9528
rect 44088 9036 44140 9042
rect 44088 8978 44140 8984
rect 44100 8906 44128 8978
rect 44088 8900 44140 8906
rect 44088 8842 44140 8848
rect 44192 7886 44220 9522
rect 44284 8498 44312 9590
rect 44456 9444 44508 9450
rect 44456 9386 44508 9392
rect 44468 9042 44496 9386
rect 44456 9036 44508 9042
rect 44456 8978 44508 8984
rect 44272 8492 44324 8498
rect 44272 8434 44324 8440
rect 44548 8492 44600 8498
rect 44548 8434 44600 8440
rect 43996 7880 44048 7886
rect 43996 7822 44048 7828
rect 44180 7880 44232 7886
rect 44180 7822 44232 7828
rect 43904 7812 43956 7818
rect 43904 7754 43956 7760
rect 44456 7812 44508 7818
rect 44456 7754 44508 7760
rect 43916 7410 43944 7754
rect 44468 7546 44496 7754
rect 44456 7540 44508 7546
rect 44456 7482 44508 7488
rect 44560 7410 44588 8434
rect 43904 7404 43956 7410
rect 43904 7346 43956 7352
rect 44548 7404 44600 7410
rect 44548 7346 44600 7352
rect 44560 6798 44588 7346
rect 44548 6792 44600 6798
rect 44548 6734 44600 6740
rect 44180 5228 44232 5234
rect 44180 5170 44232 5176
rect 44548 5228 44600 5234
rect 44548 5170 44600 5176
rect 43628 4820 43680 4826
rect 43628 4762 43680 4768
rect 43640 4690 43944 4706
rect 43640 4684 43956 4690
rect 43640 4678 43904 4684
rect 43640 4622 43668 4678
rect 43904 4626 43956 4632
rect 43628 4616 43680 4622
rect 43996 4616 44048 4622
rect 43628 4558 43680 4564
rect 43994 4584 43996 4593
rect 44048 4584 44050 4593
rect 44050 4542 44128 4570
rect 43994 4519 44050 4528
rect 43536 4004 43588 4010
rect 43536 3946 43588 3952
rect 43628 3936 43680 3942
rect 43628 3878 43680 3884
rect 43996 3936 44048 3942
rect 43996 3878 44048 3884
rect 43442 3768 43498 3777
rect 43442 3703 43498 3712
rect 43352 3596 43404 3602
rect 43352 3538 43404 3544
rect 43640 3482 43668 3878
rect 43720 3732 43772 3738
rect 43720 3674 43772 3680
rect 43548 3454 43668 3482
rect 43260 3392 43312 3398
rect 43260 3334 43312 3340
rect 43168 3052 43220 3058
rect 43168 2994 43220 3000
rect 43272 2774 43300 3334
rect 43548 2990 43576 3454
rect 43628 3392 43680 3398
rect 43628 3334 43680 3340
rect 43640 3058 43668 3334
rect 43628 3052 43680 3058
rect 43628 2994 43680 3000
rect 43352 2984 43404 2990
rect 43352 2926 43404 2932
rect 43536 2984 43588 2990
rect 43536 2926 43588 2932
rect 43180 2746 43300 2774
rect 43076 1760 43128 1766
rect 43076 1702 43128 1708
rect 43180 800 43208 2746
rect 43364 2689 43392 2926
rect 43444 2916 43496 2922
rect 43444 2858 43496 2864
rect 43350 2680 43406 2689
rect 43350 2615 43406 2624
rect 43352 2304 43404 2310
rect 43352 2246 43404 2252
rect 43364 2106 43392 2246
rect 43352 2100 43404 2106
rect 43352 2042 43404 2048
rect 43456 800 43484 2858
rect 43548 2446 43576 2926
rect 43626 2680 43682 2689
rect 43626 2615 43682 2624
rect 43536 2440 43588 2446
rect 43536 2382 43588 2388
rect 43640 2106 43668 2615
rect 43628 2100 43680 2106
rect 43628 2042 43680 2048
rect 43732 800 43760 3674
rect 43810 3632 43866 3641
rect 43810 3567 43812 3576
rect 43864 3567 43866 3576
rect 43812 3538 43864 3544
rect 43904 2372 43956 2378
rect 43904 2314 43956 2320
rect 43916 1698 43944 2314
rect 43904 1692 43956 1698
rect 43904 1634 43956 1640
rect 44008 800 44036 3878
rect 44100 3602 44128 4542
rect 44192 3738 44220 5170
rect 44456 5092 44508 5098
rect 44456 5034 44508 5040
rect 44272 5024 44324 5030
rect 44272 4966 44324 4972
rect 44284 4826 44312 4966
rect 44272 4820 44324 4826
rect 44272 4762 44324 4768
rect 44364 4480 44416 4486
rect 44364 4422 44416 4428
rect 44376 4146 44404 4422
rect 44364 4140 44416 4146
rect 44364 4082 44416 4088
rect 44364 4004 44416 4010
rect 44364 3946 44416 3952
rect 44376 3738 44404 3946
rect 44180 3732 44232 3738
rect 44180 3674 44232 3680
rect 44364 3732 44416 3738
rect 44364 3674 44416 3680
rect 44178 3632 44234 3641
rect 44088 3596 44140 3602
rect 44178 3567 44234 3576
rect 44088 3538 44140 3544
rect 44192 3534 44220 3567
rect 44180 3528 44232 3534
rect 44180 3470 44232 3476
rect 44364 3052 44416 3058
rect 44364 2994 44416 3000
rect 44180 2848 44232 2854
rect 44180 2790 44232 2796
rect 44192 2310 44220 2790
rect 44180 2304 44232 2310
rect 44180 2246 44232 2252
rect 44376 1442 44404 2994
rect 44468 2446 44496 5034
rect 44456 2440 44508 2446
rect 44456 2382 44508 2388
rect 44284 1414 44404 1442
rect 44284 800 44312 1414
rect 44560 800 44588 5170
rect 44652 5098 44680 12310
rect 44640 5092 44692 5098
rect 44640 5034 44692 5040
rect 44744 4078 44772 16594
rect 45112 12434 45140 40394
rect 45284 20324 45336 20330
rect 45284 20266 45336 20272
rect 45296 19786 45324 20266
rect 45376 19848 45428 19854
rect 45376 19790 45428 19796
rect 45284 19780 45336 19786
rect 45284 19722 45336 19728
rect 45388 19378 45416 19790
rect 45560 19780 45612 19786
rect 45560 19722 45612 19728
rect 45376 19372 45428 19378
rect 45376 19314 45428 19320
rect 45284 18896 45336 18902
rect 45284 18838 45336 18844
rect 45296 18630 45324 18838
rect 45284 18624 45336 18630
rect 45284 18566 45336 18572
rect 45296 18358 45324 18566
rect 45284 18352 45336 18358
rect 45284 18294 45336 18300
rect 45192 16652 45244 16658
rect 45192 16594 45244 16600
rect 44928 12406 45140 12434
rect 44824 10464 44876 10470
rect 44824 10406 44876 10412
rect 44836 10130 44864 10406
rect 44824 10124 44876 10130
rect 44824 10066 44876 10072
rect 44824 8492 44876 8498
rect 44824 8434 44876 8440
rect 44836 8294 44864 8434
rect 44824 8288 44876 8294
rect 44824 8230 44876 8236
rect 44732 4072 44784 4078
rect 44732 4014 44784 4020
rect 44824 4004 44876 4010
rect 44824 3946 44876 3952
rect 44836 800 44864 3946
rect 44928 3194 44956 12406
rect 45204 11762 45232 16594
rect 45388 16250 45416 19314
rect 45572 18698 45600 19722
rect 45652 19372 45704 19378
rect 45652 19314 45704 19320
rect 45664 18970 45692 19314
rect 45652 18964 45704 18970
rect 45652 18906 45704 18912
rect 45560 18692 45612 18698
rect 45560 18634 45612 18640
rect 45376 16244 45428 16250
rect 45376 16186 45428 16192
rect 45192 11756 45244 11762
rect 45192 11698 45244 11704
rect 45468 11756 45520 11762
rect 45468 11698 45520 11704
rect 45560 11756 45612 11762
rect 45560 11698 45612 11704
rect 45100 11144 45152 11150
rect 45100 11086 45152 11092
rect 45008 9036 45060 9042
rect 45008 8978 45060 8984
rect 45020 6361 45048 8978
rect 45112 8974 45140 11086
rect 45192 10464 45244 10470
rect 45192 10406 45244 10412
rect 45204 9586 45232 10406
rect 45480 10266 45508 11698
rect 45468 10260 45520 10266
rect 45468 10202 45520 10208
rect 45468 9920 45520 9926
rect 45468 9862 45520 9868
rect 45480 9654 45508 9862
rect 45468 9648 45520 9654
rect 45468 9590 45520 9596
rect 45192 9580 45244 9586
rect 45192 9522 45244 9528
rect 45100 8968 45152 8974
rect 45100 8910 45152 8916
rect 45204 8566 45232 9522
rect 45192 8560 45244 8566
rect 45192 8502 45244 8508
rect 45204 7426 45232 8502
rect 45376 8424 45428 8430
rect 45376 8366 45428 8372
rect 45468 8424 45520 8430
rect 45468 8366 45520 8372
rect 45388 7886 45416 8366
rect 45480 8294 45508 8366
rect 45468 8288 45520 8294
rect 45468 8230 45520 8236
rect 45284 7880 45336 7886
rect 45284 7822 45336 7828
rect 45376 7880 45428 7886
rect 45376 7822 45428 7828
rect 45112 7410 45232 7426
rect 45100 7404 45232 7410
rect 45152 7398 45232 7404
rect 45100 7346 45152 7352
rect 45296 7002 45324 7822
rect 45284 6996 45336 7002
rect 45284 6938 45336 6944
rect 45480 6798 45508 8230
rect 45468 6792 45520 6798
rect 45468 6734 45520 6740
rect 45006 6352 45062 6361
rect 45006 6287 45062 6296
rect 45192 5092 45244 5098
rect 45192 5034 45244 5040
rect 45008 5024 45060 5030
rect 45008 4966 45060 4972
rect 45020 4185 45048 4966
rect 45100 4548 45152 4554
rect 45100 4490 45152 4496
rect 45006 4176 45062 4185
rect 45006 4111 45062 4120
rect 45112 3754 45140 4490
rect 45204 4162 45232 5034
rect 45376 4208 45428 4214
rect 45204 4134 45324 4162
rect 45376 4150 45428 4156
rect 45190 4040 45246 4049
rect 45190 3975 45246 3984
rect 45020 3726 45140 3754
rect 44916 3188 44968 3194
rect 44916 3130 44968 3136
rect 45020 3058 45048 3726
rect 45100 3664 45152 3670
rect 45100 3606 45152 3612
rect 45008 3052 45060 3058
rect 45008 2994 45060 3000
rect 45008 2644 45060 2650
rect 45008 2586 45060 2592
rect 45020 2514 45048 2586
rect 45008 2508 45060 2514
rect 45008 2450 45060 2456
rect 45112 800 45140 3606
rect 45204 3194 45232 3975
rect 45192 3188 45244 3194
rect 45192 3130 45244 3136
rect 45296 2990 45324 4134
rect 45284 2984 45336 2990
rect 45284 2926 45336 2932
rect 45388 2922 45416 4150
rect 45468 4072 45520 4078
rect 45468 4014 45520 4020
rect 45480 3913 45508 4014
rect 45466 3904 45522 3913
rect 45466 3839 45522 3848
rect 45468 3392 45520 3398
rect 45468 3334 45520 3340
rect 45376 2916 45428 2922
rect 45376 2858 45428 2864
rect 45374 2680 45430 2689
rect 45374 2615 45376 2624
rect 45428 2615 45430 2624
rect 45376 2586 45428 2592
rect 45192 2440 45244 2446
rect 45192 2382 45244 2388
rect 45204 1086 45232 2382
rect 45480 1442 45508 3334
rect 45572 3126 45600 11698
rect 45652 10464 45704 10470
rect 45652 10406 45704 10412
rect 45664 10130 45692 10406
rect 45652 10124 45704 10130
rect 45652 10066 45704 10072
rect 45652 5228 45704 5234
rect 45652 5170 45704 5176
rect 45560 3120 45612 3126
rect 45560 3062 45612 3068
rect 45388 1414 45508 1442
rect 45192 1080 45244 1086
rect 45192 1022 45244 1028
rect 45388 800 45416 1414
rect 45664 800 45692 5170
rect 45756 2774 45784 44338
rect 47584 40384 47636 40390
rect 47584 40326 47636 40332
rect 46848 38344 46900 38350
rect 46848 38286 46900 38292
rect 46296 34060 46348 34066
rect 46296 34002 46348 34008
rect 46308 23594 46336 34002
rect 46480 28552 46532 28558
rect 46480 28494 46532 28500
rect 46296 23588 46348 23594
rect 46296 23530 46348 23536
rect 46296 19712 46348 19718
rect 46296 19654 46348 19660
rect 46308 18766 46336 19654
rect 46386 19272 46442 19281
rect 46386 19207 46388 19216
rect 46440 19207 46442 19216
rect 46388 19178 46440 19184
rect 45928 18760 45980 18766
rect 45928 18702 45980 18708
rect 46020 18760 46072 18766
rect 46020 18702 46072 18708
rect 46296 18760 46348 18766
rect 46296 18702 46348 18708
rect 46388 18760 46440 18766
rect 46388 18702 46440 18708
rect 45836 18624 45888 18630
rect 45836 18566 45888 18572
rect 45848 18426 45876 18566
rect 45940 18426 45968 18702
rect 45836 18420 45888 18426
rect 45836 18362 45888 18368
rect 45928 18420 45980 18426
rect 45928 18362 45980 18368
rect 46032 17882 46060 18702
rect 46400 18290 46428 18702
rect 46388 18284 46440 18290
rect 46388 18226 46440 18232
rect 46020 17876 46072 17882
rect 46020 17818 46072 17824
rect 46388 16516 46440 16522
rect 46388 16458 46440 16464
rect 46400 16250 46428 16458
rect 46388 16244 46440 16250
rect 46388 16186 46440 16192
rect 46296 11892 46348 11898
rect 46296 11834 46348 11840
rect 46112 11756 46164 11762
rect 46112 11698 46164 11704
rect 46124 11354 46152 11698
rect 46112 11348 46164 11354
rect 46112 11290 46164 11296
rect 46308 11150 46336 11834
rect 46296 11144 46348 11150
rect 46296 11086 46348 11092
rect 46112 10056 46164 10062
rect 46112 9998 46164 10004
rect 46018 9208 46074 9217
rect 46018 9143 46074 9152
rect 45836 7404 45888 7410
rect 45836 7346 45888 7352
rect 45848 7002 45876 7346
rect 45928 7200 45980 7206
rect 45928 7142 45980 7148
rect 45940 7002 45968 7142
rect 45836 6996 45888 7002
rect 45836 6938 45888 6944
rect 45928 6996 45980 7002
rect 45928 6938 45980 6944
rect 46032 6780 46060 9143
rect 46124 8974 46152 9998
rect 46296 9920 46348 9926
rect 46296 9862 46348 9868
rect 46308 9586 46336 9862
rect 46296 9580 46348 9586
rect 46296 9522 46348 9528
rect 46204 9036 46256 9042
rect 46204 8978 46256 8984
rect 46112 8968 46164 8974
rect 46112 8910 46164 8916
rect 46124 8634 46152 8910
rect 46216 8634 46244 8978
rect 46308 8974 46336 9522
rect 46296 8968 46348 8974
rect 46296 8910 46348 8916
rect 46112 8628 46164 8634
rect 46112 8570 46164 8576
rect 46204 8628 46256 8634
rect 46204 8570 46256 8576
rect 46388 8492 46440 8498
rect 46388 8434 46440 8440
rect 46400 8090 46428 8434
rect 46388 8084 46440 8090
rect 46388 8026 46440 8032
rect 46388 7200 46440 7206
rect 46388 7142 46440 7148
rect 46400 6866 46428 7142
rect 46388 6860 46440 6866
rect 46388 6802 46440 6808
rect 46032 6752 46152 6780
rect 46020 4548 46072 4554
rect 46020 4490 46072 4496
rect 45928 4140 45980 4146
rect 45928 4082 45980 4088
rect 45940 3942 45968 4082
rect 45928 3936 45980 3942
rect 45928 3878 45980 3884
rect 46032 3670 46060 4490
rect 46124 4214 46152 6752
rect 46112 4208 46164 4214
rect 46112 4150 46164 4156
rect 46020 3664 46072 3670
rect 46020 3606 46072 3612
rect 46492 3194 46520 28494
rect 46860 26234 46888 38286
rect 47308 28416 47360 28422
rect 47308 28358 47360 28364
rect 46676 26206 46888 26234
rect 46676 19174 46704 26206
rect 47032 20460 47084 20466
rect 47032 20402 47084 20408
rect 46848 20392 46900 20398
rect 46848 20334 46900 20340
rect 46860 19786 46888 20334
rect 46848 19780 46900 19786
rect 46848 19722 46900 19728
rect 46664 19168 46716 19174
rect 46664 19110 46716 19116
rect 46940 19168 46992 19174
rect 46940 19110 46992 19116
rect 46570 18592 46626 18601
rect 46570 18527 46626 18536
rect 46584 18426 46612 18527
rect 46572 18420 46624 18426
rect 46572 18362 46624 18368
rect 46676 18358 46704 19110
rect 46952 18850 46980 19110
rect 47044 18970 47072 20402
rect 47216 20256 47268 20262
rect 47216 20198 47268 20204
rect 47228 19854 47256 20198
rect 47216 19848 47268 19854
rect 47216 19790 47268 19796
rect 47032 18964 47084 18970
rect 47032 18906 47084 18912
rect 46768 18822 46980 18850
rect 46768 18698 46796 18822
rect 46756 18692 46808 18698
rect 46756 18634 46808 18640
rect 46848 18692 46900 18698
rect 46848 18634 46900 18640
rect 46664 18352 46716 18358
rect 46664 18294 46716 18300
rect 46572 16448 46624 16454
rect 46572 16390 46624 16396
rect 46584 16250 46612 16390
rect 46572 16244 46624 16250
rect 46572 16186 46624 16192
rect 46584 16153 46612 16186
rect 46570 16144 46626 16153
rect 46570 16079 46626 16088
rect 46756 16108 46808 16114
rect 46756 16050 46808 16056
rect 46572 16040 46624 16046
rect 46572 15982 46624 15988
rect 46584 11286 46612 15982
rect 46768 15638 46796 16050
rect 46756 15632 46808 15638
rect 46756 15574 46808 15580
rect 46664 12980 46716 12986
rect 46664 12922 46716 12928
rect 46572 11280 46624 11286
rect 46572 11222 46624 11228
rect 46584 10606 46612 11222
rect 46572 10600 46624 10606
rect 46572 10542 46624 10548
rect 46584 9602 46612 10542
rect 46676 10130 46704 12922
rect 46860 11642 46888 18634
rect 46940 18352 46992 18358
rect 46938 18320 46940 18329
rect 46992 18320 46994 18329
rect 46938 18255 46994 18264
rect 47124 16584 47176 16590
rect 47124 16526 47176 16532
rect 46768 11614 46888 11642
rect 46768 11150 46796 11614
rect 46848 11552 46900 11558
rect 46848 11494 46900 11500
rect 46756 11144 46808 11150
rect 46756 11086 46808 11092
rect 46664 10124 46716 10130
rect 46664 10066 46716 10072
rect 46676 9722 46704 10066
rect 46664 9716 46716 9722
rect 46664 9658 46716 9664
rect 46584 9574 46704 9602
rect 46572 8424 46624 8430
rect 46572 8366 46624 8372
rect 46584 7954 46612 8366
rect 46676 7954 46704 9574
rect 46768 9178 46796 11086
rect 46860 11082 46888 11494
rect 46848 11076 46900 11082
rect 46848 11018 46900 11024
rect 46848 10668 46900 10674
rect 46848 10610 46900 10616
rect 46860 10062 46888 10610
rect 46848 10056 46900 10062
rect 46848 9998 46900 10004
rect 46938 9480 46994 9489
rect 46938 9415 46994 9424
rect 46756 9172 46808 9178
rect 46756 9114 46808 9120
rect 46848 8968 46900 8974
rect 46848 8910 46900 8916
rect 46572 7948 46624 7954
rect 46572 7890 46624 7896
rect 46664 7948 46716 7954
rect 46664 7890 46716 7896
rect 46676 6866 46704 7890
rect 46756 7812 46808 7818
rect 46756 7754 46808 7760
rect 46664 6860 46716 6866
rect 46664 6802 46716 6808
rect 46768 6458 46796 7754
rect 46756 6452 46808 6458
rect 46756 6394 46808 6400
rect 46768 5166 46796 6394
rect 46860 6322 46888 8910
rect 46848 6316 46900 6322
rect 46848 6258 46900 6264
rect 46756 5160 46808 5166
rect 46756 5102 46808 5108
rect 46860 4078 46888 6258
rect 46848 4072 46900 4078
rect 46848 4014 46900 4020
rect 46846 3768 46902 3777
rect 46846 3703 46902 3712
rect 46860 3602 46888 3703
rect 46848 3596 46900 3602
rect 46848 3538 46900 3544
rect 46756 3460 46808 3466
rect 46756 3402 46808 3408
rect 46480 3188 46532 3194
rect 46480 3130 46532 3136
rect 46204 3052 46256 3058
rect 46204 2994 46256 3000
rect 45756 2746 46152 2774
rect 46124 2650 46152 2746
rect 46112 2644 46164 2650
rect 46112 2586 46164 2592
rect 45928 2372 45980 2378
rect 45928 2314 45980 2320
rect 45940 800 45968 2314
rect 46216 800 46244 2994
rect 46480 2440 46532 2446
rect 46480 2382 46532 2388
rect 46492 800 46520 2382
rect 46768 800 46796 3402
rect 46952 1358 46980 9415
rect 47032 3936 47084 3942
rect 47032 3878 47084 3884
rect 47044 3738 47072 3878
rect 47032 3732 47084 3738
rect 47032 3674 47084 3680
rect 47032 3052 47084 3058
rect 47032 2994 47084 3000
rect 46940 1352 46992 1358
rect 46940 1294 46992 1300
rect 47044 800 47072 2994
rect 47136 2650 47164 16526
rect 47216 15904 47268 15910
rect 47216 15846 47268 15852
rect 47228 3618 47256 15846
rect 47320 3942 47348 28358
rect 47492 26988 47544 26994
rect 47492 26930 47544 26936
rect 47400 15700 47452 15706
rect 47400 15642 47452 15648
rect 47412 9738 47440 15642
rect 47504 12434 47532 26930
rect 47596 23526 47624 40326
rect 49976 37120 50028 37126
rect 49976 37062 50028 37068
rect 49988 36650 50016 37062
rect 49976 36644 50028 36650
rect 49976 36586 50028 36592
rect 48964 35556 49016 35562
rect 48964 35498 49016 35504
rect 47676 35284 47728 35290
rect 47676 35226 47728 35232
rect 47688 23526 47716 35226
rect 48872 25696 48924 25702
rect 48872 25638 48924 25644
rect 47860 23588 47912 23594
rect 47860 23530 47912 23536
rect 47584 23520 47636 23526
rect 47584 23462 47636 23468
rect 47676 23520 47728 23526
rect 47676 23462 47728 23468
rect 47872 22094 47900 23530
rect 48596 23520 48648 23526
rect 48596 23462 48648 23468
rect 47872 22066 47992 22094
rect 47860 20936 47912 20942
rect 47860 20878 47912 20884
rect 47676 20868 47728 20874
rect 47676 20810 47728 20816
rect 47688 19922 47716 20810
rect 47676 19916 47728 19922
rect 47676 19858 47728 19864
rect 47584 19372 47636 19378
rect 47584 19314 47636 19320
rect 47596 18698 47624 19314
rect 47688 19174 47716 19858
rect 47872 19378 47900 20878
rect 47860 19372 47912 19378
rect 47860 19314 47912 19320
rect 47676 19168 47728 19174
rect 47676 19110 47728 19116
rect 47584 18692 47636 18698
rect 47584 18634 47636 18640
rect 47596 16522 47624 18634
rect 47688 17610 47716 19110
rect 47872 18766 47900 19314
rect 47860 18760 47912 18766
rect 47860 18702 47912 18708
rect 47676 17604 47728 17610
rect 47676 17546 47728 17552
rect 47584 16516 47636 16522
rect 47584 16458 47636 16464
rect 47768 15904 47820 15910
rect 47768 15846 47820 15852
rect 47780 14346 47808 15846
rect 47768 14340 47820 14346
rect 47768 14282 47820 14288
rect 47504 12406 47808 12434
rect 47412 9710 47716 9738
rect 47308 3936 47360 3942
rect 47308 3878 47360 3884
rect 47492 3936 47544 3942
rect 47492 3878 47544 3884
rect 47400 3664 47452 3670
rect 47228 3612 47400 3618
rect 47504 3641 47532 3878
rect 47228 3606 47452 3612
rect 47490 3632 47546 3641
rect 47228 3590 47440 3606
rect 47490 3567 47546 3576
rect 47584 3528 47636 3534
rect 47584 3470 47636 3476
rect 47124 2644 47176 2650
rect 47124 2586 47176 2592
rect 47308 2372 47360 2378
rect 47308 2314 47360 2320
rect 47320 800 47348 2314
rect 47596 800 47624 3470
rect 47688 2990 47716 9710
rect 47676 2984 47728 2990
rect 47676 2926 47728 2932
rect 47780 2650 47808 12406
rect 47858 8120 47914 8129
rect 47858 8055 47914 8064
rect 47872 3738 47900 8055
rect 47860 3732 47912 3738
rect 47860 3674 47912 3680
rect 47964 3194 47992 22066
rect 48228 20800 48280 20806
rect 48228 20742 48280 20748
rect 48136 20392 48188 20398
rect 48136 20334 48188 20340
rect 48148 18222 48176 20334
rect 48240 19854 48268 20742
rect 48412 20460 48464 20466
rect 48412 20402 48464 20408
rect 48424 19990 48452 20402
rect 48412 19984 48464 19990
rect 48412 19926 48464 19932
rect 48228 19848 48280 19854
rect 48228 19790 48280 19796
rect 48320 19780 48372 19786
rect 48320 19722 48372 19728
rect 48228 19372 48280 19378
rect 48228 19314 48280 19320
rect 48136 18216 48188 18222
rect 48136 18158 48188 18164
rect 48148 15978 48176 18158
rect 48240 17678 48268 19314
rect 48332 19310 48360 19722
rect 48320 19304 48372 19310
rect 48320 19246 48372 19252
rect 48332 18766 48360 19246
rect 48320 18760 48372 18766
rect 48320 18702 48372 18708
rect 48504 18760 48556 18766
rect 48504 18702 48556 18708
rect 48516 17882 48544 18702
rect 48504 17876 48556 17882
rect 48504 17818 48556 17824
rect 48228 17672 48280 17678
rect 48228 17614 48280 17620
rect 48320 17672 48372 17678
rect 48320 17614 48372 17620
rect 48332 17066 48360 17614
rect 48320 17060 48372 17066
rect 48320 17002 48372 17008
rect 48228 16040 48280 16046
rect 48228 15982 48280 15988
rect 48136 15972 48188 15978
rect 48136 15914 48188 15920
rect 48148 15366 48176 15914
rect 48136 15360 48188 15366
rect 48136 15302 48188 15308
rect 48148 14414 48176 15302
rect 48240 14618 48268 15982
rect 48320 14884 48372 14890
rect 48320 14826 48372 14832
rect 48332 14618 48360 14826
rect 48228 14612 48280 14618
rect 48228 14554 48280 14560
rect 48320 14612 48372 14618
rect 48320 14554 48372 14560
rect 48136 14408 48188 14414
rect 48136 14350 48188 14356
rect 48240 6798 48268 14554
rect 48412 13456 48464 13462
rect 48412 13398 48464 13404
rect 48320 11552 48372 11558
rect 48320 11494 48372 11500
rect 48228 6792 48280 6798
rect 48228 6734 48280 6740
rect 48332 5914 48360 11494
rect 48320 5908 48372 5914
rect 48320 5850 48372 5856
rect 48136 4140 48188 4146
rect 48136 4082 48188 4088
rect 47952 3188 48004 3194
rect 47952 3130 48004 3136
rect 47860 2848 47912 2854
rect 47860 2790 47912 2796
rect 47768 2644 47820 2650
rect 47768 2586 47820 2592
rect 47872 800 47900 2790
rect 48148 800 48176 4082
rect 48424 4010 48452 13398
rect 48412 4004 48464 4010
rect 48412 3946 48464 3952
rect 48608 3738 48636 23462
rect 48688 22772 48740 22778
rect 48688 22714 48740 22720
rect 48596 3732 48648 3738
rect 48596 3674 48648 3680
rect 48412 3052 48464 3058
rect 48412 2994 48464 3000
rect 48424 800 48452 2994
rect 48700 2650 48728 22714
rect 48780 18624 48832 18630
rect 48780 18566 48832 18572
rect 48792 18290 48820 18566
rect 48780 18284 48832 18290
rect 48780 18226 48832 18232
rect 48780 10260 48832 10266
rect 48780 10202 48832 10208
rect 48792 6866 48820 10202
rect 48780 6860 48832 6866
rect 48780 6802 48832 6808
rect 48792 5234 48820 6802
rect 48780 5228 48832 5234
rect 48780 5170 48832 5176
rect 48780 3528 48832 3534
rect 48780 3470 48832 3476
rect 48688 2644 48740 2650
rect 48688 2586 48740 2592
rect 48792 1034 48820 3470
rect 48884 3194 48912 25638
rect 48976 12434 49004 35498
rect 49148 31816 49200 31822
rect 49148 31758 49200 31764
rect 49056 29300 49108 29306
rect 49056 29242 49108 29248
rect 49068 13802 49096 29242
rect 49160 20874 49188 31758
rect 49792 31136 49844 31142
rect 49792 31078 49844 31084
rect 49516 23588 49568 23594
rect 49516 23530 49568 23536
rect 49148 20868 49200 20874
rect 49148 20810 49200 20816
rect 49160 20602 49188 20810
rect 49148 20596 49200 20602
rect 49148 20538 49200 20544
rect 49528 19718 49556 23530
rect 49700 19848 49752 19854
rect 49700 19790 49752 19796
rect 49516 19712 49568 19718
rect 49516 19654 49568 19660
rect 49712 18698 49740 19790
rect 49700 18692 49752 18698
rect 49700 18634 49752 18640
rect 49608 18284 49660 18290
rect 49608 18226 49660 18232
rect 49620 18086 49648 18226
rect 49608 18080 49660 18086
rect 49608 18022 49660 18028
rect 49620 17610 49648 18022
rect 49608 17604 49660 17610
rect 49608 17546 49660 17552
rect 49056 13796 49108 13802
rect 49056 13738 49108 13744
rect 48976 12406 49096 12434
rect 48872 3188 48924 3194
rect 48872 3130 48924 3136
rect 48964 3052 49016 3058
rect 48964 2994 49016 3000
rect 48700 1006 48820 1034
rect 48700 800 48728 1006
rect 48976 800 49004 2994
rect 49068 2650 49096 12406
rect 49424 10804 49476 10810
rect 49424 10746 49476 10752
rect 49436 3738 49464 10746
rect 49424 3732 49476 3738
rect 49424 3674 49476 3680
rect 49332 3528 49384 3534
rect 49332 3470 49384 3476
rect 49344 3126 49372 3470
rect 49804 3194 49832 31078
rect 50172 26234 50200 55186
rect 50294 54428 50602 54437
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54363 50602 54372
rect 50294 53340 50602 53349
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53275 50602 53284
rect 50294 52252 50602 52261
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52187 50602 52196
rect 50294 51164 50602 51173
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51099 50602 51108
rect 50294 50076 50602 50085
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50011 50602 50020
rect 50294 48988 50602 48997
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48923 50602 48932
rect 50294 47900 50602 47909
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47835 50602 47844
rect 50294 46812 50602 46821
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46747 50602 46756
rect 50294 45724 50602 45733
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45659 50602 45668
rect 50294 44636 50602 44645
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44571 50602 44580
rect 50294 43548 50602 43557
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43483 50602 43492
rect 50294 42460 50602 42469
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42395 50602 42404
rect 50294 41372 50602 41381
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41307 50602 41316
rect 50294 40284 50602 40293
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40219 50602 40228
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 50712 39092 50764 39098
rect 50712 39034 50764 39040
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 50724 35894 50752 39034
rect 50724 35866 50844 35894
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 50080 26206 50200 26234
rect 49974 20088 50030 20097
rect 49974 20023 50030 20032
rect 49988 19718 50016 20023
rect 49976 19712 50028 19718
rect 49976 19654 50028 19660
rect 50080 18358 50108 26206
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 50712 20868 50764 20874
rect 50712 20810 50764 20816
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 50528 20460 50580 20466
rect 50528 20402 50580 20408
rect 50158 19816 50214 19825
rect 50158 19751 50214 19760
rect 50172 19378 50200 19751
rect 50540 19700 50568 20402
rect 50724 19854 50752 20810
rect 50712 19848 50764 19854
rect 50710 19816 50712 19825
rect 50764 19816 50766 19825
rect 50710 19751 50766 19760
rect 50712 19712 50764 19718
rect 50540 19672 50660 19700
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 50160 19372 50212 19378
rect 50160 19314 50212 19320
rect 50632 19174 50660 19672
rect 50712 19654 50764 19660
rect 50724 19378 50752 19654
rect 50712 19372 50764 19378
rect 50712 19314 50764 19320
rect 50620 19168 50672 19174
rect 50620 19110 50672 19116
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 50068 18352 50120 18358
rect 50068 18294 50120 18300
rect 50620 17604 50672 17610
rect 50620 17546 50672 17552
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 50632 16658 50660 17546
rect 50816 17252 50844 35866
rect 51632 35080 51684 35086
rect 51632 35022 51684 35028
rect 50988 27056 51040 27062
rect 50988 26998 51040 27004
rect 51000 22094 51028 26998
rect 50724 17224 50844 17252
rect 50908 22066 51028 22094
rect 50620 16652 50672 16658
rect 50620 16594 50672 16600
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 50724 11830 50752 17224
rect 50908 12434 50936 22066
rect 50988 21344 51040 21350
rect 50988 21286 51040 21292
rect 51000 20262 51028 21286
rect 51448 20528 51500 20534
rect 51448 20470 51500 20476
rect 50988 20256 51040 20262
rect 50988 20198 51040 20204
rect 51460 19922 51488 20470
rect 51644 20330 51672 35022
rect 51736 29714 51764 56714
rect 53208 47598 53236 60998
rect 53932 60172 53984 60178
rect 53932 60114 53984 60120
rect 53380 47796 53432 47802
rect 53380 47738 53432 47744
rect 53196 47592 53248 47598
rect 53196 47534 53248 47540
rect 53196 35216 53248 35222
rect 53196 35158 53248 35164
rect 51724 29708 51776 29714
rect 51724 29650 51776 29656
rect 53208 22094 53236 35158
rect 53208 22066 53328 22094
rect 52736 21412 52788 21418
rect 52736 21354 52788 21360
rect 53196 21412 53248 21418
rect 53196 21354 53248 21360
rect 52092 21344 52144 21350
rect 52092 21286 52144 21292
rect 52104 21010 52132 21286
rect 52092 21004 52144 21010
rect 52092 20946 52144 20952
rect 51632 20324 51684 20330
rect 51632 20266 51684 20272
rect 51644 20097 51672 20266
rect 51630 20088 51686 20097
rect 51630 20023 51686 20032
rect 51080 19916 51132 19922
rect 51080 19858 51132 19864
rect 51448 19916 51500 19922
rect 51448 19858 51500 19864
rect 51092 19378 51120 19858
rect 51264 19712 51316 19718
rect 51264 19654 51316 19660
rect 51172 19440 51224 19446
rect 51276 19428 51304 19654
rect 51224 19400 51304 19428
rect 51172 19382 51224 19388
rect 51080 19372 51132 19378
rect 51080 19314 51132 19320
rect 51368 19310 51396 19341
rect 51356 19304 51408 19310
rect 51540 19304 51592 19310
rect 51408 19252 51540 19258
rect 51356 19246 51592 19252
rect 51368 19230 51580 19246
rect 51368 18766 51396 19230
rect 51356 18760 51408 18766
rect 51356 18702 51408 18708
rect 51080 17672 51132 17678
rect 51080 17614 51132 17620
rect 50988 16652 51040 16658
rect 50988 16594 51040 16600
rect 51000 15722 51028 16594
rect 51092 16114 51120 17614
rect 51170 17232 51226 17241
rect 51368 17202 51396 18702
rect 51724 17604 51776 17610
rect 51724 17546 51776 17552
rect 51540 17536 51592 17542
rect 51540 17478 51592 17484
rect 51552 17202 51580 17478
rect 51736 17338 51764 17546
rect 51724 17332 51776 17338
rect 51724 17274 51776 17280
rect 51170 17167 51172 17176
rect 51224 17167 51226 17176
rect 51356 17196 51408 17202
rect 51172 17138 51224 17144
rect 51356 17138 51408 17144
rect 51540 17196 51592 17202
rect 51540 17138 51592 17144
rect 52104 17134 52132 20946
rect 52748 20942 52776 21354
rect 53208 21078 53236 21354
rect 53196 21072 53248 21078
rect 53196 21014 53248 21020
rect 52736 20936 52788 20942
rect 52736 20878 52788 20884
rect 53104 20936 53156 20942
rect 53104 20878 53156 20884
rect 53116 20262 53144 20878
rect 53104 20256 53156 20262
rect 53104 20198 53156 20204
rect 52276 19780 52328 19786
rect 52276 19722 52328 19728
rect 52288 19378 52316 19722
rect 52460 19440 52512 19446
rect 52460 19382 52512 19388
rect 52276 19372 52328 19378
rect 52276 19314 52328 19320
rect 52184 18080 52236 18086
rect 52184 18022 52236 18028
rect 51448 17128 51500 17134
rect 51448 17070 51500 17076
rect 52092 17128 52144 17134
rect 52092 17070 52144 17076
rect 51356 16584 51408 16590
rect 51460 16572 51488 17070
rect 51408 16544 51488 16572
rect 51540 16584 51592 16590
rect 51356 16526 51408 16532
rect 51540 16526 51592 16532
rect 51080 16108 51132 16114
rect 51080 16050 51132 16056
rect 51172 15904 51224 15910
rect 51172 15846 51224 15852
rect 51184 15722 51212 15846
rect 51000 15694 51212 15722
rect 51184 15502 51212 15694
rect 51172 15496 51224 15502
rect 51172 15438 51224 15444
rect 50908 12406 51028 12434
rect 50712 11824 50764 11830
rect 50712 11766 50764 11772
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 50712 4752 50764 4758
rect 50712 4694 50764 4700
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 49884 3460 49936 3466
rect 49884 3402 49936 3408
rect 50620 3460 50672 3466
rect 50620 3402 50672 3408
rect 49792 3188 49844 3194
rect 49792 3130 49844 3136
rect 49332 3120 49384 3126
rect 49332 3062 49384 3068
rect 49516 3120 49568 3126
rect 49516 3062 49568 3068
rect 49056 2644 49108 2650
rect 49056 2586 49108 2592
rect 49240 2508 49292 2514
rect 49240 2450 49292 2456
rect 49252 800 49280 2450
rect 49528 800 49556 3062
rect 49608 2916 49660 2922
rect 49608 2858 49660 2864
rect 49700 2916 49752 2922
rect 49700 2858 49752 2864
rect 49620 2825 49648 2858
rect 49606 2816 49662 2825
rect 49606 2751 49662 2760
rect 49712 2446 49740 2858
rect 49896 2774 49924 3402
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 50160 3052 50212 3058
rect 50160 2994 50212 3000
rect 49804 2746 49924 2774
rect 49700 2440 49752 2446
rect 49700 2382 49752 2388
rect 49804 800 49832 2746
rect 50068 2304 50120 2310
rect 50068 2246 50120 2252
rect 50080 800 50108 2246
rect 50172 1442 50200 2994
rect 50436 2848 50488 2854
rect 50528 2848 50580 2854
rect 50436 2790 50488 2796
rect 50526 2816 50528 2825
rect 50580 2816 50582 2825
rect 50448 2446 50476 2790
rect 50526 2751 50582 2760
rect 50436 2440 50488 2446
rect 50436 2382 50488 2388
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 50172 1414 50384 1442
rect 50356 800 50384 1414
rect 50632 800 50660 3402
rect 50724 3194 50752 4694
rect 50804 3392 50856 3398
rect 50804 3334 50856 3340
rect 50712 3188 50764 3194
rect 50712 3130 50764 3136
rect 50816 2922 50844 3334
rect 50896 3120 50948 3126
rect 50896 3062 50948 3068
rect 50804 2916 50856 2922
rect 50804 2858 50856 2864
rect 50712 2576 50764 2582
rect 50712 2518 50764 2524
rect 50724 2106 50752 2518
rect 50712 2100 50764 2106
rect 50712 2042 50764 2048
rect 50908 800 50936 3062
rect 51000 2514 51028 12406
rect 51368 6390 51396 16526
rect 51552 15706 51580 16526
rect 51724 16448 51776 16454
rect 51724 16390 51776 16396
rect 51736 16182 51764 16390
rect 51724 16176 51776 16182
rect 51724 16118 51776 16124
rect 51540 15700 51592 15706
rect 51540 15642 51592 15648
rect 51724 9920 51776 9926
rect 51724 9862 51776 9868
rect 51356 6384 51408 6390
rect 51356 6326 51408 6332
rect 51368 5930 51396 6326
rect 51276 5902 51396 5930
rect 51276 4622 51304 5902
rect 51448 5024 51500 5030
rect 51448 4966 51500 4972
rect 51460 4622 51488 4966
rect 51264 4616 51316 4622
rect 51264 4558 51316 4564
rect 51448 4616 51500 4622
rect 51448 4558 51500 4564
rect 51736 4146 51764 9862
rect 52000 4208 52052 4214
rect 52000 4150 52052 4156
rect 51724 4140 51776 4146
rect 51724 4082 51776 4088
rect 51724 3528 51776 3534
rect 51724 3470 51776 3476
rect 51264 3460 51316 3466
rect 51264 3402 51316 3408
rect 50988 2508 51040 2514
rect 50988 2450 51040 2456
rect 51276 2394 51304 3402
rect 51448 3052 51500 3058
rect 51448 2994 51500 3000
rect 51184 2366 51304 2394
rect 51184 800 51212 2366
rect 51264 2304 51316 2310
rect 51264 2246 51316 2252
rect 51276 1970 51304 2246
rect 51264 1964 51316 1970
rect 51264 1906 51316 1912
rect 51460 800 51488 2994
rect 51736 800 51764 3470
rect 52012 800 52040 4150
rect 52196 3194 52224 18022
rect 52472 17678 52500 19382
rect 52460 17672 52512 17678
rect 52460 17614 52512 17620
rect 52368 17604 52420 17610
rect 52368 17546 52420 17552
rect 52276 17332 52328 17338
rect 52276 17274 52328 17280
rect 52288 16794 52316 17274
rect 52380 17270 52408 17546
rect 52472 17270 52500 17614
rect 53104 17536 53156 17542
rect 53104 17478 53156 17484
rect 52368 17264 52420 17270
rect 52368 17206 52420 17212
rect 52460 17264 52512 17270
rect 52460 17206 52512 17212
rect 52472 16794 52500 17206
rect 52276 16788 52328 16794
rect 52276 16730 52328 16736
rect 52460 16788 52512 16794
rect 52460 16730 52512 16736
rect 53116 16590 53144 17478
rect 53104 16584 53156 16590
rect 53104 16526 53156 16532
rect 52368 15904 52420 15910
rect 52368 15846 52420 15852
rect 52380 15502 52408 15846
rect 52368 15496 52420 15502
rect 52368 15438 52420 15444
rect 52460 14816 52512 14822
rect 52460 14758 52512 14764
rect 52472 7546 52500 14758
rect 53116 8566 53144 16526
rect 53104 8560 53156 8566
rect 53104 8502 53156 8508
rect 52460 7540 52512 7546
rect 52460 7482 52512 7488
rect 53104 4684 53156 4690
rect 53104 4626 53156 4632
rect 53116 4282 53144 4626
rect 52460 4276 52512 4282
rect 52460 4218 52512 4224
rect 53104 4276 53156 4282
rect 53104 4218 53156 4224
rect 52472 3738 52500 4218
rect 52828 4208 52880 4214
rect 52828 4150 52880 4156
rect 52460 3732 52512 3738
rect 52460 3674 52512 3680
rect 52276 3460 52328 3466
rect 52276 3402 52328 3408
rect 52184 3188 52236 3194
rect 52184 3130 52236 3136
rect 52288 800 52316 3402
rect 52552 2372 52604 2378
rect 52552 2314 52604 2320
rect 52564 800 52592 2314
rect 52840 800 52868 4150
rect 53196 3528 53248 3534
rect 53196 3470 53248 3476
rect 53104 2304 53156 2310
rect 53104 2246 53156 2252
rect 53116 1902 53144 2246
rect 53104 1896 53156 1902
rect 53104 1838 53156 1844
rect 53208 1714 53236 3470
rect 53300 2990 53328 22066
rect 53392 10742 53420 47738
rect 53840 37256 53892 37262
rect 53840 37198 53892 37204
rect 53656 36780 53708 36786
rect 53656 36722 53708 36728
rect 53380 10736 53432 10742
rect 53380 10678 53432 10684
rect 53472 10668 53524 10674
rect 53472 10610 53524 10616
rect 53484 10470 53512 10610
rect 53472 10464 53524 10470
rect 53472 10406 53524 10412
rect 53564 4480 53616 4486
rect 53564 4422 53616 4428
rect 53380 4208 53432 4214
rect 53380 4150 53432 4156
rect 53288 2984 53340 2990
rect 53288 2926 53340 2932
rect 53116 1686 53236 1714
rect 53116 800 53144 1686
rect 53392 800 53420 4150
rect 53472 4072 53524 4078
rect 53472 4014 53524 4020
rect 53484 2922 53512 4014
rect 53576 3466 53604 4422
rect 53668 4010 53696 36722
rect 53852 36582 53880 37198
rect 53944 36854 53972 60114
rect 54116 59968 54168 59974
rect 54116 59910 54168 59916
rect 54128 37262 54156 59910
rect 54312 42634 54340 60998
rect 54680 60722 54708 63294
rect 55310 63294 55536 63322
rect 55310 63200 55366 63294
rect 55402 61568 55458 61577
rect 55402 61503 55458 61512
rect 55416 60722 55444 61503
rect 55508 61198 55536 63294
rect 56046 63200 56102 64000
rect 56782 63322 56838 64000
rect 56782 63294 56916 63322
rect 56782 63200 56838 63294
rect 56060 61198 56088 63200
rect 56414 62656 56470 62665
rect 56414 62591 56470 62600
rect 56138 62112 56194 62121
rect 56138 62047 56194 62056
rect 55496 61192 55548 61198
rect 55496 61134 55548 61140
rect 56048 61192 56100 61198
rect 56048 61134 56100 61140
rect 55772 61124 55824 61130
rect 55772 61066 55824 61072
rect 54668 60716 54720 60722
rect 54668 60658 54720 60664
rect 55404 60716 55456 60722
rect 55404 60658 55456 60664
rect 54852 60512 54904 60518
rect 54852 60454 54904 60460
rect 55588 60512 55640 60518
rect 55588 60454 55640 60460
rect 54864 43382 54892 60454
rect 55600 60314 55628 60454
rect 55588 60308 55640 60314
rect 55588 60250 55640 60256
rect 55784 50386 55812 61066
rect 56152 60722 56180 62047
rect 56140 60716 56192 60722
rect 56140 60658 56192 60664
rect 56428 59702 56456 62591
rect 56692 61056 56744 61062
rect 56506 61024 56562 61033
rect 56692 60998 56744 61004
rect 56506 60959 56562 60968
rect 56520 60110 56548 60959
rect 56508 60104 56560 60110
rect 56508 60046 56560 60052
rect 56416 59696 56468 59702
rect 56416 59638 56468 59644
rect 56704 58546 56732 60998
rect 56888 60722 56916 63294
rect 57518 63200 57574 64000
rect 58254 63322 58310 64000
rect 57992 63294 58310 63322
rect 57532 61198 57560 63200
rect 57520 61192 57572 61198
rect 57520 61134 57572 61140
rect 56876 60716 56928 60722
rect 56876 60658 56928 60664
rect 57060 60512 57112 60518
rect 57060 60454 57112 60460
rect 57242 60480 57298 60489
rect 56692 58540 56744 58546
rect 56692 58482 56744 58488
rect 55772 50380 55824 50386
rect 55772 50322 55824 50328
rect 57072 45490 57100 60454
rect 57242 60415 57298 60424
rect 57256 60110 57284 60415
rect 57992 60110 58020 63294
rect 58254 63200 58310 63294
rect 58990 63200 59046 64000
rect 58072 60716 58124 60722
rect 58072 60658 58124 60664
rect 57244 60104 57296 60110
rect 57244 60046 57296 60052
rect 57980 60104 58032 60110
rect 57980 60046 58032 60052
rect 58084 59945 58112 60658
rect 58256 60512 58308 60518
rect 58256 60454 58308 60460
rect 58268 60217 58296 60454
rect 58254 60208 58310 60217
rect 58254 60143 58310 60152
rect 58256 60036 58308 60042
rect 58256 59978 58308 59984
rect 58070 59936 58126 59945
rect 58070 59871 58126 59880
rect 58072 59628 58124 59634
rect 58072 59570 58124 59576
rect 57152 59424 57204 59430
rect 58084 59401 58112 59570
rect 57152 59366 57204 59372
rect 58070 59392 58126 59401
rect 57164 59022 57192 59366
rect 58070 59327 58126 59336
rect 58072 59084 58124 59090
rect 58072 59026 58124 59032
rect 57152 59016 57204 59022
rect 57152 58958 57204 58964
rect 57888 59016 57940 59022
rect 58084 58993 58112 59026
rect 57888 58958 57940 58964
rect 58070 58984 58126 58993
rect 57900 58313 57928 58958
rect 58070 58919 58126 58928
rect 58162 58848 58218 58857
rect 58162 58783 58218 58792
rect 58176 58614 58204 58783
rect 58164 58608 58216 58614
rect 58164 58550 58216 58556
rect 57886 58304 57942 58313
rect 57886 58239 57942 58248
rect 57980 57860 58032 57866
rect 57980 57802 58032 57808
rect 57992 57769 58020 57802
rect 58072 57792 58124 57798
rect 57978 57760 58034 57769
rect 58072 57734 58124 57740
rect 57978 57695 58034 57704
rect 57886 57216 57942 57225
rect 57886 57151 57942 57160
rect 57900 56846 57928 57151
rect 57888 56840 57940 56846
rect 57888 56782 57940 56788
rect 57428 50312 57480 50318
rect 57428 50254 57480 50260
rect 57060 45484 57112 45490
rect 57060 45426 57112 45432
rect 56784 44872 56836 44878
rect 56784 44814 56836 44820
rect 54852 43376 54904 43382
rect 54852 43318 54904 43324
rect 54300 42628 54352 42634
rect 54300 42570 54352 42576
rect 54668 41608 54720 41614
rect 54668 41550 54720 41556
rect 54208 37460 54260 37466
rect 54208 37402 54260 37408
rect 54116 37256 54168 37262
rect 54116 37198 54168 37204
rect 54024 37188 54076 37194
rect 54024 37130 54076 37136
rect 53932 36848 53984 36854
rect 53932 36790 53984 36796
rect 54036 36650 54064 37130
rect 54220 36650 54248 37402
rect 54300 37256 54352 37262
rect 54300 37198 54352 37204
rect 54484 37256 54536 37262
rect 54484 37198 54536 37204
rect 54024 36644 54076 36650
rect 54024 36586 54076 36592
rect 54208 36644 54260 36650
rect 54208 36586 54260 36592
rect 53840 36576 53892 36582
rect 53840 36518 53892 36524
rect 53840 19848 53892 19854
rect 53840 19790 53892 19796
rect 53852 18902 53880 19790
rect 53840 18896 53892 18902
rect 53840 18838 53892 18844
rect 53932 18828 53984 18834
rect 53932 18770 53984 18776
rect 53840 18692 53892 18698
rect 53840 18634 53892 18640
rect 53852 18426 53880 18634
rect 53944 18426 53972 18770
rect 53840 18420 53892 18426
rect 53840 18362 53892 18368
rect 53932 18420 53984 18426
rect 53932 18362 53984 18368
rect 53932 17128 53984 17134
rect 53930 17096 53932 17105
rect 53984 17096 53986 17105
rect 53930 17031 53986 17040
rect 53748 16244 53800 16250
rect 53748 16186 53800 16192
rect 53760 15910 53788 16186
rect 53932 16108 53984 16114
rect 53932 16050 53984 16056
rect 53748 15904 53800 15910
rect 53748 15846 53800 15852
rect 53944 15570 53972 16050
rect 53932 15564 53984 15570
rect 53932 15506 53984 15512
rect 54036 10810 54064 36586
rect 54312 26234 54340 37198
rect 54220 26206 54340 26234
rect 54116 21004 54168 21010
rect 54116 20946 54168 20952
rect 54128 20466 54156 20946
rect 54116 20460 54168 20466
rect 54116 20402 54168 20408
rect 54116 16992 54168 16998
rect 54116 16934 54168 16940
rect 54128 16250 54156 16934
rect 54116 16244 54168 16250
rect 54116 16186 54168 16192
rect 54220 12434 54248 26206
rect 54496 20942 54524 37198
rect 54484 20936 54536 20942
rect 54484 20878 54536 20884
rect 54496 20602 54524 20878
rect 54484 20596 54536 20602
rect 54484 20538 54536 20544
rect 54392 20256 54444 20262
rect 54392 20198 54444 20204
rect 54300 19848 54352 19854
rect 54300 19790 54352 19796
rect 54312 19446 54340 19790
rect 54300 19440 54352 19446
rect 54300 19382 54352 19388
rect 54404 18154 54432 20198
rect 54576 19916 54628 19922
rect 54576 19858 54628 19864
rect 54588 18290 54616 19858
rect 54680 19718 54708 41550
rect 55036 36576 55088 36582
rect 55036 36518 55088 36524
rect 54944 24132 54996 24138
rect 54944 24074 54996 24080
rect 54760 20936 54812 20942
rect 54760 20878 54812 20884
rect 54852 20936 54904 20942
rect 54852 20878 54904 20884
rect 54772 20058 54800 20878
rect 54760 20052 54812 20058
rect 54760 19994 54812 20000
rect 54668 19712 54720 19718
rect 54668 19654 54720 19660
rect 54576 18284 54628 18290
rect 54576 18226 54628 18232
rect 54392 18148 54444 18154
rect 54392 18090 54444 18096
rect 54298 17232 54354 17241
rect 54298 17167 54300 17176
rect 54352 17167 54354 17176
rect 54300 17138 54352 17144
rect 54300 16992 54352 16998
rect 54300 16934 54352 16940
rect 54312 16590 54340 16934
rect 54300 16584 54352 16590
rect 54300 16526 54352 16532
rect 54404 16114 54432 18090
rect 54588 17814 54616 18226
rect 54576 17808 54628 17814
rect 54576 17750 54628 17756
rect 54576 17672 54628 17678
rect 54576 17614 54628 17620
rect 54588 16522 54616 17614
rect 54668 17332 54720 17338
rect 54668 17274 54720 17280
rect 54760 17332 54812 17338
rect 54760 17274 54812 17280
rect 54680 16726 54708 17274
rect 54668 16720 54720 16726
rect 54668 16662 54720 16668
rect 54576 16516 54628 16522
rect 54576 16458 54628 16464
rect 54588 16114 54616 16458
rect 54772 16250 54800 17274
rect 54760 16244 54812 16250
rect 54760 16186 54812 16192
rect 54392 16108 54444 16114
rect 54392 16050 54444 16056
rect 54576 16108 54628 16114
rect 54576 16050 54628 16056
rect 54772 16046 54800 16186
rect 54760 16040 54812 16046
rect 54760 15982 54812 15988
rect 54864 14958 54892 20878
rect 54852 14952 54904 14958
rect 54852 14894 54904 14900
rect 54220 12406 54340 12434
rect 54024 10804 54076 10810
rect 54024 10746 54076 10752
rect 54312 10674 54340 12406
rect 54300 10668 54352 10674
rect 54300 10610 54352 10616
rect 54208 10600 54260 10606
rect 54208 10542 54260 10548
rect 53656 4004 53708 4010
rect 53656 3946 53708 3952
rect 54220 3738 54248 10542
rect 54484 4140 54536 4146
rect 54484 4082 54536 4088
rect 54208 3732 54260 3738
rect 54208 3674 54260 3680
rect 53564 3460 53616 3466
rect 53564 3402 53616 3408
rect 53932 3052 53984 3058
rect 53932 2994 53984 3000
rect 54208 3052 54260 3058
rect 54208 2994 54260 3000
rect 53472 2916 53524 2922
rect 53472 2858 53524 2864
rect 53656 2440 53708 2446
rect 53656 2382 53708 2388
rect 53668 800 53696 2382
rect 53944 800 53972 2994
rect 54220 800 54248 2994
rect 54496 800 54524 4082
rect 54760 3528 54812 3534
rect 54760 3470 54812 3476
rect 54772 800 54800 3470
rect 54956 3126 54984 24074
rect 55048 22094 55076 36518
rect 56140 32904 56192 32910
rect 56140 32846 56192 32852
rect 55864 32768 55916 32774
rect 55864 32710 55916 32716
rect 55588 28552 55640 28558
rect 55588 28494 55640 28500
rect 55048 22066 55168 22094
rect 55036 18828 55088 18834
rect 55036 18770 55088 18776
rect 55048 18426 55076 18770
rect 55036 18420 55088 18426
rect 55036 18362 55088 18368
rect 55140 6914 55168 22066
rect 55312 21004 55364 21010
rect 55312 20946 55364 20952
rect 55220 20800 55272 20806
rect 55220 20742 55272 20748
rect 55232 20466 55260 20742
rect 55220 20460 55272 20466
rect 55220 20402 55272 20408
rect 55324 18766 55352 20946
rect 55312 18760 55364 18766
rect 55312 18702 55364 18708
rect 55600 17882 55628 28494
rect 55876 26926 55904 32710
rect 55864 26920 55916 26926
rect 55864 26862 55916 26868
rect 56048 20936 56100 20942
rect 56048 20878 56100 20884
rect 55680 20868 55732 20874
rect 55680 20810 55732 20816
rect 55692 19854 55720 20810
rect 55864 20256 55916 20262
rect 55864 20198 55916 20204
rect 55876 19854 55904 20198
rect 56060 20058 56088 20878
rect 56048 20052 56100 20058
rect 56048 19994 56100 20000
rect 55680 19848 55732 19854
rect 55680 19790 55732 19796
rect 55864 19848 55916 19854
rect 55864 19790 55916 19796
rect 55588 17876 55640 17882
rect 55588 17818 55640 17824
rect 55692 17338 55720 19790
rect 56152 19786 56180 32846
rect 56692 20800 56744 20806
rect 56692 20742 56744 20748
rect 56600 20596 56652 20602
rect 56600 20538 56652 20544
rect 56508 20528 56560 20534
rect 56508 20470 56560 20476
rect 56520 19922 56548 20470
rect 56508 19916 56560 19922
rect 56508 19858 56560 19864
rect 56140 19780 56192 19786
rect 56140 19722 56192 19728
rect 55864 18624 55916 18630
rect 55864 18566 55916 18572
rect 55876 18290 55904 18566
rect 56520 18358 56548 19858
rect 56612 19718 56640 20538
rect 56704 19854 56732 20742
rect 56692 19848 56744 19854
rect 56692 19790 56744 19796
rect 56600 19712 56652 19718
rect 56600 19654 56652 19660
rect 56600 18760 56652 18766
rect 56600 18702 56652 18708
rect 56508 18352 56560 18358
rect 56508 18294 56560 18300
rect 55864 18284 55916 18290
rect 55864 18226 55916 18232
rect 56520 17746 56548 18294
rect 56508 17740 56560 17746
rect 56508 17682 56560 17688
rect 56140 17604 56192 17610
rect 56140 17546 56192 17552
rect 56152 17338 56180 17546
rect 55680 17332 55732 17338
rect 55680 17274 55732 17280
rect 56140 17332 56192 17338
rect 56140 17274 56192 17280
rect 56048 17196 56100 17202
rect 56048 17138 56100 17144
rect 55772 17128 55824 17134
rect 55770 17096 55772 17105
rect 55824 17096 55826 17105
rect 55770 17031 55826 17040
rect 56060 16454 56088 17138
rect 56520 16794 56548 17682
rect 56508 16788 56560 16794
rect 56508 16730 56560 16736
rect 55220 16448 55272 16454
rect 55220 16390 55272 16396
rect 56048 16448 56100 16454
rect 56048 16390 56100 16396
rect 55232 16182 55260 16390
rect 55220 16176 55272 16182
rect 55220 16118 55272 16124
rect 56612 14618 56640 18702
rect 56600 14612 56652 14618
rect 56600 14554 56652 14560
rect 56796 14550 56824 44814
rect 57244 44804 57296 44810
rect 57244 44746 57296 44752
rect 57256 44713 57284 44746
rect 57242 44704 57298 44713
rect 57242 44639 57298 44648
rect 57060 42628 57112 42634
rect 57060 42570 57112 42576
rect 57072 42537 57100 42570
rect 57336 42560 57388 42566
rect 57058 42528 57114 42537
rect 57336 42502 57388 42508
rect 57058 42463 57114 42472
rect 57348 41585 57376 42502
rect 57334 41576 57390 41585
rect 57244 41540 57296 41546
rect 57334 41511 57390 41520
rect 57244 41482 57296 41488
rect 57256 41449 57284 41482
rect 57242 41440 57298 41449
rect 57242 41375 57298 41384
rect 57060 40452 57112 40458
rect 57060 40394 57112 40400
rect 57072 40361 57100 40394
rect 57058 40352 57114 40361
rect 57058 40287 57114 40296
rect 57060 39364 57112 39370
rect 57060 39306 57112 39312
rect 57072 39273 57100 39306
rect 57058 39264 57114 39273
rect 57058 39199 57114 39208
rect 57060 32836 57112 32842
rect 57060 32778 57112 32784
rect 57072 32745 57100 32778
rect 57058 32736 57114 32745
rect 57058 32671 57114 32680
rect 57152 29640 57204 29646
rect 57152 29582 57204 29588
rect 57060 29572 57112 29578
rect 57060 29514 57112 29520
rect 57072 29481 57100 29514
rect 57058 29472 57114 29481
rect 57058 29407 57114 29416
rect 57060 22024 57112 22030
rect 57060 21966 57112 21972
rect 57072 17882 57100 21966
rect 57164 18426 57192 29582
rect 57336 22092 57388 22098
rect 57336 22034 57388 22040
rect 57244 18692 57296 18698
rect 57244 18634 57296 18640
rect 57256 18601 57284 18634
rect 57242 18592 57298 18601
rect 57242 18527 57298 18536
rect 57152 18420 57204 18426
rect 57152 18362 57204 18368
rect 57060 17876 57112 17882
rect 57060 17818 57112 17824
rect 57072 17338 57100 17818
rect 57060 17332 57112 17338
rect 57060 17274 57112 17280
rect 57348 17218 57376 22034
rect 57256 17190 57376 17218
rect 57060 16516 57112 16522
rect 57060 16458 57112 16464
rect 56968 16448 57020 16454
rect 57072 16425 57100 16458
rect 57152 16448 57204 16454
rect 56968 16390 57020 16396
rect 57058 16416 57114 16425
rect 56980 16266 57008 16390
rect 57152 16390 57204 16396
rect 57058 16351 57114 16360
rect 56980 16238 57100 16266
rect 56784 14544 56836 14550
rect 56784 14486 56836 14492
rect 55220 13796 55272 13802
rect 55220 13738 55272 13744
rect 55048 6886 55168 6914
rect 55048 3738 55076 6886
rect 55036 3732 55088 3738
rect 55036 3674 55088 3680
rect 55232 3194 55260 13738
rect 56968 13320 57020 13326
rect 56968 13262 57020 13268
rect 55864 13252 55916 13258
rect 55864 13194 55916 13200
rect 55496 8288 55548 8294
rect 55496 8230 55548 8236
rect 55508 7886 55536 8230
rect 55496 7880 55548 7886
rect 55496 7822 55548 7828
rect 55772 7880 55824 7886
rect 55772 7822 55824 7828
rect 55784 7478 55812 7822
rect 55772 7472 55824 7478
rect 55772 7414 55824 7420
rect 55876 5710 55904 13194
rect 56980 13161 57008 13262
rect 56966 13152 57022 13161
rect 56966 13087 57022 13096
rect 56876 11144 56928 11150
rect 56876 11086 56928 11092
rect 56140 11076 56192 11082
rect 56140 11018 56192 11024
rect 56152 8974 56180 11018
rect 56508 10056 56560 10062
rect 56508 9998 56560 10004
rect 56324 9376 56376 9382
rect 56324 9318 56376 9324
rect 56336 8974 56364 9318
rect 56140 8968 56192 8974
rect 56140 8910 56192 8916
rect 56324 8968 56376 8974
rect 56324 8910 56376 8916
rect 55956 8016 56008 8022
rect 55956 7958 56008 7964
rect 55968 7410 55996 7958
rect 56152 7818 56180 8910
rect 56232 8492 56284 8498
rect 56232 8434 56284 8440
rect 56244 8265 56272 8434
rect 56520 8362 56548 9998
rect 56888 9042 56916 11086
rect 56968 11076 57020 11082
rect 56968 11018 57020 11024
rect 56980 10810 57008 11018
rect 56968 10804 57020 10810
rect 56968 10746 57020 10752
rect 57072 10674 57100 16238
rect 57164 15473 57192 16390
rect 57150 15464 57206 15473
rect 57150 15399 57206 15408
rect 57256 13870 57284 17190
rect 57336 17128 57388 17134
rect 57336 17070 57388 17076
rect 57348 16969 57376 17070
rect 57334 16960 57390 16969
rect 57334 16895 57390 16904
rect 57244 13864 57296 13870
rect 57244 13806 57296 13812
rect 57152 11756 57204 11762
rect 57152 11698 57204 11704
rect 57164 11529 57192 11698
rect 57440 11626 57468 50254
rect 57888 50176 57940 50182
rect 57888 50118 57940 50124
rect 57900 49609 57928 50118
rect 57886 49600 57942 49609
rect 57886 49535 57942 49544
rect 57980 49156 58032 49162
rect 57980 49098 58032 49104
rect 57992 49065 58020 49098
rect 57978 49056 58034 49065
rect 57978 48991 58034 49000
rect 57796 48136 57848 48142
rect 57796 48078 57848 48084
rect 57704 45960 57756 45966
rect 57704 45902 57756 45908
rect 57612 43784 57664 43790
rect 57612 43726 57664 43732
rect 57520 40520 57572 40526
rect 57520 40462 57572 40468
rect 57532 23594 57560 40462
rect 57520 23588 57572 23594
rect 57520 23530 57572 23536
rect 57624 18086 57652 43726
rect 57716 22098 57744 45902
rect 57704 22092 57756 22098
rect 57704 22034 57756 22040
rect 57808 21978 57836 48078
rect 58084 47802 58112 57734
rect 58162 56672 58218 56681
rect 58162 56607 58218 56616
rect 58176 56438 58204 56607
rect 58164 56432 58216 56438
rect 58164 56374 58216 56380
rect 58164 48068 58216 48074
rect 58164 48010 58216 48016
rect 58176 47977 58204 48010
rect 58162 47968 58218 47977
rect 58162 47903 58218 47912
rect 58072 47796 58124 47802
rect 58072 47738 58124 47744
rect 58072 47660 58124 47666
rect 58072 47602 58124 47608
rect 58084 47433 58112 47602
rect 58070 47424 58126 47433
rect 58070 47359 58126 47368
rect 58162 46336 58218 46345
rect 58162 46271 58218 46280
rect 58176 46034 58204 46271
rect 58164 46028 58216 46034
rect 58164 45970 58216 45976
rect 58070 45792 58126 45801
rect 58070 45727 58126 45736
rect 58084 45490 58112 45727
rect 58072 45484 58124 45490
rect 58072 45426 58124 45432
rect 57888 44804 57940 44810
rect 57888 44746 57940 44752
rect 57900 44169 57928 44746
rect 57886 44160 57942 44169
rect 57886 44095 57942 44104
rect 58164 43716 58216 43722
rect 58164 43658 58216 43664
rect 58176 43081 58204 43658
rect 58162 43072 58218 43081
rect 58162 43007 58218 43016
rect 57980 42628 58032 42634
rect 57980 42570 58032 42576
rect 57992 41993 58020 42570
rect 57978 41984 58034 41993
rect 57978 41919 58034 41928
rect 57888 41540 57940 41546
rect 57888 41482 57940 41488
rect 57900 40905 57928 41482
rect 57886 40896 57942 40905
rect 57886 40831 57942 40840
rect 57888 40384 57940 40390
rect 57888 40326 57940 40332
rect 57900 39817 57928 40326
rect 57886 39808 57942 39817
rect 57886 39743 57942 39752
rect 57980 39364 58032 39370
rect 57980 39306 58032 39312
rect 57992 38729 58020 39306
rect 58072 39296 58124 39302
rect 58072 39238 58124 39244
rect 58084 39098 58112 39238
rect 58072 39092 58124 39098
rect 58072 39034 58124 39040
rect 57978 38720 58034 38729
rect 57978 38655 58034 38664
rect 58164 38276 58216 38282
rect 58164 38218 58216 38224
rect 58176 38185 58204 38218
rect 58162 38176 58218 38185
rect 58162 38111 58218 38120
rect 58072 37868 58124 37874
rect 58072 37810 58124 37816
rect 58084 37641 58112 37810
rect 58070 37632 58126 37641
rect 58070 37567 58126 37576
rect 58164 37188 58216 37194
rect 58164 37130 58216 37136
rect 58176 36553 58204 37130
rect 58162 36544 58218 36553
rect 58162 36479 58218 36488
rect 57980 36100 58032 36106
rect 57980 36042 58032 36048
rect 57992 36009 58020 36042
rect 57978 36000 58034 36009
rect 57978 35935 58034 35944
rect 58164 35012 58216 35018
rect 58164 34954 58216 34960
rect 58176 34921 58204 34954
rect 58162 34912 58218 34921
rect 58162 34847 58218 34856
rect 57888 34604 57940 34610
rect 57888 34546 57940 34552
rect 57900 34377 57928 34546
rect 57886 34368 57942 34377
rect 57886 34303 57942 34312
rect 58162 33280 58218 33289
rect 58162 33215 58218 33224
rect 58176 32978 58204 33215
rect 58164 32972 58216 32978
rect 58164 32914 58216 32920
rect 58268 31958 58296 59978
rect 59004 59430 59032 63200
rect 58992 59424 59044 59430
rect 58992 59366 59044 59372
rect 58346 56128 58402 56137
rect 58346 56063 58402 56072
rect 58360 55962 58388 56063
rect 58348 55956 58400 55962
rect 58348 55898 58400 55904
rect 58348 54664 58400 54670
rect 58348 54606 58400 54612
rect 58360 54505 58388 54606
rect 58346 54496 58402 54505
rect 58346 54431 58402 54440
rect 58348 52896 58400 52902
rect 58346 52864 58348 52873
rect 58400 52864 58402 52873
rect 58346 52799 58402 52808
rect 58348 51400 58400 51406
rect 58348 51342 58400 51348
rect 58360 51241 58388 51342
rect 58346 51232 58402 51241
rect 58346 51167 58402 51176
rect 59084 49156 59136 49162
rect 59084 49098 59136 49104
rect 58808 47456 58860 47462
rect 58808 47398 58860 47404
rect 58624 45280 58676 45286
rect 58624 45222 58676 45228
rect 58348 42628 58400 42634
rect 58348 42570 58400 42576
rect 58256 31952 58308 31958
rect 58256 31894 58308 31900
rect 58164 31816 58216 31822
rect 58164 31758 58216 31764
rect 58176 31657 58204 31758
rect 58162 31648 58218 31657
rect 58162 31583 58218 31592
rect 58072 31340 58124 31346
rect 58072 31282 58124 31288
rect 58084 31113 58112 31282
rect 58070 31104 58126 31113
rect 58070 31039 58126 31048
rect 58162 30016 58218 30025
rect 58162 29951 58218 29960
rect 58176 29714 58204 29951
rect 58164 29708 58216 29714
rect 58164 29650 58216 29656
rect 58164 28484 58216 28490
rect 58164 28426 58216 28432
rect 58176 28393 58204 28426
rect 58162 28384 58218 28393
rect 58162 28319 58218 28328
rect 57978 27840 58034 27849
rect 57978 27775 58034 27784
rect 57992 27470 58020 27775
rect 57980 27464 58032 27470
rect 57980 27406 58032 27412
rect 58072 27328 58124 27334
rect 58072 27270 58124 27276
rect 58084 26738 58112 27270
rect 57992 26710 58112 26738
rect 58162 26752 58218 26761
rect 57888 26376 57940 26382
rect 57888 26318 57940 26324
rect 57716 21950 57836 21978
rect 57612 18080 57664 18086
rect 57612 18022 57664 18028
rect 57716 15094 57744 21950
rect 57900 20602 57928 26318
rect 57992 25786 58020 26710
rect 58162 26687 58218 26696
rect 58176 26450 58204 26687
rect 58164 26444 58216 26450
rect 58164 26386 58216 26392
rect 58070 26208 58126 26217
rect 58070 26143 58126 26152
rect 58084 25906 58112 26143
rect 58072 25900 58124 25906
rect 58072 25842 58124 25848
rect 57992 25758 58112 25786
rect 57980 25696 58032 25702
rect 57980 25638 58032 25644
rect 57992 21690 58020 25638
rect 58084 24970 58112 25758
rect 58164 25220 58216 25226
rect 58164 25162 58216 25168
rect 58176 25129 58204 25162
rect 58162 25120 58218 25129
rect 58162 25055 58218 25064
rect 58084 24942 58204 24970
rect 58072 24812 58124 24818
rect 58072 24754 58124 24760
rect 58084 24585 58112 24754
rect 58070 24576 58126 24585
rect 58070 24511 58126 24520
rect 58176 23610 58204 24942
rect 58256 24608 58308 24614
rect 58256 24550 58308 24556
rect 58084 23582 58204 23610
rect 58084 21706 58112 23582
rect 58162 23488 58218 23497
rect 58162 23423 58218 23432
rect 58176 23186 58204 23423
rect 58164 23180 58216 23186
rect 58164 23122 58216 23128
rect 58162 22944 58218 22953
rect 58162 22879 58218 22888
rect 58176 22710 58204 22879
rect 58164 22704 58216 22710
rect 58164 22646 58216 22652
rect 58164 21956 58216 21962
rect 58164 21898 58216 21904
rect 58176 21865 58204 21898
rect 58162 21856 58218 21865
rect 58162 21791 58218 21800
rect 57980 21684 58032 21690
rect 58084 21678 58204 21706
rect 57980 21626 58032 21632
rect 58072 21548 58124 21554
rect 58072 21490 58124 21496
rect 58084 21321 58112 21490
rect 58176 21418 58204 21678
rect 58268 21622 58296 24550
rect 58256 21616 58308 21622
rect 58256 21558 58308 21564
rect 58164 21412 58216 21418
rect 58164 21354 58216 21360
rect 58256 21344 58308 21350
rect 58070 21312 58126 21321
rect 58256 21286 58308 21292
rect 58070 21247 58126 21256
rect 58268 21146 58296 21286
rect 58256 21140 58308 21146
rect 58256 21082 58308 21088
rect 58164 20868 58216 20874
rect 58164 20810 58216 20816
rect 57888 20596 57940 20602
rect 57888 20538 57940 20544
rect 58176 20233 58204 20810
rect 58162 20224 58218 20233
rect 58162 20159 58218 20168
rect 57978 19680 58034 19689
rect 57978 19615 58034 19624
rect 57992 18766 58020 19615
rect 58072 19168 58124 19174
rect 58072 19110 58124 19116
rect 58084 18970 58112 19110
rect 58072 18964 58124 18970
rect 58072 18906 58124 18912
rect 57980 18760 58032 18766
rect 57980 18702 58032 18708
rect 57978 18048 58034 18057
rect 57978 17983 58034 17992
rect 57992 16590 58020 17983
rect 58360 17542 58388 42570
rect 58440 41540 58492 41546
rect 58440 41482 58492 41488
rect 58452 18834 58480 41482
rect 58532 37664 58584 37670
rect 58532 37606 58584 37612
rect 58440 18828 58492 18834
rect 58440 18770 58492 18776
rect 58348 17536 58400 17542
rect 58348 17478 58400 17484
rect 58544 16726 58572 37606
rect 58532 16720 58584 16726
rect 58532 16662 58584 16668
rect 57980 16584 58032 16590
rect 57980 16526 58032 16532
rect 58072 16448 58124 16454
rect 58072 16390 58124 16396
rect 57704 15088 57756 15094
rect 57704 15030 57756 15036
rect 57978 14784 58034 14793
rect 57978 14719 58034 14728
rect 57992 14414 58020 14719
rect 57980 14408 58032 14414
rect 57980 14350 58032 14356
rect 58084 13841 58112 16390
rect 58636 15910 58664 45222
rect 58716 44804 58768 44810
rect 58716 44746 58768 44752
rect 58624 15904 58676 15910
rect 58624 15846 58676 15852
rect 58164 15428 58216 15434
rect 58164 15370 58216 15376
rect 58176 15337 58204 15370
rect 58162 15328 58218 15337
rect 58162 15263 58218 15272
rect 58070 13832 58126 13841
rect 58070 13767 58126 13776
rect 58162 13696 58218 13705
rect 58162 13631 58218 13640
rect 58176 13394 58204 13631
rect 58164 13388 58216 13394
rect 58164 13330 58216 13336
rect 57888 13320 57940 13326
rect 57888 13262 57940 13268
rect 57900 12986 57928 13262
rect 57888 12980 57940 12986
rect 57888 12922 57940 12928
rect 57888 12232 57940 12238
rect 57888 12174 57940 12180
rect 57428 11620 57480 11626
rect 57428 11562 57480 11568
rect 57150 11520 57206 11529
rect 57150 11455 57206 11464
rect 57900 11286 57928 12174
rect 58164 12164 58216 12170
rect 58164 12106 58216 12112
rect 58176 12073 58204 12106
rect 58162 12064 58218 12073
rect 58162 11999 58218 12008
rect 57888 11280 57940 11286
rect 57888 11222 57940 11228
rect 57900 10674 57928 11222
rect 57060 10668 57112 10674
rect 57060 10610 57112 10616
rect 57888 10668 57940 10674
rect 57888 10610 57940 10616
rect 57072 10282 57100 10610
rect 58162 10432 58218 10441
rect 58162 10367 58218 10376
rect 56980 10254 57100 10282
rect 56980 9586 57008 10254
rect 58176 10130 58204 10367
rect 58164 10124 58216 10130
rect 58164 10066 58216 10072
rect 57060 9988 57112 9994
rect 57060 9930 57112 9936
rect 57072 9897 57100 9930
rect 57152 9920 57204 9926
rect 57058 9888 57114 9897
rect 57152 9862 57204 9868
rect 57058 9823 57114 9832
rect 56968 9580 57020 9586
rect 56968 9522 57020 9528
rect 57060 9580 57112 9586
rect 57060 9522 57112 9528
rect 56876 9036 56928 9042
rect 56876 8978 56928 8984
rect 56508 8356 56560 8362
rect 56508 8298 56560 8304
rect 56230 8256 56286 8265
rect 56230 8191 56286 8200
rect 56888 7954 56916 8978
rect 56980 8294 57008 9522
rect 57072 8838 57100 9522
rect 57060 8832 57112 8838
rect 57060 8774 57112 8780
rect 57072 8498 57100 8774
rect 57060 8492 57112 8498
rect 57060 8434 57112 8440
rect 56968 8288 57020 8294
rect 56968 8230 57020 8236
rect 56876 7948 56928 7954
rect 56876 7890 56928 7896
rect 56140 7812 56192 7818
rect 56140 7754 56192 7760
rect 55956 7404 56008 7410
rect 55956 7346 56008 7352
rect 56152 7342 56180 7754
rect 56508 7540 56560 7546
rect 56508 7482 56560 7488
rect 56520 7410 56548 7482
rect 56508 7404 56560 7410
rect 56508 7346 56560 7352
rect 56140 7336 56192 7342
rect 56140 7278 56192 7284
rect 55864 5704 55916 5710
rect 55864 5646 55916 5652
rect 56520 4826 56548 7346
rect 56888 6798 56916 7890
rect 56980 7410 57008 8230
rect 56968 7404 57020 7410
rect 56968 7346 57020 7352
rect 56968 7200 57020 7206
rect 56968 7142 57020 7148
rect 56980 6798 57008 7142
rect 57164 6914 57192 9862
rect 57334 8800 57390 8809
rect 57334 8735 57390 8744
rect 57348 8566 57376 8735
rect 57336 8560 57388 8566
rect 57336 8502 57388 8508
rect 57796 8084 57848 8090
rect 57796 8026 57848 8032
rect 57072 6886 57192 6914
rect 56876 6792 56928 6798
rect 56876 6734 56928 6740
rect 56968 6792 57020 6798
rect 56968 6734 57020 6740
rect 56508 4820 56560 4826
rect 56508 4762 56560 4768
rect 56888 3602 56916 6734
rect 57072 6225 57100 6886
rect 57150 6624 57206 6633
rect 57150 6559 57206 6568
rect 57164 6390 57192 6559
rect 57152 6384 57204 6390
rect 57152 6326 57204 6332
rect 57058 6216 57114 6225
rect 57058 6151 57114 6160
rect 57808 5710 57836 8026
rect 58256 7404 58308 7410
rect 58256 7346 58308 7352
rect 58162 7168 58218 7177
rect 58162 7103 58218 7112
rect 57980 6656 58032 6662
rect 57980 6598 58032 6604
rect 57992 5778 58020 6598
rect 58176 5778 58204 7103
rect 58268 6662 58296 7346
rect 58348 6996 58400 7002
rect 58348 6938 58400 6944
rect 58256 6656 58308 6662
rect 58256 6598 58308 6604
rect 57980 5772 58032 5778
rect 57980 5714 58032 5720
rect 58164 5772 58216 5778
rect 58164 5714 58216 5720
rect 57796 5704 57848 5710
rect 57796 5646 57848 5652
rect 57244 5636 57296 5642
rect 57244 5578 57296 5584
rect 57256 5545 57284 5578
rect 57242 5536 57298 5545
rect 57242 5471 57298 5480
rect 58072 5228 58124 5234
rect 58072 5170 58124 5176
rect 58084 5001 58112 5170
rect 58070 4992 58126 5001
rect 58070 4927 58126 4936
rect 57796 4616 57848 4622
rect 57796 4558 57848 4564
rect 56876 3596 56928 3602
rect 56876 3538 56928 3544
rect 57244 3392 57296 3398
rect 57244 3334 57296 3340
rect 55220 3188 55272 3194
rect 55220 3130 55272 3136
rect 54944 3120 54996 3126
rect 54944 3062 54996 3068
rect 55312 3052 55364 3058
rect 55312 2994 55364 3000
rect 55036 2440 55088 2446
rect 55036 2382 55088 2388
rect 55048 800 55076 2382
rect 55324 800 55352 2994
rect 57256 2446 57284 3334
rect 57244 2440 57296 2446
rect 57244 2382 57296 2388
rect 57336 2372 57388 2378
rect 57336 2314 57388 2320
rect 57348 2281 57376 2314
rect 57334 2272 57390 2281
rect 57334 2207 57390 2216
rect 57808 1737 57836 4558
rect 57888 4208 57940 4214
rect 57888 4150 57940 4156
rect 57900 3913 57928 4150
rect 58360 4146 58388 6938
rect 58728 6730 58756 44746
rect 58820 15638 58848 47398
rect 58900 36100 58952 36106
rect 58900 36042 58952 36048
rect 58912 17678 58940 36042
rect 58992 34740 59044 34746
rect 58992 34682 59044 34688
rect 59004 21894 59032 34682
rect 58992 21888 59044 21894
rect 58992 21830 59044 21836
rect 58900 17672 58952 17678
rect 58900 17614 58952 17620
rect 58808 15632 58860 15638
rect 58808 15574 58860 15580
rect 59096 11898 59124 49098
rect 59176 31136 59228 31142
rect 59176 31078 59228 31084
rect 59188 19514 59216 31078
rect 59176 19508 59228 19514
rect 59176 19450 59228 19456
rect 59084 11892 59136 11898
rect 59084 11834 59136 11840
rect 58716 6724 58768 6730
rect 58716 6666 58768 6672
rect 58348 4140 58400 4146
rect 58348 4082 58400 4088
rect 57886 3904 57942 3913
rect 57886 3839 57942 3848
rect 58162 3360 58218 3369
rect 58162 3295 58218 3304
rect 58176 3126 58204 3295
rect 58164 3120 58216 3126
rect 58164 3062 58216 3068
rect 58256 3052 58308 3058
rect 58256 2994 58308 3000
rect 58162 2816 58218 2825
rect 58162 2751 58218 2760
rect 58176 2446 58204 2751
rect 58268 2650 58296 2994
rect 58256 2644 58308 2650
rect 58256 2586 58308 2592
rect 58164 2440 58216 2446
rect 58164 2382 58216 2388
rect 57794 1728 57850 1737
rect 57794 1663 57850 1672
rect 55956 1352 56008 1358
rect 55956 1294 56008 1300
rect 55968 1193 55996 1294
rect 55954 1184 56010 1193
rect 55954 1119 56010 1128
rect 4526 0 4582 800
rect 4802 0 4858 800
rect 5078 0 5134 800
rect 5354 0 5410 800
rect 5630 0 5686 800
rect 5906 0 5962 800
rect 6182 0 6238 800
rect 6458 0 6514 800
rect 6734 0 6790 800
rect 7010 0 7066 800
rect 7286 0 7342 800
rect 7562 0 7618 800
rect 7838 0 7894 800
rect 8114 0 8170 800
rect 8390 0 8446 800
rect 8666 0 8722 800
rect 8942 0 8998 800
rect 9218 0 9274 800
rect 9494 0 9550 800
rect 9770 0 9826 800
rect 10046 0 10102 800
rect 10322 0 10378 800
rect 10598 0 10654 800
rect 10874 0 10930 800
rect 11150 0 11206 800
rect 11426 0 11482 800
rect 11702 0 11758 800
rect 11978 0 12034 800
rect 12254 0 12310 800
rect 12530 0 12586 800
rect 12806 0 12862 800
rect 13082 0 13138 800
rect 13358 0 13414 800
rect 13634 0 13690 800
rect 13910 0 13966 800
rect 14186 0 14242 800
rect 14462 0 14518 800
rect 14738 0 14794 800
rect 15014 0 15070 800
rect 15290 0 15346 800
rect 15566 0 15622 800
rect 15842 0 15898 800
rect 16118 0 16174 800
rect 16394 0 16450 800
rect 16670 0 16726 800
rect 16946 0 17002 800
rect 17222 0 17278 800
rect 17498 0 17554 800
rect 17774 0 17830 800
rect 18050 0 18106 800
rect 18326 0 18382 800
rect 18602 0 18658 800
rect 18878 0 18934 800
rect 19154 0 19210 800
rect 19430 0 19486 800
rect 19706 0 19762 800
rect 19982 0 20038 800
rect 20258 0 20314 800
rect 20534 0 20590 800
rect 20810 0 20866 800
rect 21086 0 21142 800
rect 21362 0 21418 800
rect 21638 0 21694 800
rect 21914 0 21970 800
rect 22190 0 22246 800
rect 22466 0 22522 800
rect 22742 0 22798 800
rect 23018 0 23074 800
rect 23294 0 23350 800
rect 23570 0 23626 800
rect 23846 0 23902 800
rect 24122 0 24178 800
rect 24398 0 24454 800
rect 24674 0 24730 800
rect 24950 0 25006 800
rect 25226 0 25282 800
rect 25502 0 25558 800
rect 25778 0 25834 800
rect 26054 0 26110 800
rect 26330 0 26386 800
rect 26606 0 26662 800
rect 26882 0 26938 800
rect 27158 0 27214 800
rect 27434 0 27490 800
rect 27710 0 27766 800
rect 27986 0 28042 800
rect 28262 0 28318 800
rect 28538 0 28594 800
rect 28814 0 28870 800
rect 29090 0 29146 800
rect 29366 0 29422 800
rect 29642 0 29698 800
rect 29918 0 29974 800
rect 30194 0 30250 800
rect 30470 0 30526 800
rect 30746 0 30802 800
rect 31022 0 31078 800
rect 31298 0 31354 800
rect 31574 0 31630 800
rect 31850 0 31906 800
rect 32126 0 32182 800
rect 32402 0 32458 800
rect 32678 0 32734 800
rect 32954 0 33010 800
rect 33230 0 33286 800
rect 33506 0 33562 800
rect 33782 0 33838 800
rect 34058 0 34114 800
rect 34334 0 34390 800
rect 34610 0 34666 800
rect 34886 0 34942 800
rect 35162 0 35218 800
rect 35438 0 35494 800
rect 35714 0 35770 800
rect 35990 0 36046 800
rect 36266 0 36322 800
rect 36542 0 36598 800
rect 36818 0 36874 800
rect 37094 0 37150 800
rect 37370 0 37426 800
rect 37646 0 37702 800
rect 37922 0 37978 800
rect 38198 0 38254 800
rect 38474 0 38530 800
rect 38750 0 38806 800
rect 39026 0 39082 800
rect 39302 0 39358 800
rect 39578 0 39634 800
rect 39854 0 39910 800
rect 40130 0 40186 800
rect 40406 0 40462 800
rect 40682 0 40738 800
rect 40958 0 41014 800
rect 41234 0 41290 800
rect 41510 0 41566 800
rect 41786 0 41842 800
rect 42062 0 42118 800
rect 42338 0 42394 800
rect 42614 0 42670 800
rect 42890 0 42946 800
rect 43166 0 43222 800
rect 43442 0 43498 800
rect 43718 0 43774 800
rect 43994 0 44050 800
rect 44270 0 44326 800
rect 44546 0 44602 800
rect 44822 0 44878 800
rect 45098 0 45154 800
rect 45374 0 45430 800
rect 45650 0 45706 800
rect 45926 0 45982 800
rect 46202 0 46258 800
rect 46478 0 46534 800
rect 46754 0 46810 800
rect 47030 0 47086 800
rect 47306 0 47362 800
rect 47582 0 47638 800
rect 47858 0 47914 800
rect 48134 0 48190 800
rect 48410 0 48466 800
rect 48686 0 48742 800
rect 48962 0 49018 800
rect 49238 0 49294 800
rect 49514 0 49570 800
rect 49790 0 49846 800
rect 50066 0 50122 800
rect 50342 0 50398 800
rect 50618 0 50674 800
rect 50894 0 50950 800
rect 51170 0 51226 800
rect 51446 0 51502 800
rect 51722 0 51778 800
rect 51998 0 52054 800
rect 52274 0 52330 800
rect 52550 0 52606 800
rect 52826 0 52882 800
rect 53102 0 53158 800
rect 53378 0 53434 800
rect 53654 0 53710 800
rect 53930 0 53986 800
rect 54206 0 54262 800
rect 54482 0 54538 800
rect 54758 0 54814 800
rect 55034 0 55090 800
rect 55310 0 55366 800
<< via2 >>
rect 1674 61784 1730 61840
rect 1582 60424 1638 60480
rect 1674 59744 1730 59800
rect 2778 61140 2780 61160
rect 2780 61140 2832 61160
rect 2832 61140 2834 61160
rect 2778 61104 2834 61140
rect 4220 61498 4276 61500
rect 4300 61498 4356 61500
rect 4380 61498 4436 61500
rect 4460 61498 4516 61500
rect 4220 61446 4266 61498
rect 4266 61446 4276 61498
rect 4300 61446 4330 61498
rect 4330 61446 4342 61498
rect 4342 61446 4356 61498
rect 4380 61446 4394 61498
rect 4394 61446 4406 61498
rect 4406 61446 4436 61498
rect 4460 61446 4470 61498
rect 4470 61446 4516 61498
rect 4220 61444 4276 61446
rect 4300 61444 4356 61446
rect 4380 61444 4436 61446
rect 4460 61444 4516 61446
rect 4220 60410 4276 60412
rect 4300 60410 4356 60412
rect 4380 60410 4436 60412
rect 4460 60410 4516 60412
rect 4220 60358 4266 60410
rect 4266 60358 4276 60410
rect 4300 60358 4330 60410
rect 4330 60358 4342 60410
rect 4342 60358 4356 60410
rect 4380 60358 4394 60410
rect 4394 60358 4406 60410
rect 4406 60358 4436 60410
rect 4460 60358 4470 60410
rect 4470 60358 4516 60410
rect 4220 60356 4276 60358
rect 4300 60356 4356 60358
rect 4380 60356 4436 60358
rect 4460 60356 4516 60358
rect 1674 59064 1730 59120
rect 1582 58384 1638 58440
rect 1582 57704 1638 57760
rect 1582 57024 1638 57080
rect 1674 56344 1730 56400
rect 1674 55684 1730 55720
rect 1674 55664 1676 55684
rect 1676 55664 1728 55684
rect 1728 55664 1730 55684
rect 1582 54984 1638 55040
rect 1674 54304 1730 54360
rect 1582 53624 1638 53680
rect 1674 52944 1730 53000
rect 1582 52264 1638 52320
rect 1674 51584 1730 51640
rect 1674 50904 1730 50960
rect 1674 50244 1730 50280
rect 1674 50224 1676 50244
rect 1676 50224 1728 50244
rect 1728 50224 1730 50244
rect 1582 49544 1638 49600
rect 1582 48864 1638 48920
rect 1674 48184 1730 48240
rect 1674 47504 1730 47560
rect 1582 46824 1638 46880
rect 1582 46144 1638 46200
rect 1674 45464 1730 45520
rect 1582 44820 1584 44840
rect 1584 44820 1636 44840
rect 1636 44820 1638 44840
rect 1582 44784 1638 44820
rect 1674 44104 1730 44160
rect 1674 43424 1730 43480
rect 1582 42744 1638 42800
rect 1582 42064 1638 42120
rect 1674 41384 1730 41440
rect 1674 40704 1730 40760
rect 1674 40024 1730 40080
rect 1674 39364 1730 39400
rect 1674 39344 1676 39364
rect 1676 39344 1728 39364
rect 1728 39344 1730 39364
rect 1674 38664 1730 38720
rect 1674 37984 1730 38040
rect 1674 37304 1730 37360
rect 1582 36624 1638 36680
rect 1674 35944 1730 36000
rect 1674 35264 1730 35320
rect 1674 34584 1730 34640
rect 1674 33924 1730 33960
rect 1674 33904 1676 33924
rect 1676 33904 1728 33924
rect 1728 33904 1730 33924
rect 1674 33224 1730 33280
rect 1674 32544 1730 32600
rect 1674 31864 1730 31920
rect 1674 31184 1730 31240
rect 1674 30504 1730 30560
rect 1766 29824 1822 29880
rect 1858 29144 1914 29200
rect 1858 28484 1914 28520
rect 1858 28464 1860 28484
rect 1860 28464 1912 28484
rect 1912 28464 1914 28484
rect 1766 27784 1822 27840
rect 1858 27104 1914 27160
rect 1766 26424 1822 26480
rect 1766 25780 1768 25800
rect 1768 25780 1820 25800
rect 1820 25780 1822 25800
rect 1766 25744 1822 25780
rect 1858 25064 1914 25120
rect 1766 24384 1822 24440
rect 1858 23704 1914 23760
rect 1858 23044 1914 23080
rect 1858 23024 1860 23044
rect 1860 23024 1912 23044
rect 1912 23024 1914 23044
rect 1766 22344 1822 22400
rect 1858 21664 1914 21720
rect 1766 20984 1822 21040
rect 1766 20340 1768 20360
rect 1768 20340 1820 20360
rect 1820 20340 1822 20360
rect 1766 20304 1822 20340
rect 1858 19624 1914 19680
rect 1858 18944 1914 19000
rect 1858 18264 1914 18320
rect 1858 17604 1914 17640
rect 1858 17584 1860 17604
rect 1860 17584 1912 17604
rect 1912 17584 1914 17604
rect 1766 16904 1822 16960
rect 1858 16224 1914 16280
rect 1766 15544 1822 15600
rect 1766 14900 1768 14920
rect 1768 14900 1820 14920
rect 1820 14900 1822 14920
rect 1766 14864 1822 14900
rect 1858 14184 1914 14240
rect 1766 13504 1822 13560
rect 1858 12824 1914 12880
rect 1858 12144 1914 12200
rect 1766 11464 1822 11520
rect 1858 10784 1914 10840
rect 1766 10124 1822 10160
rect 1766 10104 1768 10124
rect 1768 10104 1820 10124
rect 1820 10104 1822 10124
rect 1582 9968 1638 10024
rect 4220 59322 4276 59324
rect 4300 59322 4356 59324
rect 4380 59322 4436 59324
rect 4460 59322 4516 59324
rect 4220 59270 4266 59322
rect 4266 59270 4276 59322
rect 4300 59270 4330 59322
rect 4330 59270 4342 59322
rect 4342 59270 4356 59322
rect 4380 59270 4394 59322
rect 4394 59270 4406 59322
rect 4406 59270 4436 59322
rect 4460 59270 4470 59322
rect 4470 59270 4516 59322
rect 4220 59268 4276 59270
rect 4300 59268 4356 59270
rect 4380 59268 4436 59270
rect 4460 59268 4516 59270
rect 4220 58234 4276 58236
rect 4300 58234 4356 58236
rect 4380 58234 4436 58236
rect 4460 58234 4516 58236
rect 4220 58182 4266 58234
rect 4266 58182 4276 58234
rect 4300 58182 4330 58234
rect 4330 58182 4342 58234
rect 4342 58182 4356 58234
rect 4380 58182 4394 58234
rect 4394 58182 4406 58234
rect 4406 58182 4436 58234
rect 4460 58182 4470 58234
rect 4470 58182 4516 58234
rect 4220 58180 4276 58182
rect 4300 58180 4356 58182
rect 4380 58180 4436 58182
rect 4460 58180 4516 58182
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 2410 18808 2466 18864
rect 2410 18692 2466 18728
rect 2410 18672 2412 18692
rect 2412 18672 2464 18692
rect 2464 18672 2466 18692
rect 2410 17196 2466 17232
rect 2410 17176 2412 17196
rect 2412 17176 2464 17196
rect 2464 17176 2466 17196
rect 2410 15988 2412 16008
rect 2412 15988 2464 16008
rect 2464 15988 2466 16008
rect 2410 15952 2466 15988
rect 2410 14476 2466 14512
rect 2410 14456 2412 14476
rect 2412 14456 2464 14476
rect 2464 14456 2466 14476
rect 1766 9460 1768 9480
rect 1768 9460 1820 9480
rect 1820 9460 1822 9480
rect 1766 9424 1822 9460
rect 1858 8744 1914 8800
rect 1766 8064 1822 8120
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 12990 61140 12992 61160
rect 12992 61140 13044 61160
rect 13044 61140 13046 61160
rect 12990 61104 13046 61140
rect 15290 42064 15346 42120
rect 6918 13232 6974 13288
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 6826 10240 6882 10296
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 1858 7384 1914 7440
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 1858 6724 1914 6760
rect 1858 6704 1860 6724
rect 1860 6704 1912 6724
rect 1912 6704 1914 6724
rect 1766 6024 1822 6080
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 1858 5344 1914 5400
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 1766 4664 1822 4720
rect 1766 4020 1768 4040
rect 1768 4020 1820 4040
rect 1820 4020 1822 4040
rect 1766 3984 1822 4020
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 1858 3304 1914 3360
rect 5906 3984 5962 4040
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 1766 2624 1822 2680
rect 1858 1944 1914 2000
rect 6642 2760 6698 2816
rect 7010 3732 7066 3768
rect 7010 3712 7012 3732
rect 7012 3712 7064 3732
rect 7064 3712 7066 3732
rect 8298 8916 8300 8936
rect 8300 8916 8352 8936
rect 8352 8916 8354 8936
rect 8298 8880 8354 8916
rect 7930 7928 7986 7984
rect 9494 10548 9496 10568
rect 9496 10548 9548 10568
rect 9548 10548 9550 10568
rect 9494 10512 9550 10548
rect 7654 3848 7710 3904
rect 11058 21256 11114 21312
rect 9770 7112 9826 7168
rect 8206 2932 8208 2952
rect 8208 2932 8260 2952
rect 8260 2932 8262 2952
rect 8206 2896 8262 2932
rect 8574 3984 8630 4040
rect 9862 4664 9918 4720
rect 9402 3848 9458 3904
rect 8942 2488 8998 2544
rect 9586 3052 9642 3088
rect 9586 3032 9588 3052
rect 9588 3032 9640 3052
rect 9640 3032 9642 3052
rect 11886 12960 11942 13016
rect 12070 12180 12072 12200
rect 12072 12180 12124 12200
rect 12124 12180 12126 12200
rect 12070 12144 12126 12180
rect 11886 11756 11942 11792
rect 11886 11736 11888 11756
rect 11888 11736 11940 11756
rect 11940 11736 11942 11756
rect 10322 2896 10378 2952
rect 12530 7520 12586 7576
rect 12530 3848 12586 3904
rect 12898 8744 12954 8800
rect 12990 3848 13046 3904
rect 12898 3440 12954 3496
rect 14462 5888 14518 5944
rect 15382 16108 15438 16144
rect 15382 16088 15384 16108
rect 15384 16088 15436 16108
rect 15436 16088 15438 16108
rect 15106 13368 15162 13424
rect 14738 11600 14794 11656
rect 14830 11464 14886 11520
rect 14830 11212 14886 11248
rect 14830 11192 14832 11212
rect 14832 11192 14884 11212
rect 14884 11192 14886 11212
rect 15290 11636 15292 11656
rect 15292 11636 15344 11656
rect 15344 11636 15346 11656
rect 15290 11600 15346 11636
rect 15290 9424 15346 9480
rect 16118 11736 16174 11792
rect 15106 8200 15162 8256
rect 14830 6024 14886 6080
rect 15290 8064 15346 8120
rect 15198 7268 15254 7304
rect 15198 7248 15200 7268
rect 15200 7248 15252 7268
rect 15252 7248 15254 7268
rect 15382 6332 15384 6352
rect 15384 6332 15436 6352
rect 15436 6332 15438 6352
rect 15382 6296 15438 6332
rect 15934 9580 15990 9616
rect 15934 9560 15936 9580
rect 15936 9560 15988 9580
rect 15988 9560 15990 9580
rect 15842 9424 15898 9480
rect 15750 8200 15806 8256
rect 16670 11600 16726 11656
rect 18602 59336 18658 59392
rect 17498 50224 17554 50280
rect 19580 60954 19636 60956
rect 19660 60954 19716 60956
rect 19740 60954 19796 60956
rect 19820 60954 19876 60956
rect 19580 60902 19626 60954
rect 19626 60902 19636 60954
rect 19660 60902 19690 60954
rect 19690 60902 19702 60954
rect 19702 60902 19716 60954
rect 19740 60902 19754 60954
rect 19754 60902 19766 60954
rect 19766 60902 19796 60954
rect 19820 60902 19830 60954
rect 19830 60902 19876 60954
rect 19580 60900 19636 60902
rect 19660 60900 19716 60902
rect 19740 60900 19796 60902
rect 19820 60900 19876 60902
rect 19580 59866 19636 59868
rect 19660 59866 19716 59868
rect 19740 59866 19796 59868
rect 19820 59866 19876 59868
rect 19580 59814 19626 59866
rect 19626 59814 19636 59866
rect 19660 59814 19690 59866
rect 19690 59814 19702 59866
rect 19702 59814 19716 59866
rect 19740 59814 19754 59866
rect 19754 59814 19766 59866
rect 19766 59814 19796 59866
rect 19820 59814 19830 59866
rect 19830 59814 19876 59866
rect 19580 59812 19636 59814
rect 19660 59812 19716 59814
rect 19740 59812 19796 59814
rect 19820 59812 19876 59814
rect 19580 58778 19636 58780
rect 19660 58778 19716 58780
rect 19740 58778 19796 58780
rect 19820 58778 19876 58780
rect 19580 58726 19626 58778
rect 19626 58726 19636 58778
rect 19660 58726 19690 58778
rect 19690 58726 19702 58778
rect 19702 58726 19716 58778
rect 19740 58726 19754 58778
rect 19754 58726 19766 58778
rect 19766 58726 19796 58778
rect 19820 58726 19830 58778
rect 19830 58726 19876 58778
rect 19580 58724 19636 58726
rect 19660 58724 19716 58726
rect 19740 58724 19796 58726
rect 19820 58724 19876 58726
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 22742 60696 22798 60752
rect 20718 37848 20774 37904
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 18510 20460 18566 20496
rect 18510 20440 18512 20460
rect 18512 20440 18564 20460
rect 18564 20440 18566 20460
rect 17038 11736 17094 11792
rect 16302 7792 16358 7848
rect 16854 11056 16910 11112
rect 16118 6296 16174 6352
rect 17406 11464 17462 11520
rect 17038 8608 17094 8664
rect 17958 12960 18014 13016
rect 17866 11212 17922 11248
rect 17866 11192 17868 11212
rect 17868 11192 17920 11212
rect 17920 11192 17922 11212
rect 17774 10376 17830 10432
rect 17682 10240 17738 10296
rect 17498 8472 17554 8528
rect 17222 6976 17278 7032
rect 16946 4800 17002 4856
rect 16762 2896 16818 2952
rect 17774 4936 17830 4992
rect 17958 3848 18014 3904
rect 18694 13776 18750 13832
rect 18418 13404 18420 13424
rect 18420 13404 18472 13424
rect 18472 13404 18474 13424
rect 18418 13368 18474 13404
rect 18510 8336 18566 8392
rect 18602 7384 18658 7440
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19614 14340 19670 14376
rect 19614 14320 19616 14340
rect 19616 14320 19668 14340
rect 19668 14320 19670 14340
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19246 11620 19302 11656
rect 19246 11600 19248 11620
rect 19248 11600 19300 11620
rect 19300 11600 19302 11620
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19522 12552 19578 12608
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19982 11872 20038 11928
rect 20166 12552 20222 12608
rect 22098 60288 22154 60344
rect 22098 60152 22154 60208
rect 22558 60288 22614 60344
rect 21546 34076 21548 34096
rect 21548 34076 21600 34096
rect 21600 34076 21602 34096
rect 21546 34040 21602 34076
rect 21454 33360 21510 33416
rect 22006 59608 22062 59664
rect 20718 25200 20774 25256
rect 22558 37748 22560 37768
rect 22560 37748 22612 37768
rect 22612 37748 22614 37768
rect 22558 37712 22614 37748
rect 20902 18536 20958 18592
rect 21638 18284 21694 18320
rect 21638 18264 21640 18284
rect 21640 18264 21692 18284
rect 21692 18264 21694 18284
rect 20718 15952 20774 16008
rect 20442 15136 20498 15192
rect 19798 11600 19854 11656
rect 19706 11328 19762 11384
rect 20074 11464 20130 11520
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19614 10648 19670 10704
rect 19246 9288 19302 9344
rect 19154 9016 19210 9072
rect 19154 8744 19210 8800
rect 19798 10240 19854 10296
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 18970 7520 19026 7576
rect 19982 8064 20038 8120
rect 19154 7656 19210 7712
rect 19154 7268 19210 7304
rect 19154 7248 19156 7268
rect 19156 7248 19208 7268
rect 19208 7248 19210 7268
rect 19062 7112 19118 7168
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19522 7420 19524 7440
rect 19524 7420 19576 7440
rect 19576 7420 19578 7440
rect 19522 7384 19578 7420
rect 19890 7284 19892 7304
rect 19892 7284 19944 7304
rect 19944 7284 19946 7304
rect 19890 7248 19946 7284
rect 19062 6160 19118 6216
rect 18878 5616 18934 5672
rect 18970 4684 19026 4720
rect 18970 4664 18972 4684
rect 18972 4664 19024 4684
rect 19024 4664 19026 4684
rect 18418 3576 18474 3632
rect 17498 2624 17554 2680
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19522 5752 19578 5808
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19430 5208 19486 5264
rect 19430 4564 19432 4584
rect 19432 4564 19484 4584
rect 19484 4564 19486 4584
rect 19430 4528 19486 4564
rect 19890 4548 19946 4584
rect 19890 4528 19892 4548
rect 19892 4528 19944 4548
rect 19944 4528 19946 4548
rect 19338 4392 19394 4448
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19338 4276 19394 4312
rect 19338 4256 19340 4276
rect 19340 4256 19392 4276
rect 19392 4256 19394 4276
rect 19522 4156 19524 4176
rect 19524 4156 19576 4176
rect 19576 4156 19578 4176
rect 19522 4120 19578 4156
rect 20350 8608 20406 8664
rect 20902 15680 20958 15736
rect 20718 14592 20774 14648
rect 19430 4020 19432 4040
rect 19432 4020 19484 4040
rect 19484 4020 19486 4040
rect 19430 3984 19486 4020
rect 19522 3596 19578 3632
rect 19522 3576 19524 3596
rect 19524 3576 19576 3596
rect 19576 3576 19578 3596
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19890 2624 19946 2680
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 19706 1944 19762 2000
rect 21546 15816 21602 15872
rect 21454 14340 21510 14376
rect 21454 14320 21456 14340
rect 21456 14320 21508 14340
rect 21508 14320 21510 14340
rect 21270 12144 21326 12200
rect 21086 8336 21142 8392
rect 20626 6160 20682 6216
rect 20902 5244 20904 5264
rect 20904 5244 20956 5264
rect 20956 5244 20958 5264
rect 20902 5208 20958 5244
rect 20810 4528 20866 4584
rect 20718 3732 20774 3768
rect 20718 3712 20720 3732
rect 20720 3712 20772 3732
rect 20772 3712 20774 3732
rect 21454 11328 21510 11384
rect 22742 59628 22798 59664
rect 22742 59608 22744 59628
rect 22744 59608 22796 59628
rect 22796 59608 22798 59628
rect 22834 53896 22890 53952
rect 23386 59644 23388 59664
rect 23388 59644 23440 59664
rect 23440 59644 23442 59664
rect 23386 59608 23442 59644
rect 22926 37884 22928 37904
rect 22928 37884 22980 37904
rect 22980 37884 22982 37904
rect 22926 37848 22982 37884
rect 23018 37712 23074 37768
rect 22742 34040 22798 34096
rect 22558 25492 22614 25528
rect 22558 25472 22560 25492
rect 22560 25472 22612 25492
rect 22612 25472 22614 25492
rect 22558 21256 22614 21312
rect 22466 18400 22522 18456
rect 21914 15816 21970 15872
rect 22190 13776 22246 13832
rect 21822 12416 21878 12472
rect 21730 11056 21786 11112
rect 21914 10104 21970 10160
rect 21546 7248 21602 7304
rect 21454 5072 21510 5128
rect 21086 4120 21142 4176
rect 21178 3984 21234 4040
rect 20902 3576 20958 3632
rect 20994 2388 20996 2408
rect 20996 2388 21048 2408
rect 21048 2388 21050 2408
rect 20994 2352 21050 2388
rect 21822 5616 21878 5672
rect 22466 15952 22522 16008
rect 22190 11600 22246 11656
rect 22098 10104 22154 10160
rect 22466 8916 22468 8936
rect 22468 8916 22520 8936
rect 22520 8916 22522 8936
rect 22466 8880 22522 8916
rect 22374 7112 22430 7168
rect 22374 5480 22430 5536
rect 22282 3168 22338 3224
rect 21730 2896 21786 2952
rect 22650 8880 22706 8936
rect 22742 8744 22798 8800
rect 23018 11600 23074 11656
rect 23386 18264 23442 18320
rect 23386 15408 23442 15464
rect 23294 11872 23350 11928
rect 23110 10376 23166 10432
rect 23018 10104 23074 10160
rect 23386 9832 23442 9888
rect 23386 9696 23442 9752
rect 27342 48864 27398 48920
rect 24858 34584 24914 34640
rect 24398 17176 24454 17232
rect 24858 29552 24914 29608
rect 23846 13096 23902 13152
rect 24030 12008 24086 12064
rect 23662 10920 23718 10976
rect 23386 9288 23442 9344
rect 23570 9288 23626 9344
rect 23938 11076 23994 11112
rect 23938 11056 23940 11076
rect 23940 11056 23992 11076
rect 23992 11056 23994 11076
rect 23846 9288 23902 9344
rect 23386 5344 23442 5400
rect 23570 5072 23626 5128
rect 23662 4936 23718 4992
rect 24122 8744 24178 8800
rect 24398 13812 24400 13832
rect 24400 13812 24452 13832
rect 24452 13812 24454 13832
rect 24398 13776 24454 13812
rect 24306 12044 24308 12064
rect 24308 12044 24360 12064
rect 24360 12044 24362 12064
rect 24306 12008 24362 12044
rect 24950 19796 24952 19816
rect 24952 19796 25004 19816
rect 25004 19796 25006 19816
rect 24950 19760 25006 19796
rect 24766 18400 24822 18456
rect 25134 20440 25190 20496
rect 25042 17484 25044 17504
rect 25044 17484 25096 17504
rect 25096 17484 25098 17504
rect 25042 17448 25098 17484
rect 25226 17212 25228 17232
rect 25228 17212 25280 17232
rect 25280 17212 25282 17232
rect 25226 17176 25282 17212
rect 24858 16396 24860 16416
rect 24860 16396 24912 16416
rect 24912 16396 24914 16416
rect 24858 16360 24914 16396
rect 24674 15136 24730 15192
rect 25226 16360 25282 16416
rect 24490 11600 24546 11656
rect 24398 11192 24454 11248
rect 24306 9288 24362 9344
rect 24490 11092 24492 11112
rect 24492 11092 24544 11112
rect 24544 11092 24546 11112
rect 24490 11056 24546 11092
rect 24674 10956 24676 10976
rect 24676 10956 24728 10976
rect 24728 10956 24730 10976
rect 24398 9152 24454 9208
rect 24306 8608 24362 8664
rect 23846 7112 23902 7168
rect 23570 2896 23626 2952
rect 24674 10920 24730 10956
rect 24674 9016 24730 9072
rect 24674 8336 24730 8392
rect 24950 10784 25006 10840
rect 25318 15428 25374 15464
rect 25318 15408 25320 15428
rect 25320 15408 25372 15428
rect 25372 15408 25374 15428
rect 25962 20440 26018 20496
rect 25686 15544 25742 15600
rect 24950 8200 25006 8256
rect 24398 4528 24454 4584
rect 25594 10784 25650 10840
rect 25962 16360 26018 16416
rect 28630 59608 28686 59664
rect 26514 18536 26570 18592
rect 26146 13912 26202 13968
rect 26054 11464 26110 11520
rect 25778 9832 25834 9888
rect 25594 9696 25650 9752
rect 25318 9152 25374 9208
rect 25502 9288 25558 9344
rect 26054 10376 26110 10432
rect 25686 7792 25742 7848
rect 26698 15272 26754 15328
rect 26974 12300 27030 12336
rect 26974 12280 26976 12300
rect 26976 12280 27028 12300
rect 27028 12280 27030 12300
rect 26422 9560 26478 9616
rect 26146 8472 26202 8528
rect 26606 9560 26662 9616
rect 26698 8336 26754 8392
rect 26238 5752 26294 5808
rect 24214 2760 24270 2816
rect 24858 3576 24914 3632
rect 27526 16904 27582 16960
rect 30378 60052 30380 60072
rect 30380 60052 30432 60072
rect 30432 60052 30434 60072
rect 30378 60016 30434 60052
rect 30654 59880 30710 59936
rect 28998 27512 29054 27568
rect 27894 16532 27896 16552
rect 27896 16532 27948 16552
rect 27948 16532 27950 16552
rect 27894 16496 27950 16532
rect 28170 17312 28226 17368
rect 27618 13096 27674 13152
rect 27342 12280 27398 12336
rect 27342 11736 27398 11792
rect 27342 11056 27398 11112
rect 27250 10376 27306 10432
rect 27158 9288 27214 9344
rect 27158 5888 27214 5944
rect 27802 11056 27858 11112
rect 27618 9988 27674 10024
rect 27618 9968 27620 9988
rect 27620 9968 27672 9988
rect 27672 9968 27674 9988
rect 27894 10104 27950 10160
rect 27802 9560 27858 9616
rect 27526 9288 27582 9344
rect 27986 8916 27988 8936
rect 27988 8916 28040 8936
rect 28040 8916 28042 8936
rect 27526 7112 27582 7168
rect 27986 8880 28042 8916
rect 27618 5072 27674 5128
rect 27158 4664 27214 4720
rect 27066 3712 27122 3768
rect 27250 3460 27306 3496
rect 27802 5752 27858 5808
rect 27710 3732 27766 3768
rect 27710 3712 27712 3732
rect 27712 3712 27764 3732
rect 27764 3712 27766 3732
rect 27250 3440 27252 3460
rect 27252 3440 27304 3460
rect 27304 3440 27306 3460
rect 27158 3032 27214 3088
rect 27526 3052 27582 3088
rect 27526 3032 27528 3052
rect 27528 3032 27580 3052
rect 27580 3032 27582 3052
rect 28170 12416 28226 12472
rect 28906 17856 28962 17912
rect 29090 17176 29146 17232
rect 28722 17040 28778 17096
rect 28446 15680 28502 15736
rect 28446 15408 28502 15464
rect 28170 11056 28226 11112
rect 28170 8472 28226 8528
rect 28354 12008 28410 12064
rect 28538 9832 28594 9888
rect 28446 9580 28502 9616
rect 28446 9560 28448 9580
rect 28448 9560 28500 9580
rect 28500 9560 28502 9580
rect 28170 6296 28226 6352
rect 28078 3576 28134 3632
rect 28078 3032 28134 3088
rect 28998 13912 29054 13968
rect 29550 17856 29606 17912
rect 29182 11192 29238 11248
rect 28998 10648 29054 10704
rect 29182 10648 29238 10704
rect 28906 10240 28962 10296
rect 28722 9968 28778 10024
rect 28814 9560 28870 9616
rect 30378 18400 30434 18456
rect 30654 18536 30710 18592
rect 29826 15020 29882 15056
rect 29826 15000 29828 15020
rect 29828 15000 29880 15020
rect 29880 15000 29882 15020
rect 30838 17312 30894 17368
rect 29458 10104 29514 10160
rect 29550 9716 29606 9752
rect 29550 9696 29552 9716
rect 29552 9696 29604 9716
rect 29604 9696 29606 9716
rect 29550 9424 29606 9480
rect 29550 8508 29552 8528
rect 29552 8508 29604 8528
rect 29604 8508 29606 8528
rect 29550 8472 29606 8508
rect 28814 5208 28870 5264
rect 28722 4664 28778 4720
rect 27894 2488 27950 2544
rect 30010 10920 30066 10976
rect 30470 15308 30472 15328
rect 30472 15308 30524 15328
rect 30524 15308 30526 15328
rect 30470 15272 30526 15308
rect 30470 15000 30526 15056
rect 30194 10784 30250 10840
rect 30010 9696 30066 9752
rect 29734 9596 29736 9616
rect 29736 9596 29788 9616
rect 29788 9596 29790 9616
rect 29734 9560 29790 9596
rect 29090 3032 29146 3088
rect 29642 6296 29698 6352
rect 30194 9560 30250 9616
rect 29918 7112 29974 7168
rect 29734 5752 29790 5808
rect 31298 17992 31354 18048
rect 31482 17992 31538 18048
rect 31758 17992 31814 18048
rect 31666 16768 31722 16824
rect 31850 15816 31906 15872
rect 31574 13388 31630 13424
rect 31574 13368 31576 13388
rect 31576 13368 31628 13388
rect 31628 13368 31630 13388
rect 31390 12844 31446 12880
rect 31390 12824 31392 12844
rect 31392 12824 31444 12844
rect 31444 12824 31446 12844
rect 31390 11056 31446 11112
rect 30654 9560 30710 9616
rect 30562 7656 30618 7712
rect 30378 6976 30434 7032
rect 30194 5208 30250 5264
rect 30378 3848 30434 3904
rect 30930 8200 30986 8256
rect 32034 14320 32090 14376
rect 31758 11192 31814 11248
rect 31758 10648 31814 10704
rect 31574 10376 31630 10432
rect 32126 13252 32182 13288
rect 32126 13232 32128 13252
rect 32128 13232 32180 13252
rect 32180 13232 32182 13252
rect 32678 59880 32734 59936
rect 32770 43152 32826 43208
rect 32402 17740 32458 17776
rect 32402 17720 32404 17740
rect 32404 17720 32456 17740
rect 32456 17720 32458 17740
rect 32586 17584 32642 17640
rect 32402 15952 32458 16008
rect 32310 12008 32366 12064
rect 32586 15816 32642 15872
rect 32678 13096 32734 13152
rect 32034 10784 32090 10840
rect 32126 10648 32182 10704
rect 31298 8372 31300 8392
rect 31300 8372 31352 8392
rect 31352 8372 31354 8392
rect 31298 8336 31354 8372
rect 31206 7656 31262 7712
rect 30838 6976 30894 7032
rect 30838 5344 30894 5400
rect 31850 9152 31906 9208
rect 31574 8744 31630 8800
rect 31666 8608 31722 8664
rect 31666 8336 31722 8392
rect 31482 7520 31538 7576
rect 31482 6740 31484 6760
rect 31484 6740 31536 6760
rect 31536 6740 31538 6760
rect 31482 6704 31538 6740
rect 31298 5228 31354 5264
rect 31298 5208 31300 5228
rect 31300 5208 31352 5228
rect 31352 5208 31354 5228
rect 31942 4684 31998 4720
rect 32218 9968 32274 10024
rect 32862 14456 32918 14512
rect 34940 61498 34996 61500
rect 35020 61498 35076 61500
rect 35100 61498 35156 61500
rect 35180 61498 35236 61500
rect 34940 61446 34986 61498
rect 34986 61446 34996 61498
rect 35020 61446 35050 61498
rect 35050 61446 35062 61498
rect 35062 61446 35076 61498
rect 35100 61446 35114 61498
rect 35114 61446 35126 61498
rect 35126 61446 35156 61498
rect 35180 61446 35190 61498
rect 35190 61446 35236 61498
rect 34940 61444 34996 61446
rect 35020 61444 35076 61446
rect 35100 61444 35156 61446
rect 35180 61444 35236 61446
rect 34940 60410 34996 60412
rect 35020 60410 35076 60412
rect 35100 60410 35156 60412
rect 35180 60410 35236 60412
rect 34940 60358 34986 60410
rect 34986 60358 34996 60410
rect 35020 60358 35050 60410
rect 35050 60358 35062 60410
rect 35062 60358 35076 60410
rect 35100 60358 35114 60410
rect 35114 60358 35126 60410
rect 35126 60358 35156 60410
rect 35180 60358 35190 60410
rect 35190 60358 35236 60410
rect 34940 60356 34996 60358
rect 35020 60356 35076 60358
rect 35100 60356 35156 60358
rect 35180 60356 35236 60358
rect 34940 59322 34996 59324
rect 35020 59322 35076 59324
rect 35100 59322 35156 59324
rect 35180 59322 35236 59324
rect 34940 59270 34986 59322
rect 34986 59270 34996 59322
rect 35020 59270 35050 59322
rect 35050 59270 35062 59322
rect 35062 59270 35076 59322
rect 35100 59270 35114 59322
rect 35114 59270 35126 59322
rect 35126 59270 35156 59322
rect 35180 59270 35190 59322
rect 35190 59270 35236 59322
rect 34940 59268 34996 59270
rect 35020 59268 35076 59270
rect 35100 59268 35156 59270
rect 35180 59268 35236 59270
rect 34940 58234 34996 58236
rect 35020 58234 35076 58236
rect 35100 58234 35156 58236
rect 35180 58234 35236 58236
rect 34940 58182 34986 58234
rect 34986 58182 34996 58234
rect 35020 58182 35050 58234
rect 35050 58182 35062 58234
rect 35062 58182 35076 58234
rect 35100 58182 35114 58234
rect 35114 58182 35126 58234
rect 35126 58182 35156 58234
rect 35180 58182 35190 58234
rect 35190 58182 35236 58234
rect 34940 58180 34996 58182
rect 35020 58180 35076 58182
rect 35100 58180 35156 58182
rect 35180 58180 35236 58182
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 33138 18400 33194 18456
rect 33046 17176 33102 17232
rect 33782 17856 33838 17912
rect 33598 16788 33654 16824
rect 33598 16768 33600 16788
rect 33600 16768 33652 16788
rect 33652 16768 33654 16788
rect 32310 9016 32366 9072
rect 32218 5616 32274 5672
rect 31942 4664 31944 4684
rect 31944 4664 31996 4684
rect 31996 4664 31998 4684
rect 31482 4528 31538 4584
rect 32218 4428 32220 4448
rect 32220 4428 32272 4448
rect 32272 4428 32274 4448
rect 32218 4392 32274 4428
rect 32494 8200 32550 8256
rect 32770 8492 32826 8528
rect 32770 8472 32772 8492
rect 32772 8472 32824 8492
rect 32824 8472 32826 8492
rect 32586 6296 32642 6352
rect 33414 10648 33470 10704
rect 33230 9152 33286 9208
rect 33414 9580 33470 9616
rect 33414 9560 33416 9580
rect 33416 9560 33468 9580
rect 33468 9560 33470 9580
rect 32954 8744 33010 8800
rect 32862 5888 32918 5944
rect 32586 5616 32642 5672
rect 32586 5344 32642 5400
rect 32770 4020 32772 4040
rect 32772 4020 32824 4040
rect 32824 4020 32826 4040
rect 32770 3984 32826 4020
rect 32770 2896 32826 2952
rect 33138 4392 33194 4448
rect 33690 7112 33746 7168
rect 34518 17312 34574 17368
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 35070 19896 35126 19952
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 35162 17584 35218 17640
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34242 12688 34298 12744
rect 33874 8492 33930 8528
rect 33874 8472 33876 8492
rect 33876 8472 33928 8492
rect 33928 8472 33930 8492
rect 34426 10376 34482 10432
rect 34334 8880 34390 8936
rect 33506 5480 33562 5536
rect 33414 4800 33470 4856
rect 35254 14320 35310 14376
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 35346 12180 35348 12200
rect 35348 12180 35400 12200
rect 35400 12180 35402 12200
rect 35346 12144 35402 12180
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 35254 10784 35310 10840
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34150 5344 34206 5400
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 35530 10104 35586 10160
rect 35530 9288 35586 9344
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 35438 7540 35494 7576
rect 35438 7520 35440 7540
rect 35440 7520 35492 7540
rect 35492 7520 35494 7540
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34610 4664 34666 4720
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 36542 17448 36598 17504
rect 36266 13268 36268 13288
rect 36268 13268 36320 13288
rect 36320 13268 36322 13288
rect 36266 13232 36322 13268
rect 36450 12844 36506 12880
rect 36450 12824 36452 12844
rect 36452 12824 36504 12844
rect 36504 12824 36506 12844
rect 35806 12008 35862 12064
rect 36082 12144 36138 12200
rect 36082 10648 36138 10704
rect 36174 9968 36230 10024
rect 35806 6724 35862 6760
rect 35806 6704 35808 6724
rect 35808 6704 35860 6724
rect 35860 6704 35862 6724
rect 35990 3984 36046 4040
rect 37278 42644 37280 42664
rect 37280 42644 37332 42664
rect 37332 42644 37334 42664
rect 37278 42608 37334 42644
rect 37002 18536 37058 18592
rect 36726 11872 36782 11928
rect 36542 10512 36598 10568
rect 36450 9052 36452 9072
rect 36452 9052 36504 9072
rect 36504 9052 36506 9072
rect 36450 9016 36506 9052
rect 36634 8744 36690 8800
rect 36542 7928 36598 7984
rect 36358 5344 36414 5400
rect 36266 3984 36322 4040
rect 36358 3304 36414 3360
rect 36542 2896 36598 2952
rect 37278 13232 37334 13288
rect 37462 13096 37518 13152
rect 37094 8916 37096 8936
rect 37096 8916 37148 8936
rect 37148 8916 37150 8936
rect 37094 8880 37150 8916
rect 37462 8608 37518 8664
rect 38014 45328 38070 45384
rect 38290 17040 38346 17096
rect 38566 17448 38622 17504
rect 38658 17312 38714 17368
rect 38750 17176 38806 17232
rect 38474 17060 38530 17096
rect 38474 17040 38476 17060
rect 38476 17040 38528 17060
rect 38528 17040 38530 17060
rect 38382 16904 38438 16960
rect 38842 16904 38898 16960
rect 38842 16224 38898 16280
rect 38566 13368 38622 13424
rect 38106 12008 38162 12064
rect 37830 11056 37886 11112
rect 37462 8336 37518 8392
rect 38750 10260 38806 10296
rect 38750 10240 38752 10260
rect 38752 10240 38804 10260
rect 38804 10240 38806 10260
rect 38658 10140 38666 10160
rect 38666 10140 38714 10160
rect 38658 10104 38714 10140
rect 39026 12688 39082 12744
rect 38842 9968 38898 10024
rect 38382 9152 38438 9208
rect 38658 9832 38714 9888
rect 38750 9696 38806 9752
rect 38750 9560 38806 9616
rect 38566 9036 38622 9072
rect 38566 9016 38568 9036
rect 38568 9016 38620 9036
rect 38620 9016 38622 9036
rect 38290 8608 38346 8664
rect 37370 3848 37426 3904
rect 37370 3032 37426 3088
rect 37278 2896 37334 2952
rect 38106 6160 38162 6216
rect 38474 8472 38530 8528
rect 38658 8064 38714 8120
rect 38658 7948 38714 7984
rect 38658 7928 38660 7948
rect 38660 7928 38712 7948
rect 38712 7928 38714 7948
rect 38382 6432 38438 6488
rect 38290 3032 38346 3088
rect 39210 12552 39266 12608
rect 39118 9696 39174 9752
rect 39394 8880 39450 8936
rect 38566 3340 38568 3360
rect 38568 3340 38620 3360
rect 38620 3340 38622 3360
rect 38566 3304 38622 3340
rect 39210 7928 39266 7984
rect 39670 17484 39672 17504
rect 39672 17484 39724 17504
rect 39724 17484 39726 17504
rect 39670 17448 39726 17484
rect 39762 17060 39818 17096
rect 39762 17040 39764 17060
rect 39764 17040 39816 17060
rect 39816 17040 39818 17060
rect 39578 6840 39634 6896
rect 40038 18828 40094 18864
rect 40038 18808 40040 18828
rect 40040 18808 40092 18828
rect 40092 18808 40094 18828
rect 40038 15544 40094 15600
rect 40130 11736 40186 11792
rect 40038 11328 40094 11384
rect 40222 8916 40224 8936
rect 40224 8916 40276 8936
rect 40276 8916 40278 8936
rect 40222 8880 40278 8916
rect 39946 3848 40002 3904
rect 40130 3984 40186 4040
rect 41970 59336 42026 59392
rect 41142 18808 41198 18864
rect 40958 18572 40960 18592
rect 40960 18572 41012 18592
rect 41012 18572 41014 18592
rect 40958 18536 41014 18572
rect 40958 15852 40960 15872
rect 40960 15852 41012 15872
rect 41012 15852 41014 15872
rect 40958 15816 41014 15852
rect 41050 15544 41106 15600
rect 41326 17212 41328 17232
rect 41328 17212 41380 17232
rect 41380 17212 41382 17232
rect 41326 17176 41382 17212
rect 41878 19116 41880 19136
rect 41880 19116 41932 19136
rect 41932 19116 41934 19136
rect 41878 19080 41934 19116
rect 41418 11192 41474 11248
rect 40682 5072 40738 5128
rect 41694 11736 41750 11792
rect 42246 19236 42302 19272
rect 42246 19216 42248 19236
rect 42248 19216 42300 19236
rect 42300 19216 42302 19236
rect 42154 12416 42210 12472
rect 42706 57296 42762 57352
rect 42798 18300 42800 18320
rect 42800 18300 42852 18320
rect 42852 18300 42854 18320
rect 42798 18264 42854 18300
rect 42890 16496 42946 16552
rect 42522 14456 42578 14512
rect 41878 9288 41934 9344
rect 41970 5752 42026 5808
rect 42430 11328 42486 11384
rect 42890 10104 42946 10160
rect 43626 19080 43682 19136
rect 42614 3984 42670 4040
rect 42706 3848 42762 3904
rect 42614 2624 42670 2680
rect 43350 4528 43406 4584
rect 43350 3984 43406 4040
rect 50300 60954 50356 60956
rect 50380 60954 50436 60956
rect 50460 60954 50516 60956
rect 50540 60954 50596 60956
rect 50300 60902 50346 60954
rect 50346 60902 50356 60954
rect 50380 60902 50410 60954
rect 50410 60902 50422 60954
rect 50422 60902 50436 60954
rect 50460 60902 50474 60954
rect 50474 60902 50486 60954
rect 50486 60902 50516 60954
rect 50540 60902 50550 60954
rect 50550 60902 50596 60954
rect 50300 60900 50356 60902
rect 50380 60900 50436 60902
rect 50460 60900 50516 60902
rect 50540 60900 50596 60902
rect 53378 61104 53434 61160
rect 50300 59866 50356 59868
rect 50380 59866 50436 59868
rect 50460 59866 50516 59868
rect 50540 59866 50596 59868
rect 50300 59814 50346 59866
rect 50346 59814 50356 59866
rect 50380 59814 50410 59866
rect 50410 59814 50422 59866
rect 50422 59814 50436 59866
rect 50460 59814 50474 59866
rect 50474 59814 50486 59866
rect 50486 59814 50516 59866
rect 50540 59814 50550 59866
rect 50550 59814 50596 59866
rect 50300 59812 50356 59814
rect 50380 59812 50436 59814
rect 50460 59812 50516 59814
rect 50540 59812 50596 59814
rect 50300 58778 50356 58780
rect 50380 58778 50436 58780
rect 50460 58778 50516 58780
rect 50540 58778 50596 58780
rect 50300 58726 50346 58778
rect 50346 58726 50356 58778
rect 50380 58726 50410 58778
rect 50410 58726 50422 58778
rect 50422 58726 50436 58778
rect 50460 58726 50474 58778
rect 50474 58726 50486 58778
rect 50486 58726 50516 58778
rect 50540 58726 50550 58778
rect 50550 58726 50596 58778
rect 50300 58724 50356 58726
rect 50380 58724 50436 58726
rect 50460 58724 50516 58726
rect 50540 58724 50596 58726
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 44546 10240 44602 10296
rect 43994 4564 43996 4584
rect 43996 4564 44048 4584
rect 44048 4564 44050 4584
rect 43994 4528 44050 4564
rect 43442 3712 43498 3768
rect 43350 2624 43406 2680
rect 43626 2624 43682 2680
rect 43810 3596 43866 3632
rect 43810 3576 43812 3596
rect 43812 3576 43864 3596
rect 43864 3576 43866 3596
rect 44178 3576 44234 3632
rect 45006 6296 45062 6352
rect 45006 4120 45062 4176
rect 45190 3984 45246 4040
rect 45466 3848 45522 3904
rect 45374 2644 45430 2680
rect 45374 2624 45376 2644
rect 45376 2624 45428 2644
rect 45428 2624 45430 2644
rect 46386 19236 46442 19272
rect 46386 19216 46388 19236
rect 46388 19216 46440 19236
rect 46440 19216 46442 19236
rect 46018 9152 46074 9208
rect 46570 18536 46626 18592
rect 46570 16088 46626 16144
rect 46938 18300 46940 18320
rect 46940 18300 46992 18320
rect 46992 18300 46994 18320
rect 46938 18264 46994 18300
rect 46938 9424 46994 9480
rect 46846 3712 46902 3768
rect 47490 3576 47546 3632
rect 47858 8064 47914 8120
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 49974 20032 50030 20088
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 50158 19760 50214 19816
rect 50710 19796 50712 19816
rect 50712 19796 50764 19816
rect 50764 19796 50766 19816
rect 50710 19760 50766 19796
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 51630 20032 51686 20088
rect 51170 17196 51226 17232
rect 51170 17176 51172 17196
rect 51172 17176 51224 17196
rect 51224 17176 51226 17196
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 49606 2760 49662 2816
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50526 2796 50528 2816
rect 50528 2796 50580 2816
rect 50580 2796 50582 2816
rect 50526 2760 50582 2796
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 55402 61512 55458 61568
rect 56414 62600 56470 62656
rect 56138 62056 56194 62112
rect 56506 60968 56562 61024
rect 57242 60424 57298 60480
rect 58254 60152 58310 60208
rect 58070 59880 58126 59936
rect 58070 59336 58126 59392
rect 58070 58928 58126 58984
rect 58162 58792 58218 58848
rect 57886 58248 57942 58304
rect 57978 57704 58034 57760
rect 57886 57160 57942 57216
rect 53930 17076 53932 17096
rect 53932 17076 53984 17096
rect 53984 17076 53986 17096
rect 53930 17040 53986 17076
rect 54298 17196 54354 17232
rect 54298 17176 54300 17196
rect 54300 17176 54352 17196
rect 54352 17176 54354 17196
rect 55770 17076 55772 17096
rect 55772 17076 55824 17096
rect 55824 17076 55826 17096
rect 55770 17040 55826 17076
rect 57242 44648 57298 44704
rect 57058 42472 57114 42528
rect 57334 41520 57390 41576
rect 57242 41384 57298 41440
rect 57058 40296 57114 40352
rect 57058 39208 57114 39264
rect 57058 32680 57114 32736
rect 57058 29416 57114 29472
rect 57242 18536 57298 18592
rect 57058 16360 57114 16416
rect 56966 13096 57022 13152
rect 57150 15408 57206 15464
rect 57334 16904 57390 16960
rect 57886 49544 57942 49600
rect 57978 49000 58034 49056
rect 58162 56616 58218 56672
rect 58162 47912 58218 47968
rect 58070 47368 58126 47424
rect 58162 46280 58218 46336
rect 58070 45736 58126 45792
rect 57886 44104 57942 44160
rect 58162 43016 58218 43072
rect 57978 41928 58034 41984
rect 57886 40840 57942 40896
rect 57886 39752 57942 39808
rect 57978 38664 58034 38720
rect 58162 38120 58218 38176
rect 58070 37576 58126 37632
rect 58162 36488 58218 36544
rect 57978 35944 58034 36000
rect 58162 34856 58218 34912
rect 57886 34312 57942 34368
rect 58162 33224 58218 33280
rect 58346 56072 58402 56128
rect 58346 54440 58402 54496
rect 58346 52844 58348 52864
rect 58348 52844 58400 52864
rect 58400 52844 58402 52864
rect 58346 52808 58402 52844
rect 58346 51176 58402 51232
rect 58162 31592 58218 31648
rect 58070 31048 58126 31104
rect 58162 29960 58218 30016
rect 58162 28328 58218 28384
rect 57978 27784 58034 27840
rect 58162 26696 58218 26752
rect 58070 26152 58126 26208
rect 58162 25064 58218 25120
rect 58070 24520 58126 24576
rect 58162 23432 58218 23488
rect 58162 22888 58218 22944
rect 58162 21800 58218 21856
rect 58070 21256 58126 21312
rect 58162 20168 58218 20224
rect 57978 19624 58034 19680
rect 57978 17992 58034 18048
rect 57978 14728 58034 14784
rect 58162 15272 58218 15328
rect 58070 13776 58126 13832
rect 58162 13640 58218 13696
rect 57150 11464 57206 11520
rect 58162 12008 58218 12064
rect 58162 10376 58218 10432
rect 57058 9832 57114 9888
rect 56230 8200 56286 8256
rect 57334 8744 57390 8800
rect 57150 6568 57206 6624
rect 57058 6160 57114 6216
rect 58162 7112 58218 7168
rect 57242 5480 57298 5536
rect 58070 4936 58126 4992
rect 57334 2216 57390 2272
rect 57886 3848 57942 3904
rect 58162 3304 58218 3360
rect 58162 2760 58218 2816
rect 57794 1672 57850 1728
rect 55954 1128 56010 1184
<< metal3 >>
rect 56409 62658 56475 62661
rect 59200 62658 60000 62688
rect 56409 62656 60000 62658
rect 56409 62600 56414 62656
rect 56470 62600 60000 62656
rect 56409 62598 60000 62600
rect 56409 62595 56475 62598
rect 59200 62568 60000 62598
rect 56133 62114 56199 62117
rect 59200 62114 60000 62144
rect 56133 62112 60000 62114
rect 56133 62056 56138 62112
rect 56194 62056 60000 62112
rect 56133 62054 60000 62056
rect 56133 62051 56199 62054
rect 59200 62024 60000 62054
rect 0 61842 800 61872
rect 1669 61842 1735 61845
rect 0 61840 1735 61842
rect 0 61784 1674 61840
rect 1730 61784 1735 61840
rect 0 61782 1735 61784
rect 0 61752 800 61782
rect 1669 61779 1735 61782
rect 55397 61570 55463 61573
rect 59200 61570 60000 61600
rect 55397 61568 60000 61570
rect 55397 61512 55402 61568
rect 55458 61512 60000 61568
rect 55397 61510 60000 61512
rect 55397 61507 55463 61510
rect 4210 61504 4526 61505
rect 4210 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4526 61504
rect 4210 61439 4526 61440
rect 34930 61504 35246 61505
rect 34930 61440 34936 61504
rect 35000 61440 35016 61504
rect 35080 61440 35096 61504
rect 35160 61440 35176 61504
rect 35240 61440 35246 61504
rect 59200 61480 60000 61510
rect 34930 61439 35246 61440
rect 0 61162 800 61192
rect 2773 61162 2839 61165
rect 0 61160 2839 61162
rect 0 61104 2778 61160
rect 2834 61104 2839 61160
rect 0 61102 2839 61104
rect 0 61072 800 61102
rect 2773 61099 2839 61102
rect 12985 61162 13051 61165
rect 28574 61162 28580 61164
rect 12985 61160 28580 61162
rect 12985 61104 12990 61160
rect 13046 61104 28580 61160
rect 12985 61102 28580 61104
rect 12985 61099 13051 61102
rect 28574 61100 28580 61102
rect 28644 61100 28650 61164
rect 30046 61100 30052 61164
rect 30116 61162 30122 61164
rect 53373 61162 53439 61165
rect 30116 61160 53439 61162
rect 30116 61104 53378 61160
rect 53434 61104 53439 61160
rect 30116 61102 53439 61104
rect 30116 61100 30122 61102
rect 53373 61099 53439 61102
rect 56501 61026 56567 61029
rect 59200 61026 60000 61056
rect 56501 61024 60000 61026
rect 56501 60968 56506 61024
rect 56562 60968 60000 61024
rect 56501 60966 60000 60968
rect 56501 60963 56567 60966
rect 19570 60960 19886 60961
rect 19570 60896 19576 60960
rect 19640 60896 19656 60960
rect 19720 60896 19736 60960
rect 19800 60896 19816 60960
rect 19880 60896 19886 60960
rect 19570 60895 19886 60896
rect 50290 60960 50606 60961
rect 50290 60896 50296 60960
rect 50360 60896 50376 60960
rect 50440 60896 50456 60960
rect 50520 60896 50536 60960
rect 50600 60896 50606 60960
rect 59200 60936 60000 60966
rect 50290 60895 50606 60896
rect 22737 60754 22803 60757
rect 28758 60754 28764 60756
rect 22737 60752 28764 60754
rect 22737 60696 22742 60752
rect 22798 60696 28764 60752
rect 22737 60694 28764 60696
rect 22737 60691 22803 60694
rect 28758 60692 28764 60694
rect 28828 60692 28834 60756
rect 0 60482 800 60512
rect 1577 60482 1643 60485
rect 0 60480 1643 60482
rect 0 60424 1582 60480
rect 1638 60424 1643 60480
rect 0 60422 1643 60424
rect 0 60392 800 60422
rect 1577 60419 1643 60422
rect 57237 60482 57303 60485
rect 59200 60482 60000 60512
rect 57237 60480 60000 60482
rect 57237 60424 57242 60480
rect 57298 60424 60000 60480
rect 57237 60422 60000 60424
rect 57237 60419 57303 60422
rect 4210 60416 4526 60417
rect 4210 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4526 60416
rect 4210 60351 4526 60352
rect 34930 60416 35246 60417
rect 34930 60352 34936 60416
rect 35000 60352 35016 60416
rect 35080 60352 35096 60416
rect 35160 60352 35176 60416
rect 35240 60352 35246 60416
rect 59200 60392 60000 60422
rect 34930 60351 35246 60352
rect 22093 60346 22159 60349
rect 22553 60348 22619 60349
rect 22502 60346 22508 60348
rect 22093 60344 22508 60346
rect 22572 60346 22619 60348
rect 22572 60344 22700 60346
rect 22093 60288 22098 60344
rect 22154 60288 22508 60344
rect 22614 60288 22700 60344
rect 22093 60286 22508 60288
rect 22093 60283 22159 60286
rect 22502 60284 22508 60286
rect 22572 60286 22700 60288
rect 22572 60284 22619 60286
rect 22553 60283 22619 60284
rect 22093 60210 22159 60213
rect 58249 60210 58315 60213
rect 22093 60208 58315 60210
rect 22093 60152 22098 60208
rect 22154 60152 58254 60208
rect 58310 60152 58315 60208
rect 22093 60150 58315 60152
rect 22093 60147 22159 60150
rect 58249 60147 58315 60150
rect 30373 60074 30439 60077
rect 40534 60074 40540 60076
rect 30373 60072 40540 60074
rect 30373 60016 30378 60072
rect 30434 60016 40540 60072
rect 30373 60014 40540 60016
rect 30373 60011 30439 60014
rect 40534 60012 40540 60014
rect 40604 60012 40610 60076
rect 30649 59938 30715 59941
rect 32673 59938 32739 59941
rect 30649 59936 32739 59938
rect 30649 59880 30654 59936
rect 30710 59880 32678 59936
rect 32734 59880 32739 59936
rect 30649 59878 32739 59880
rect 30649 59875 30715 59878
rect 32673 59875 32739 59878
rect 58065 59938 58131 59941
rect 59200 59938 60000 59968
rect 58065 59936 60000 59938
rect 58065 59880 58070 59936
rect 58126 59880 60000 59936
rect 58065 59878 60000 59880
rect 58065 59875 58131 59878
rect 19570 59872 19886 59873
rect 0 59802 800 59832
rect 19570 59808 19576 59872
rect 19640 59808 19656 59872
rect 19720 59808 19736 59872
rect 19800 59808 19816 59872
rect 19880 59808 19886 59872
rect 19570 59807 19886 59808
rect 50290 59872 50606 59873
rect 50290 59808 50296 59872
rect 50360 59808 50376 59872
rect 50440 59808 50456 59872
rect 50520 59808 50536 59872
rect 50600 59808 50606 59872
rect 59200 59848 60000 59878
rect 50290 59807 50606 59808
rect 1669 59802 1735 59805
rect 0 59800 1735 59802
rect 0 59744 1674 59800
rect 1730 59744 1735 59800
rect 0 59742 1735 59744
rect 0 59712 800 59742
rect 1669 59739 1735 59742
rect 22001 59666 22067 59669
rect 22737 59666 22803 59669
rect 23381 59666 23447 59669
rect 28625 59666 28691 59669
rect 22001 59664 28691 59666
rect 22001 59608 22006 59664
rect 22062 59608 22742 59664
rect 22798 59608 23386 59664
rect 23442 59608 28630 59664
rect 28686 59608 28691 59664
rect 22001 59606 28691 59608
rect 22001 59603 22067 59606
rect 22737 59603 22803 59606
rect 23381 59603 23447 59606
rect 28625 59603 28691 59606
rect 18597 59394 18663 59397
rect 19190 59394 19196 59396
rect 18597 59392 19196 59394
rect 18597 59336 18602 59392
rect 18658 59336 19196 59392
rect 18597 59334 19196 59336
rect 18597 59331 18663 59334
rect 19190 59332 19196 59334
rect 19260 59332 19266 59396
rect 41965 59394 42031 59397
rect 42558 59394 42564 59396
rect 41965 59392 42564 59394
rect 41965 59336 41970 59392
rect 42026 59336 42564 59392
rect 41965 59334 42564 59336
rect 41965 59331 42031 59334
rect 42558 59332 42564 59334
rect 42628 59332 42634 59396
rect 58065 59394 58131 59397
rect 59200 59394 60000 59424
rect 58065 59392 60000 59394
rect 58065 59336 58070 59392
rect 58126 59336 60000 59392
rect 58065 59334 60000 59336
rect 58065 59331 58131 59334
rect 4210 59328 4526 59329
rect 4210 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4526 59328
rect 4210 59263 4526 59264
rect 34930 59328 35246 59329
rect 34930 59264 34936 59328
rect 35000 59264 35016 59328
rect 35080 59264 35096 59328
rect 35160 59264 35176 59328
rect 35240 59264 35246 59328
rect 59200 59304 60000 59334
rect 34930 59263 35246 59264
rect 0 59122 800 59152
rect 1669 59122 1735 59125
rect 0 59120 1735 59122
rect 0 59064 1674 59120
rect 1730 59064 1735 59120
rect 0 59062 1735 59064
rect 0 59032 800 59062
rect 1669 59059 1735 59062
rect 39246 58924 39252 58988
rect 39316 58986 39322 58988
rect 58065 58986 58131 58989
rect 39316 58984 58131 58986
rect 39316 58928 58070 58984
rect 58126 58928 58131 58984
rect 39316 58926 58131 58928
rect 39316 58924 39322 58926
rect 58065 58923 58131 58926
rect 58157 58850 58223 58853
rect 59200 58850 60000 58880
rect 58157 58848 60000 58850
rect 58157 58792 58162 58848
rect 58218 58792 60000 58848
rect 58157 58790 60000 58792
rect 58157 58787 58223 58790
rect 19570 58784 19886 58785
rect 19570 58720 19576 58784
rect 19640 58720 19656 58784
rect 19720 58720 19736 58784
rect 19800 58720 19816 58784
rect 19880 58720 19886 58784
rect 19570 58719 19886 58720
rect 50290 58784 50606 58785
rect 50290 58720 50296 58784
rect 50360 58720 50376 58784
rect 50440 58720 50456 58784
rect 50520 58720 50536 58784
rect 50600 58720 50606 58784
rect 59200 58760 60000 58790
rect 50290 58719 50606 58720
rect 0 58442 800 58472
rect 1577 58442 1643 58445
rect 0 58440 1643 58442
rect 0 58384 1582 58440
rect 1638 58384 1643 58440
rect 0 58382 1643 58384
rect 0 58352 800 58382
rect 1577 58379 1643 58382
rect 57881 58306 57947 58309
rect 59200 58306 60000 58336
rect 57881 58304 60000 58306
rect 57881 58248 57886 58304
rect 57942 58248 60000 58304
rect 57881 58246 60000 58248
rect 57881 58243 57947 58246
rect 4210 58240 4526 58241
rect 4210 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4526 58240
rect 4210 58175 4526 58176
rect 34930 58240 35246 58241
rect 34930 58176 34936 58240
rect 35000 58176 35016 58240
rect 35080 58176 35096 58240
rect 35160 58176 35176 58240
rect 35240 58176 35246 58240
rect 59200 58216 60000 58246
rect 34930 58175 35246 58176
rect 0 57762 800 57792
rect 1577 57762 1643 57765
rect 0 57760 1643 57762
rect 0 57704 1582 57760
rect 1638 57704 1643 57760
rect 0 57702 1643 57704
rect 0 57672 800 57702
rect 1577 57699 1643 57702
rect 57973 57762 58039 57765
rect 59200 57762 60000 57792
rect 57973 57760 60000 57762
rect 57973 57704 57978 57760
rect 58034 57704 60000 57760
rect 57973 57702 60000 57704
rect 57973 57699 58039 57702
rect 19570 57696 19886 57697
rect 19570 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19886 57696
rect 19570 57631 19886 57632
rect 50290 57696 50606 57697
rect 50290 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50606 57696
rect 59200 57672 60000 57702
rect 50290 57631 50606 57632
rect 42701 57354 42767 57357
rect 43662 57354 43668 57356
rect 42701 57352 43668 57354
rect 42701 57296 42706 57352
rect 42762 57296 43668 57352
rect 42701 57294 43668 57296
rect 42701 57291 42767 57294
rect 43662 57292 43668 57294
rect 43732 57292 43738 57356
rect 57881 57218 57947 57221
rect 59200 57218 60000 57248
rect 57881 57216 60000 57218
rect 57881 57160 57886 57216
rect 57942 57160 60000 57216
rect 57881 57158 60000 57160
rect 57881 57155 57947 57158
rect 4210 57152 4526 57153
rect 0 57082 800 57112
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 34930 57152 35246 57153
rect 34930 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35246 57152
rect 59200 57128 60000 57158
rect 34930 57087 35246 57088
rect 1577 57082 1643 57085
rect 0 57080 1643 57082
rect 0 57024 1582 57080
rect 1638 57024 1643 57080
rect 0 57022 1643 57024
rect 0 56992 800 57022
rect 1577 57019 1643 57022
rect 58157 56674 58223 56677
rect 59200 56674 60000 56704
rect 58157 56672 60000 56674
rect 58157 56616 58162 56672
rect 58218 56616 60000 56672
rect 58157 56614 60000 56616
rect 58157 56611 58223 56614
rect 19570 56608 19886 56609
rect 19570 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19886 56608
rect 19570 56543 19886 56544
rect 50290 56608 50606 56609
rect 50290 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50606 56608
rect 59200 56584 60000 56614
rect 50290 56543 50606 56544
rect 0 56402 800 56432
rect 1669 56402 1735 56405
rect 0 56400 1735 56402
rect 0 56344 1674 56400
rect 1730 56344 1735 56400
rect 0 56342 1735 56344
rect 0 56312 800 56342
rect 1669 56339 1735 56342
rect 58341 56130 58407 56133
rect 59200 56130 60000 56160
rect 58341 56128 60000 56130
rect 58341 56072 58346 56128
rect 58402 56072 60000 56128
rect 58341 56070 60000 56072
rect 58341 56067 58407 56070
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 34930 56064 35246 56065
rect 34930 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35246 56064
rect 59200 56040 60000 56070
rect 34930 55999 35246 56000
rect 0 55722 800 55752
rect 1669 55722 1735 55725
rect 0 55720 1735 55722
rect 0 55664 1674 55720
rect 1730 55664 1735 55720
rect 0 55662 1735 55664
rect 0 55632 800 55662
rect 1669 55659 1735 55662
rect 19570 55520 19886 55521
rect 19570 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19886 55520
rect 19570 55455 19886 55456
rect 50290 55520 50606 55521
rect 50290 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50606 55520
rect 59200 55496 60000 55616
rect 50290 55455 50606 55456
rect 0 55042 800 55072
rect 1577 55042 1643 55045
rect 0 55040 1643 55042
rect 0 54984 1582 55040
rect 1638 54984 1643 55040
rect 0 54982 1643 54984
rect 0 54952 800 54982
rect 1577 54979 1643 54982
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 59200 54952 60000 55072
rect 34930 54911 35246 54912
rect 58341 54498 58407 54501
rect 59200 54498 60000 54528
rect 58341 54496 60000 54498
rect 58341 54440 58346 54496
rect 58402 54440 60000 54496
rect 58341 54438 60000 54440
rect 58341 54435 58407 54438
rect 19570 54432 19886 54433
rect 0 54362 800 54392
rect 19570 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19886 54432
rect 19570 54367 19886 54368
rect 50290 54432 50606 54433
rect 50290 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50606 54432
rect 59200 54408 60000 54438
rect 50290 54367 50606 54368
rect 1669 54362 1735 54365
rect 0 54360 1735 54362
rect 0 54304 1674 54360
rect 1730 54304 1735 54360
rect 0 54302 1735 54304
rect 0 54272 800 54302
rect 1669 54299 1735 54302
rect 22829 53956 22895 53957
rect 22829 53952 22876 53956
rect 22940 53954 22946 53956
rect 22829 53896 22834 53952
rect 22829 53892 22876 53896
rect 22940 53894 22986 53954
rect 22940 53892 22946 53894
rect 22829 53891 22895 53892
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 59200 53864 60000 53984
rect 34930 53823 35246 53824
rect 0 53682 800 53712
rect 1577 53682 1643 53685
rect 0 53680 1643 53682
rect 0 53624 1582 53680
rect 1638 53624 1643 53680
rect 0 53622 1643 53624
rect 0 53592 800 53622
rect 1577 53619 1643 53622
rect 19570 53344 19886 53345
rect 19570 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19886 53344
rect 19570 53279 19886 53280
rect 50290 53344 50606 53345
rect 50290 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50606 53344
rect 59200 53320 60000 53440
rect 50290 53279 50606 53280
rect 0 53002 800 53032
rect 1669 53002 1735 53005
rect 0 53000 1735 53002
rect 0 52944 1674 53000
rect 1730 52944 1735 53000
rect 0 52942 1735 52944
rect 0 52912 800 52942
rect 1669 52939 1735 52942
rect 58341 52866 58407 52869
rect 59200 52866 60000 52896
rect 58341 52864 60000 52866
rect 58341 52808 58346 52864
rect 58402 52808 60000 52864
rect 58341 52806 60000 52808
rect 58341 52803 58407 52806
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 59200 52776 60000 52806
rect 34930 52735 35246 52736
rect 0 52322 800 52352
rect 1577 52322 1643 52325
rect 0 52320 1643 52322
rect 0 52264 1582 52320
rect 1638 52264 1643 52320
rect 0 52262 1643 52264
rect 0 52232 800 52262
rect 1577 52259 1643 52262
rect 19570 52256 19886 52257
rect 19570 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19886 52256
rect 19570 52191 19886 52192
rect 50290 52256 50606 52257
rect 50290 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50606 52256
rect 59200 52232 60000 52352
rect 50290 52191 50606 52192
rect 4210 51712 4526 51713
rect 0 51642 800 51672
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 59200 51688 60000 51808
rect 34930 51647 35246 51648
rect 1669 51642 1735 51645
rect 0 51640 1735 51642
rect 0 51584 1674 51640
rect 1730 51584 1735 51640
rect 0 51582 1735 51584
rect 0 51552 800 51582
rect 1669 51579 1735 51582
rect 58341 51234 58407 51237
rect 59200 51234 60000 51264
rect 58341 51232 60000 51234
rect 58341 51176 58346 51232
rect 58402 51176 60000 51232
rect 58341 51174 60000 51176
rect 58341 51171 58407 51174
rect 19570 51168 19886 51169
rect 19570 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19886 51168
rect 19570 51103 19886 51104
rect 50290 51168 50606 51169
rect 50290 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50606 51168
rect 59200 51144 60000 51174
rect 50290 51103 50606 51104
rect 0 50962 800 50992
rect 1669 50962 1735 50965
rect 0 50960 1735 50962
rect 0 50904 1674 50960
rect 1730 50904 1735 50960
rect 0 50902 1735 50904
rect 0 50872 800 50902
rect 1669 50899 1735 50902
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 59200 50600 60000 50720
rect 34930 50559 35246 50560
rect 0 50282 800 50312
rect 1669 50282 1735 50285
rect 0 50280 1735 50282
rect 0 50224 1674 50280
rect 1730 50224 1735 50280
rect 0 50222 1735 50224
rect 0 50192 800 50222
rect 1669 50219 1735 50222
rect 17493 50282 17559 50285
rect 36302 50282 36308 50284
rect 17493 50280 36308 50282
rect 17493 50224 17498 50280
rect 17554 50224 36308 50280
rect 17493 50222 36308 50224
rect 17493 50219 17559 50222
rect 36302 50220 36308 50222
rect 36372 50220 36378 50284
rect 19570 50080 19886 50081
rect 19570 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19886 50080
rect 19570 50015 19886 50016
rect 50290 50080 50606 50081
rect 50290 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50606 50080
rect 59200 50056 60000 50176
rect 50290 50015 50606 50016
rect 0 49602 800 49632
rect 1577 49602 1643 49605
rect 0 49600 1643 49602
rect 0 49544 1582 49600
rect 1638 49544 1643 49600
rect 0 49542 1643 49544
rect 0 49512 800 49542
rect 1577 49539 1643 49542
rect 57881 49602 57947 49605
rect 59200 49602 60000 49632
rect 57881 49600 60000 49602
rect 57881 49544 57886 49600
rect 57942 49544 60000 49600
rect 57881 49542 60000 49544
rect 57881 49539 57947 49542
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 59200 49512 60000 49542
rect 34930 49471 35246 49472
rect 57973 49058 58039 49061
rect 59200 49058 60000 49088
rect 57973 49056 60000 49058
rect 57973 49000 57978 49056
rect 58034 49000 60000 49056
rect 57973 48998 60000 49000
rect 57973 48995 58039 48998
rect 19570 48992 19886 48993
rect 0 48922 800 48952
rect 19570 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19886 48992
rect 19570 48927 19886 48928
rect 50290 48992 50606 48993
rect 50290 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50606 48992
rect 59200 48968 60000 48998
rect 50290 48927 50606 48928
rect 1577 48922 1643 48925
rect 0 48920 1643 48922
rect 0 48864 1582 48920
rect 1638 48864 1643 48920
rect 0 48862 1643 48864
rect 0 48832 800 48862
rect 1577 48859 1643 48862
rect 27337 48922 27403 48925
rect 42926 48922 42932 48924
rect 27337 48920 42932 48922
rect 27337 48864 27342 48920
rect 27398 48864 42932 48920
rect 27337 48862 42932 48864
rect 27337 48859 27403 48862
rect 42926 48860 42932 48862
rect 42996 48860 43002 48924
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 59200 48424 60000 48544
rect 34930 48383 35246 48384
rect 0 48242 800 48272
rect 1669 48242 1735 48245
rect 0 48240 1735 48242
rect 0 48184 1674 48240
rect 1730 48184 1735 48240
rect 0 48182 1735 48184
rect 0 48152 800 48182
rect 1669 48179 1735 48182
rect 58157 47970 58223 47973
rect 59200 47970 60000 48000
rect 58157 47968 60000 47970
rect 58157 47912 58162 47968
rect 58218 47912 60000 47968
rect 58157 47910 60000 47912
rect 58157 47907 58223 47910
rect 19570 47904 19886 47905
rect 19570 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19886 47904
rect 19570 47839 19886 47840
rect 50290 47904 50606 47905
rect 50290 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50606 47904
rect 59200 47880 60000 47910
rect 50290 47839 50606 47840
rect 0 47562 800 47592
rect 1669 47562 1735 47565
rect 0 47560 1735 47562
rect 0 47504 1674 47560
rect 1730 47504 1735 47560
rect 0 47502 1735 47504
rect 0 47472 800 47502
rect 1669 47499 1735 47502
rect 58065 47426 58131 47429
rect 59200 47426 60000 47456
rect 58065 47424 60000 47426
rect 58065 47368 58070 47424
rect 58126 47368 60000 47424
rect 58065 47366 60000 47368
rect 58065 47363 58131 47366
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 59200 47336 60000 47366
rect 34930 47295 35246 47296
rect 0 46882 800 46912
rect 1577 46882 1643 46885
rect 0 46880 1643 46882
rect 0 46824 1582 46880
rect 1638 46824 1643 46880
rect 0 46822 1643 46824
rect 0 46792 800 46822
rect 1577 46819 1643 46822
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 50290 46816 50606 46817
rect 50290 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50606 46816
rect 59200 46792 60000 46912
rect 50290 46751 50606 46752
rect 58157 46338 58223 46341
rect 59200 46338 60000 46368
rect 58157 46336 60000 46338
rect 58157 46280 58162 46336
rect 58218 46280 60000 46336
rect 58157 46278 60000 46280
rect 58157 46275 58223 46278
rect 4210 46272 4526 46273
rect 0 46202 800 46232
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 59200 46248 60000 46278
rect 34930 46207 35246 46208
rect 1577 46202 1643 46205
rect 0 46200 1643 46202
rect 0 46144 1582 46200
rect 1638 46144 1643 46200
rect 0 46142 1643 46144
rect 0 46112 800 46142
rect 1577 46139 1643 46142
rect 58065 45794 58131 45797
rect 59200 45794 60000 45824
rect 58065 45792 60000 45794
rect 58065 45736 58070 45792
rect 58126 45736 60000 45792
rect 58065 45734 60000 45736
rect 58065 45731 58131 45734
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 50290 45728 50606 45729
rect 50290 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50606 45728
rect 59200 45704 60000 45734
rect 50290 45663 50606 45664
rect 0 45522 800 45552
rect 1669 45522 1735 45525
rect 0 45520 1735 45522
rect 0 45464 1674 45520
rect 1730 45464 1735 45520
rect 0 45462 1735 45464
rect 0 45432 800 45462
rect 1669 45459 1735 45462
rect 38009 45386 38075 45389
rect 38142 45386 38148 45388
rect 38009 45384 38148 45386
rect 38009 45328 38014 45384
rect 38070 45328 38148 45384
rect 38009 45326 38148 45328
rect 38009 45323 38075 45326
rect 38142 45324 38148 45326
rect 38212 45324 38218 45388
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 59200 45160 60000 45280
rect 34930 45119 35246 45120
rect 0 44842 800 44872
rect 1577 44842 1643 44845
rect 0 44840 1643 44842
rect 0 44784 1582 44840
rect 1638 44784 1643 44840
rect 0 44782 1643 44784
rect 0 44752 800 44782
rect 1577 44779 1643 44782
rect 57237 44706 57303 44709
rect 59200 44706 60000 44736
rect 57237 44704 60000 44706
rect 57237 44648 57242 44704
rect 57298 44648 60000 44704
rect 57237 44646 60000 44648
rect 57237 44643 57303 44646
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 50290 44640 50606 44641
rect 50290 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50606 44640
rect 59200 44616 60000 44646
rect 50290 44575 50606 44576
rect 0 44162 800 44192
rect 1669 44162 1735 44165
rect 0 44160 1735 44162
rect 0 44104 1674 44160
rect 1730 44104 1735 44160
rect 0 44102 1735 44104
rect 0 44072 800 44102
rect 1669 44099 1735 44102
rect 57881 44162 57947 44165
rect 59200 44162 60000 44192
rect 57881 44160 60000 44162
rect 57881 44104 57886 44160
rect 57942 44104 60000 44160
rect 57881 44102 60000 44104
rect 57881 44099 57947 44102
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 59200 44072 60000 44102
rect 34930 44031 35246 44032
rect 19570 43552 19886 43553
rect 0 43482 800 43512
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 50290 43552 50606 43553
rect 50290 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50606 43552
rect 59200 43528 60000 43648
rect 50290 43487 50606 43488
rect 1669 43482 1735 43485
rect 0 43480 1735 43482
rect 0 43424 1674 43480
rect 1730 43424 1735 43480
rect 0 43422 1735 43424
rect 0 43392 800 43422
rect 1669 43419 1735 43422
rect 27286 43148 27292 43212
rect 27356 43210 27362 43212
rect 32765 43210 32831 43213
rect 27356 43208 32831 43210
rect 27356 43152 32770 43208
rect 32826 43152 32831 43208
rect 27356 43150 32831 43152
rect 27356 43148 27362 43150
rect 32765 43147 32831 43150
rect 58157 43074 58223 43077
rect 59200 43074 60000 43104
rect 58157 43072 60000 43074
rect 58157 43016 58162 43072
rect 58218 43016 60000 43072
rect 58157 43014 60000 43016
rect 58157 43011 58223 43014
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 59200 42984 60000 43014
rect 34930 42943 35246 42944
rect 0 42802 800 42832
rect 1577 42802 1643 42805
rect 0 42800 1643 42802
rect 0 42744 1582 42800
rect 1638 42744 1643 42800
rect 0 42742 1643 42744
rect 0 42712 800 42742
rect 1577 42739 1643 42742
rect 37273 42666 37339 42669
rect 37406 42666 37412 42668
rect 37273 42664 37412 42666
rect 37273 42608 37278 42664
rect 37334 42608 37412 42664
rect 37273 42606 37412 42608
rect 37273 42603 37339 42606
rect 37406 42604 37412 42606
rect 37476 42604 37482 42668
rect 57053 42530 57119 42533
rect 59200 42530 60000 42560
rect 57053 42528 60000 42530
rect 57053 42472 57058 42528
rect 57114 42472 60000 42528
rect 57053 42470 60000 42472
rect 57053 42467 57119 42470
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 50290 42464 50606 42465
rect 50290 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50606 42464
rect 59200 42440 60000 42470
rect 50290 42399 50606 42400
rect 0 42122 800 42152
rect 1577 42122 1643 42125
rect 0 42120 1643 42122
rect 0 42064 1582 42120
rect 1638 42064 1643 42120
rect 0 42062 1643 42064
rect 0 42032 800 42062
rect 1577 42059 1643 42062
rect 15285 42122 15351 42125
rect 39062 42122 39068 42124
rect 15285 42120 39068 42122
rect 15285 42064 15290 42120
rect 15346 42064 39068 42120
rect 15285 42062 39068 42064
rect 15285 42059 15351 42062
rect 39062 42060 39068 42062
rect 39132 42060 39138 42124
rect 57973 41986 58039 41989
rect 59200 41986 60000 42016
rect 57973 41984 60000 41986
rect 57973 41928 57978 41984
rect 58034 41928 60000 41984
rect 57973 41926 60000 41928
rect 57973 41923 58039 41926
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 59200 41896 60000 41926
rect 34930 41855 35246 41856
rect 57329 41580 57395 41581
rect 57278 41578 57284 41580
rect 57238 41518 57284 41578
rect 57348 41576 57395 41580
rect 57390 41520 57395 41576
rect 57278 41516 57284 41518
rect 57348 41516 57395 41520
rect 57329 41515 57395 41516
rect 0 41442 800 41472
rect 1669 41442 1735 41445
rect 0 41440 1735 41442
rect 0 41384 1674 41440
rect 1730 41384 1735 41440
rect 0 41382 1735 41384
rect 0 41352 800 41382
rect 1669 41379 1735 41382
rect 57237 41442 57303 41445
rect 59200 41442 60000 41472
rect 57237 41440 60000 41442
rect 57237 41384 57242 41440
rect 57298 41384 60000 41440
rect 57237 41382 60000 41384
rect 57237 41379 57303 41382
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 50290 41376 50606 41377
rect 50290 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50606 41376
rect 59200 41352 60000 41382
rect 50290 41311 50606 41312
rect 57881 40898 57947 40901
rect 59200 40898 60000 40928
rect 57881 40896 60000 40898
rect 57881 40840 57886 40896
rect 57942 40840 60000 40896
rect 57881 40838 60000 40840
rect 57881 40835 57947 40838
rect 4210 40832 4526 40833
rect 0 40762 800 40792
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 59200 40808 60000 40838
rect 34930 40767 35246 40768
rect 1669 40762 1735 40765
rect 0 40760 1735 40762
rect 0 40704 1674 40760
rect 1730 40704 1735 40760
rect 0 40702 1735 40704
rect 0 40672 800 40702
rect 1669 40699 1735 40702
rect 57053 40354 57119 40357
rect 59200 40354 60000 40384
rect 57053 40352 60000 40354
rect 57053 40296 57058 40352
rect 57114 40296 60000 40352
rect 57053 40294 60000 40296
rect 57053 40291 57119 40294
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 50290 40288 50606 40289
rect 50290 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50606 40288
rect 59200 40264 60000 40294
rect 50290 40223 50606 40224
rect 0 40082 800 40112
rect 1669 40082 1735 40085
rect 0 40080 1735 40082
rect 0 40024 1674 40080
rect 1730 40024 1735 40080
rect 0 40022 1735 40024
rect 0 39992 800 40022
rect 1669 40019 1735 40022
rect 57881 39810 57947 39813
rect 59200 39810 60000 39840
rect 57881 39808 60000 39810
rect 57881 39752 57886 39808
rect 57942 39752 60000 39808
rect 57881 39750 60000 39752
rect 57881 39747 57947 39750
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 59200 39720 60000 39750
rect 34930 39679 35246 39680
rect 0 39402 800 39432
rect 1669 39402 1735 39405
rect 0 39400 1735 39402
rect 0 39344 1674 39400
rect 1730 39344 1735 39400
rect 0 39342 1735 39344
rect 0 39312 800 39342
rect 1669 39339 1735 39342
rect 57053 39266 57119 39269
rect 59200 39266 60000 39296
rect 57053 39264 60000 39266
rect 57053 39208 57058 39264
rect 57114 39208 60000 39264
rect 57053 39206 60000 39208
rect 57053 39203 57119 39206
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 59200 39176 60000 39206
rect 50290 39135 50606 39136
rect 0 38722 800 38752
rect 1669 38722 1735 38725
rect 0 38720 1735 38722
rect 0 38664 1674 38720
rect 1730 38664 1735 38720
rect 0 38662 1735 38664
rect 0 38632 800 38662
rect 1669 38659 1735 38662
rect 57973 38722 58039 38725
rect 59200 38722 60000 38752
rect 57973 38720 60000 38722
rect 57973 38664 57978 38720
rect 58034 38664 60000 38720
rect 57973 38662 60000 38664
rect 57973 38659 58039 38662
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 59200 38632 60000 38662
rect 34930 38591 35246 38592
rect 58157 38178 58223 38181
rect 59200 38178 60000 38208
rect 58157 38176 60000 38178
rect 58157 38120 58162 38176
rect 58218 38120 60000 38176
rect 58157 38118 60000 38120
rect 58157 38115 58223 38118
rect 19570 38112 19886 38113
rect 0 38042 800 38072
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 59200 38088 60000 38118
rect 50290 38047 50606 38048
rect 1669 38042 1735 38045
rect 0 38040 1735 38042
rect 0 37984 1674 38040
rect 1730 37984 1735 38040
rect 0 37982 1735 37984
rect 0 37952 800 37982
rect 1669 37979 1735 37982
rect 20713 37906 20779 37909
rect 22921 37906 22987 37909
rect 20713 37904 22987 37906
rect 20713 37848 20718 37904
rect 20774 37848 22926 37904
rect 22982 37848 22987 37904
rect 20713 37846 22987 37848
rect 20713 37843 20779 37846
rect 22921 37843 22987 37846
rect 22553 37770 22619 37773
rect 23013 37770 23079 37773
rect 40718 37770 40724 37772
rect 22553 37768 40724 37770
rect 22553 37712 22558 37768
rect 22614 37712 23018 37768
rect 23074 37712 40724 37768
rect 22553 37710 40724 37712
rect 22553 37707 22619 37710
rect 23013 37707 23079 37710
rect 40718 37708 40724 37710
rect 40788 37708 40794 37772
rect 58065 37634 58131 37637
rect 59200 37634 60000 37664
rect 58065 37632 60000 37634
rect 58065 37576 58070 37632
rect 58126 37576 60000 37632
rect 58065 37574 60000 37576
rect 58065 37571 58131 37574
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 59200 37544 60000 37574
rect 34930 37503 35246 37504
rect 0 37362 800 37392
rect 1669 37362 1735 37365
rect 0 37360 1735 37362
rect 0 37304 1674 37360
rect 1730 37304 1735 37360
rect 0 37302 1735 37304
rect 0 37272 800 37302
rect 1669 37299 1735 37302
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 59200 37000 60000 37120
rect 50290 36959 50606 36960
rect 0 36682 800 36712
rect 1577 36682 1643 36685
rect 0 36680 1643 36682
rect 0 36624 1582 36680
rect 1638 36624 1643 36680
rect 0 36622 1643 36624
rect 0 36592 800 36622
rect 1577 36619 1643 36622
rect 58157 36546 58223 36549
rect 59200 36546 60000 36576
rect 58157 36544 60000 36546
rect 58157 36488 58162 36544
rect 58218 36488 60000 36544
rect 58157 36486 60000 36488
rect 58157 36483 58223 36486
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 59200 36456 60000 36486
rect 34930 36415 35246 36416
rect 0 36002 800 36032
rect 1669 36002 1735 36005
rect 0 36000 1735 36002
rect 0 35944 1674 36000
rect 1730 35944 1735 36000
rect 0 35942 1735 35944
rect 0 35912 800 35942
rect 1669 35939 1735 35942
rect 57973 36002 58039 36005
rect 59200 36002 60000 36032
rect 57973 36000 60000 36002
rect 57973 35944 57978 36000
rect 58034 35944 60000 36000
rect 57973 35942 60000 35944
rect 57973 35939 58039 35942
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 59200 35912 60000 35942
rect 50290 35871 50606 35872
rect 4210 35392 4526 35393
rect 0 35322 800 35352
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 59200 35368 60000 35488
rect 34930 35327 35246 35328
rect 1669 35322 1735 35325
rect 0 35320 1735 35322
rect 0 35264 1674 35320
rect 1730 35264 1735 35320
rect 0 35262 1735 35264
rect 0 35232 800 35262
rect 1669 35259 1735 35262
rect 58157 34914 58223 34917
rect 59200 34914 60000 34944
rect 58157 34912 60000 34914
rect 58157 34856 58162 34912
rect 58218 34856 60000 34912
rect 58157 34854 60000 34856
rect 58157 34851 58223 34854
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 59200 34824 60000 34854
rect 50290 34783 50606 34784
rect 0 34642 800 34672
rect 1669 34642 1735 34645
rect 0 34640 1735 34642
rect 0 34584 1674 34640
rect 1730 34584 1735 34640
rect 0 34582 1735 34584
rect 0 34552 800 34582
rect 1669 34579 1735 34582
rect 24853 34642 24919 34645
rect 25262 34642 25268 34644
rect 24853 34640 25268 34642
rect 24853 34584 24858 34640
rect 24914 34584 25268 34640
rect 24853 34582 25268 34584
rect 24853 34579 24919 34582
rect 25262 34580 25268 34582
rect 25332 34580 25338 34644
rect 57881 34370 57947 34373
rect 59200 34370 60000 34400
rect 57881 34368 60000 34370
rect 57881 34312 57886 34368
rect 57942 34312 60000 34368
rect 57881 34310 60000 34312
rect 57881 34307 57947 34310
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 59200 34280 60000 34310
rect 34930 34239 35246 34240
rect 21541 34098 21607 34101
rect 22737 34098 22803 34101
rect 21541 34096 22803 34098
rect 21541 34040 21546 34096
rect 21602 34040 22742 34096
rect 22798 34040 22803 34096
rect 21541 34038 22803 34040
rect 21541 34035 21607 34038
rect 22737 34035 22803 34038
rect 0 33962 800 33992
rect 1669 33962 1735 33965
rect 0 33960 1735 33962
rect 0 33904 1674 33960
rect 1730 33904 1735 33960
rect 0 33902 1735 33904
rect 0 33872 800 33902
rect 1669 33899 1735 33902
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 59200 33736 60000 33856
rect 50290 33695 50606 33696
rect 21449 33418 21515 33421
rect 25998 33418 26004 33420
rect 21449 33416 26004 33418
rect 21449 33360 21454 33416
rect 21510 33360 26004 33416
rect 21449 33358 26004 33360
rect 21449 33355 21515 33358
rect 25998 33356 26004 33358
rect 26068 33356 26074 33420
rect 0 33282 800 33312
rect 1669 33282 1735 33285
rect 0 33280 1735 33282
rect 0 33224 1674 33280
rect 1730 33224 1735 33280
rect 0 33222 1735 33224
rect 0 33192 800 33222
rect 1669 33219 1735 33222
rect 58157 33282 58223 33285
rect 59200 33282 60000 33312
rect 58157 33280 60000 33282
rect 58157 33224 58162 33280
rect 58218 33224 60000 33280
rect 58157 33222 60000 33224
rect 58157 33219 58223 33222
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 59200 33192 60000 33222
rect 34930 33151 35246 33152
rect 57053 32738 57119 32741
rect 59200 32738 60000 32768
rect 57053 32736 60000 32738
rect 57053 32680 57058 32736
rect 57114 32680 60000 32736
rect 57053 32678 60000 32680
rect 57053 32675 57119 32678
rect 19570 32672 19886 32673
rect 0 32602 800 32632
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 59200 32648 60000 32678
rect 50290 32607 50606 32608
rect 1669 32602 1735 32605
rect 0 32600 1735 32602
rect 0 32544 1674 32600
rect 1730 32544 1735 32600
rect 0 32542 1735 32544
rect 0 32512 800 32542
rect 1669 32539 1735 32542
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 59200 32104 60000 32224
rect 34930 32063 35246 32064
rect 0 31922 800 31952
rect 1669 31922 1735 31925
rect 0 31920 1735 31922
rect 0 31864 1674 31920
rect 1730 31864 1735 31920
rect 0 31862 1735 31864
rect 0 31832 800 31862
rect 1669 31859 1735 31862
rect 58157 31650 58223 31653
rect 59200 31650 60000 31680
rect 58157 31648 60000 31650
rect 58157 31592 58162 31648
rect 58218 31592 60000 31648
rect 58157 31590 60000 31592
rect 58157 31587 58223 31590
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 59200 31560 60000 31590
rect 50290 31519 50606 31520
rect 0 31242 800 31272
rect 1669 31242 1735 31245
rect 0 31240 1735 31242
rect 0 31184 1674 31240
rect 1730 31184 1735 31240
rect 0 31182 1735 31184
rect 0 31152 800 31182
rect 1669 31179 1735 31182
rect 58065 31106 58131 31109
rect 59200 31106 60000 31136
rect 58065 31104 60000 31106
rect 58065 31048 58070 31104
rect 58126 31048 60000 31104
rect 58065 31046 60000 31048
rect 58065 31043 58131 31046
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 59200 31016 60000 31046
rect 34930 30975 35246 30976
rect 0 30562 800 30592
rect 1669 30562 1735 30565
rect 0 30560 1735 30562
rect 0 30504 1674 30560
rect 1730 30504 1735 30560
rect 0 30502 1735 30504
rect 0 30472 800 30502
rect 1669 30499 1735 30502
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 59200 30472 60000 30592
rect 50290 30431 50606 30432
rect 58157 30018 58223 30021
rect 59200 30018 60000 30048
rect 58157 30016 60000 30018
rect 58157 29960 58162 30016
rect 58218 29960 60000 30016
rect 58157 29958 60000 29960
rect 58157 29955 58223 29958
rect 4210 29952 4526 29953
rect 0 29882 800 29912
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 59200 29928 60000 29958
rect 34930 29887 35246 29888
rect 1761 29882 1827 29885
rect 0 29880 1827 29882
rect 0 29824 1766 29880
rect 1822 29824 1827 29880
rect 0 29822 1827 29824
rect 0 29792 800 29822
rect 1761 29819 1827 29822
rect 24853 29610 24919 29613
rect 45318 29610 45324 29612
rect 24853 29608 45324 29610
rect 24853 29552 24858 29608
rect 24914 29552 45324 29608
rect 24853 29550 45324 29552
rect 24853 29547 24919 29550
rect 45318 29548 45324 29550
rect 45388 29548 45394 29612
rect 57053 29474 57119 29477
rect 59200 29474 60000 29504
rect 57053 29472 60000 29474
rect 57053 29416 57058 29472
rect 57114 29416 60000 29472
rect 57053 29414 60000 29416
rect 57053 29411 57119 29414
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 59200 29384 60000 29414
rect 50290 29343 50606 29344
rect 0 29202 800 29232
rect 1853 29202 1919 29205
rect 0 29200 1919 29202
rect 0 29144 1858 29200
rect 1914 29144 1919 29200
rect 0 29142 1919 29144
rect 0 29112 800 29142
rect 1853 29139 1919 29142
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 59200 28840 60000 28960
rect 34930 28799 35246 28800
rect 0 28522 800 28552
rect 1853 28522 1919 28525
rect 0 28520 1919 28522
rect 0 28464 1858 28520
rect 1914 28464 1919 28520
rect 0 28462 1919 28464
rect 0 28432 800 28462
rect 1853 28459 1919 28462
rect 58157 28386 58223 28389
rect 59200 28386 60000 28416
rect 58157 28384 60000 28386
rect 58157 28328 58162 28384
rect 58218 28328 60000 28384
rect 58157 28326 60000 28328
rect 58157 28323 58223 28326
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 59200 28296 60000 28326
rect 50290 28255 50606 28256
rect 0 27842 800 27872
rect 1761 27842 1827 27845
rect 0 27840 1827 27842
rect 0 27784 1766 27840
rect 1822 27784 1827 27840
rect 0 27782 1827 27784
rect 0 27752 800 27782
rect 1761 27779 1827 27782
rect 57973 27842 58039 27845
rect 59200 27842 60000 27872
rect 57973 27840 60000 27842
rect 57973 27784 57978 27840
rect 58034 27784 60000 27840
rect 57973 27782 60000 27784
rect 57973 27779 58039 27782
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 59200 27752 60000 27782
rect 34930 27711 35246 27712
rect 28993 27570 29059 27573
rect 32438 27570 32444 27572
rect 28993 27568 32444 27570
rect 28993 27512 28998 27568
rect 29054 27512 32444 27568
rect 28993 27510 32444 27512
rect 28993 27507 29059 27510
rect 32438 27508 32444 27510
rect 32508 27508 32514 27572
rect 19570 27232 19886 27233
rect 0 27162 800 27192
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 59200 27208 60000 27328
rect 50290 27167 50606 27168
rect 1853 27162 1919 27165
rect 0 27160 1919 27162
rect 0 27104 1858 27160
rect 1914 27104 1919 27160
rect 0 27102 1919 27104
rect 0 27072 800 27102
rect 1853 27099 1919 27102
rect 58157 26754 58223 26757
rect 59200 26754 60000 26784
rect 58157 26752 60000 26754
rect 58157 26696 58162 26752
rect 58218 26696 60000 26752
rect 58157 26694 60000 26696
rect 58157 26691 58223 26694
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 59200 26664 60000 26694
rect 34930 26623 35246 26624
rect 0 26482 800 26512
rect 1761 26482 1827 26485
rect 0 26480 1827 26482
rect 0 26424 1766 26480
rect 1822 26424 1827 26480
rect 0 26422 1827 26424
rect 0 26392 800 26422
rect 1761 26419 1827 26422
rect 58065 26210 58131 26213
rect 59200 26210 60000 26240
rect 58065 26208 60000 26210
rect 58065 26152 58070 26208
rect 58126 26152 60000 26208
rect 58065 26150 60000 26152
rect 58065 26147 58131 26150
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 59200 26120 60000 26150
rect 50290 26079 50606 26080
rect 0 25802 800 25832
rect 1761 25802 1827 25805
rect 0 25800 1827 25802
rect 0 25744 1766 25800
rect 1822 25744 1827 25800
rect 0 25742 1827 25744
rect 0 25712 800 25742
rect 1761 25739 1827 25742
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 59200 25576 60000 25696
rect 34930 25535 35246 25536
rect 22553 25532 22619 25533
rect 22502 25530 22508 25532
rect 22462 25470 22508 25530
rect 22572 25528 22619 25532
rect 22614 25472 22619 25528
rect 22502 25468 22508 25470
rect 22572 25468 22619 25472
rect 22553 25467 22619 25468
rect 17534 25196 17540 25260
rect 17604 25258 17610 25260
rect 20713 25258 20779 25261
rect 17604 25256 20779 25258
rect 17604 25200 20718 25256
rect 20774 25200 20779 25256
rect 17604 25198 20779 25200
rect 17604 25196 17610 25198
rect 20713 25195 20779 25198
rect 0 25122 800 25152
rect 1853 25122 1919 25125
rect 0 25120 1919 25122
rect 0 25064 1858 25120
rect 1914 25064 1919 25120
rect 0 25062 1919 25064
rect 0 25032 800 25062
rect 1853 25059 1919 25062
rect 58157 25122 58223 25125
rect 59200 25122 60000 25152
rect 58157 25120 60000 25122
rect 58157 25064 58162 25120
rect 58218 25064 60000 25120
rect 58157 25062 60000 25064
rect 58157 25059 58223 25062
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 59200 25032 60000 25062
rect 50290 24991 50606 24992
rect 58065 24578 58131 24581
rect 59200 24578 60000 24608
rect 58065 24576 60000 24578
rect 58065 24520 58070 24576
rect 58126 24520 60000 24576
rect 58065 24518 60000 24520
rect 58065 24515 58131 24518
rect 4210 24512 4526 24513
rect 0 24442 800 24472
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 59200 24488 60000 24518
rect 34930 24447 35246 24448
rect 1761 24442 1827 24445
rect 0 24440 1827 24442
rect 0 24384 1766 24440
rect 1822 24384 1827 24440
rect 0 24382 1827 24384
rect 0 24352 800 24382
rect 1761 24379 1827 24382
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 59200 23944 60000 24064
rect 50290 23903 50606 23904
rect 0 23762 800 23792
rect 1853 23762 1919 23765
rect 0 23760 1919 23762
rect 0 23704 1858 23760
rect 1914 23704 1919 23760
rect 0 23702 1919 23704
rect 0 23672 800 23702
rect 1853 23699 1919 23702
rect 58157 23490 58223 23493
rect 59200 23490 60000 23520
rect 58157 23488 60000 23490
rect 58157 23432 58162 23488
rect 58218 23432 60000 23488
rect 58157 23430 60000 23432
rect 58157 23427 58223 23430
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 59200 23400 60000 23430
rect 34930 23359 35246 23360
rect 0 23082 800 23112
rect 1853 23082 1919 23085
rect 0 23080 1919 23082
rect 0 23024 1858 23080
rect 1914 23024 1919 23080
rect 0 23022 1919 23024
rect 0 22992 800 23022
rect 1853 23019 1919 23022
rect 58157 22946 58223 22949
rect 59200 22946 60000 22976
rect 58157 22944 60000 22946
rect 58157 22888 58162 22944
rect 58218 22888 60000 22944
rect 58157 22886 60000 22888
rect 58157 22883 58223 22886
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 59200 22856 60000 22886
rect 50290 22815 50606 22816
rect 0 22402 800 22432
rect 1761 22402 1827 22405
rect 0 22400 1827 22402
rect 0 22344 1766 22400
rect 1822 22344 1827 22400
rect 0 22342 1827 22344
rect 0 22312 800 22342
rect 1761 22339 1827 22342
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 59200 22312 60000 22432
rect 34930 22271 35246 22272
rect 58157 21858 58223 21861
rect 59200 21858 60000 21888
rect 58157 21856 60000 21858
rect 58157 21800 58162 21856
rect 58218 21800 60000 21856
rect 58157 21798 60000 21800
rect 58157 21795 58223 21798
rect 19570 21792 19886 21793
rect 0 21722 800 21752
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 59200 21768 60000 21798
rect 50290 21727 50606 21728
rect 1853 21722 1919 21725
rect 0 21720 1919 21722
rect 0 21664 1858 21720
rect 1914 21664 1919 21720
rect 0 21662 1919 21664
rect 0 21632 800 21662
rect 1853 21659 1919 21662
rect 11053 21314 11119 21317
rect 22553 21314 22619 21317
rect 11053 21312 22619 21314
rect 11053 21256 11058 21312
rect 11114 21256 22558 21312
rect 22614 21256 22619 21312
rect 11053 21254 22619 21256
rect 11053 21251 11119 21254
rect 22553 21251 22619 21254
rect 58065 21314 58131 21317
rect 59200 21314 60000 21344
rect 58065 21312 60000 21314
rect 58065 21256 58070 21312
rect 58126 21256 60000 21312
rect 58065 21254 60000 21256
rect 58065 21251 58131 21254
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 59200 21224 60000 21254
rect 34930 21183 35246 21184
rect 0 21042 800 21072
rect 1761 21042 1827 21045
rect 0 21040 1827 21042
rect 0 20984 1766 21040
rect 1822 20984 1827 21040
rect 0 20982 1827 20984
rect 0 20952 800 20982
rect 1761 20979 1827 20982
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 59200 20680 60000 20800
rect 50290 20639 50606 20640
rect 18505 20498 18571 20501
rect 25129 20498 25195 20501
rect 25957 20498 26023 20501
rect 18505 20496 26023 20498
rect 18505 20440 18510 20496
rect 18566 20440 25134 20496
rect 25190 20440 25962 20496
rect 26018 20440 26023 20496
rect 18505 20438 26023 20440
rect 18505 20435 18571 20438
rect 25129 20435 25195 20438
rect 25957 20435 26023 20438
rect 0 20362 800 20392
rect 1761 20362 1827 20365
rect 0 20360 1827 20362
rect 0 20304 1766 20360
rect 1822 20304 1827 20360
rect 0 20302 1827 20304
rect 0 20272 800 20302
rect 1761 20299 1827 20302
rect 58157 20226 58223 20229
rect 59200 20226 60000 20256
rect 58157 20224 60000 20226
rect 58157 20168 58162 20224
rect 58218 20168 60000 20224
rect 58157 20166 60000 20168
rect 58157 20163 58223 20166
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 59200 20136 60000 20166
rect 34930 20095 35246 20096
rect 49969 20090 50035 20093
rect 51625 20090 51691 20093
rect 49969 20088 51691 20090
rect 49969 20032 49974 20088
rect 50030 20032 51630 20088
rect 51686 20032 51691 20088
rect 49969 20030 51691 20032
rect 49969 20027 50035 20030
rect 51625 20027 51691 20030
rect 35065 19954 35131 19957
rect 57278 19954 57284 19956
rect 35065 19952 57284 19954
rect 35065 19896 35070 19952
rect 35126 19896 57284 19952
rect 35065 19894 57284 19896
rect 35065 19891 35131 19894
rect 57278 19892 57284 19894
rect 57348 19892 57354 19956
rect 22870 19756 22876 19820
rect 22940 19818 22946 19820
rect 24945 19818 25011 19821
rect 22940 19816 25011 19818
rect 22940 19760 24950 19816
rect 25006 19760 25011 19816
rect 22940 19758 25011 19760
rect 22940 19756 22946 19758
rect 24945 19755 25011 19758
rect 50153 19818 50219 19821
rect 50705 19818 50771 19821
rect 50153 19816 50771 19818
rect 50153 19760 50158 19816
rect 50214 19760 50710 19816
rect 50766 19760 50771 19816
rect 50153 19758 50771 19760
rect 50153 19755 50219 19758
rect 50705 19755 50771 19758
rect 0 19682 800 19712
rect 1853 19682 1919 19685
rect 0 19680 1919 19682
rect 0 19624 1858 19680
rect 1914 19624 1919 19680
rect 0 19622 1919 19624
rect 0 19592 800 19622
rect 1853 19619 1919 19622
rect 57973 19682 58039 19685
rect 59200 19682 60000 19712
rect 57973 19680 60000 19682
rect 57973 19624 57978 19680
rect 58034 19624 60000 19680
rect 57973 19622 60000 19624
rect 57973 19619 58039 19622
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 59200 19592 60000 19622
rect 50290 19551 50606 19552
rect 42241 19274 42307 19277
rect 46381 19274 46447 19277
rect 42241 19272 46447 19274
rect 42241 19216 42246 19272
rect 42302 19216 46386 19272
rect 46442 19216 46447 19272
rect 42241 19214 46447 19216
rect 42241 19211 42307 19214
rect 46381 19211 46447 19214
rect 41873 19138 41939 19141
rect 43621 19138 43687 19141
rect 41873 19136 43687 19138
rect 41873 19080 41878 19136
rect 41934 19080 43626 19136
rect 43682 19080 43687 19136
rect 41873 19078 43687 19080
rect 41873 19075 41939 19078
rect 43621 19075 43687 19078
rect 4210 19072 4526 19073
rect 0 19002 800 19032
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 59200 19048 60000 19168
rect 34930 19007 35246 19008
rect 1853 19002 1919 19005
rect 0 19000 1919 19002
rect 0 18944 1858 19000
rect 1914 18944 1919 19000
rect 0 18942 1919 18944
rect 0 18912 800 18942
rect 1853 18939 1919 18942
rect 2405 18866 2471 18869
rect 30782 18866 30788 18868
rect 2405 18864 30788 18866
rect 2405 18808 2410 18864
rect 2466 18808 30788 18864
rect 2405 18806 30788 18808
rect 2405 18803 2471 18806
rect 30782 18804 30788 18806
rect 30852 18804 30858 18868
rect 40033 18866 40099 18869
rect 41137 18866 41203 18869
rect 40033 18864 41203 18866
rect 40033 18808 40038 18864
rect 40094 18808 41142 18864
rect 41198 18808 41203 18864
rect 40033 18806 41203 18808
rect 40033 18803 40099 18806
rect 41137 18803 41203 18806
rect 2405 18730 2471 18733
rect 30966 18730 30972 18732
rect 2405 18728 30972 18730
rect 2405 18672 2410 18728
rect 2466 18672 30972 18728
rect 2405 18670 30972 18672
rect 2405 18667 2471 18670
rect 30966 18668 30972 18670
rect 31036 18668 31042 18732
rect 20897 18594 20963 18597
rect 26509 18594 26575 18597
rect 20897 18592 26575 18594
rect 20897 18536 20902 18592
rect 20958 18536 26514 18592
rect 26570 18536 26575 18592
rect 20897 18534 26575 18536
rect 20897 18531 20963 18534
rect 26509 18531 26575 18534
rect 30649 18594 30715 18597
rect 36997 18594 37063 18597
rect 30649 18592 37063 18594
rect 30649 18536 30654 18592
rect 30710 18536 37002 18592
rect 37058 18536 37063 18592
rect 30649 18534 37063 18536
rect 30649 18531 30715 18534
rect 36997 18531 37063 18534
rect 40953 18594 41019 18597
rect 46565 18594 46631 18597
rect 40953 18592 46631 18594
rect 40953 18536 40958 18592
rect 41014 18536 46570 18592
rect 46626 18536 46631 18592
rect 40953 18534 46631 18536
rect 40953 18531 41019 18534
rect 46565 18531 46631 18534
rect 57237 18594 57303 18597
rect 59200 18594 60000 18624
rect 57237 18592 60000 18594
rect 57237 18536 57242 18592
rect 57298 18536 60000 18592
rect 57237 18534 60000 18536
rect 57237 18531 57303 18534
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 59200 18504 60000 18534
rect 50290 18463 50606 18464
rect 22461 18458 22527 18461
rect 24761 18458 24827 18461
rect 22461 18456 24827 18458
rect 22461 18400 22466 18456
rect 22522 18400 24766 18456
rect 24822 18400 24827 18456
rect 22461 18398 24827 18400
rect 22461 18395 22527 18398
rect 24761 18395 24827 18398
rect 30373 18458 30439 18461
rect 33133 18458 33199 18461
rect 30373 18456 33199 18458
rect 30373 18400 30378 18456
rect 30434 18400 33138 18456
rect 33194 18400 33199 18456
rect 30373 18398 33199 18400
rect 30373 18395 30439 18398
rect 33133 18395 33199 18398
rect 0 18322 800 18352
rect 1853 18322 1919 18325
rect 0 18320 1919 18322
rect 0 18264 1858 18320
rect 1914 18264 1919 18320
rect 0 18262 1919 18264
rect 0 18232 800 18262
rect 1853 18259 1919 18262
rect 21633 18322 21699 18325
rect 23381 18322 23447 18325
rect 21633 18320 23447 18322
rect 21633 18264 21638 18320
rect 21694 18264 23386 18320
rect 23442 18264 23447 18320
rect 21633 18262 23447 18264
rect 21633 18259 21699 18262
rect 23381 18259 23447 18262
rect 42793 18322 42859 18325
rect 46933 18322 46999 18325
rect 42793 18320 46999 18322
rect 42793 18264 42798 18320
rect 42854 18264 46938 18320
rect 46994 18264 46999 18320
rect 42793 18262 46999 18264
rect 42793 18259 42859 18262
rect 46933 18259 46999 18262
rect 28022 17988 28028 18052
rect 28092 18050 28098 18052
rect 31293 18050 31359 18053
rect 28092 18048 31359 18050
rect 28092 17992 31298 18048
rect 31354 17992 31359 18048
rect 28092 17990 31359 17992
rect 28092 17988 28098 17990
rect 31293 17987 31359 17990
rect 31477 18050 31543 18053
rect 31753 18050 31819 18053
rect 31477 18048 31819 18050
rect 31477 17992 31482 18048
rect 31538 17992 31758 18048
rect 31814 17992 31819 18048
rect 31477 17990 31819 17992
rect 31477 17987 31543 17990
rect 31753 17987 31819 17990
rect 57973 18050 58039 18053
rect 59200 18050 60000 18080
rect 57973 18048 60000 18050
rect 57973 17992 57978 18048
rect 58034 17992 60000 18048
rect 57973 17990 60000 17992
rect 57973 17987 58039 17990
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 59200 17960 60000 17990
rect 34930 17919 35246 17920
rect 28758 17852 28764 17916
rect 28828 17914 28834 17916
rect 28901 17914 28967 17917
rect 28828 17912 28967 17914
rect 28828 17856 28906 17912
rect 28962 17856 28967 17912
rect 28828 17854 28967 17856
rect 28828 17852 28834 17854
rect 28901 17851 28967 17854
rect 29545 17914 29611 17917
rect 33777 17914 33843 17917
rect 29545 17912 33843 17914
rect 29545 17856 29550 17912
rect 29606 17856 33782 17912
rect 33838 17856 33843 17912
rect 29545 17854 33843 17856
rect 29545 17851 29611 17854
rect 33777 17851 33843 17854
rect 32397 17780 32463 17781
rect 32397 17778 32444 17780
rect 32352 17776 32444 17778
rect 32352 17720 32402 17776
rect 32352 17718 32444 17720
rect 32397 17716 32444 17718
rect 32508 17716 32514 17780
rect 32397 17715 32463 17716
rect 0 17642 800 17672
rect 1853 17642 1919 17645
rect 0 17640 1919 17642
rect 0 17584 1858 17640
rect 1914 17584 1919 17640
rect 0 17582 1919 17584
rect 0 17552 800 17582
rect 1853 17579 1919 17582
rect 32581 17642 32647 17645
rect 35157 17642 35223 17645
rect 32581 17640 35223 17642
rect 32581 17584 32586 17640
rect 32642 17584 35162 17640
rect 35218 17584 35223 17640
rect 32581 17582 35223 17584
rect 32581 17579 32647 17582
rect 35157 17579 35223 17582
rect 25037 17506 25103 17509
rect 36537 17506 36603 17509
rect 25037 17504 36603 17506
rect 25037 17448 25042 17504
rect 25098 17448 36542 17504
rect 36598 17448 36603 17504
rect 25037 17446 36603 17448
rect 25037 17443 25103 17446
rect 36537 17443 36603 17446
rect 38561 17506 38627 17509
rect 39665 17506 39731 17509
rect 38561 17504 39731 17506
rect 38561 17448 38566 17504
rect 38622 17448 39670 17504
rect 39726 17448 39731 17504
rect 38561 17446 39731 17448
rect 38561 17443 38627 17446
rect 39665 17443 39731 17446
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 59200 17416 60000 17536
rect 50290 17375 50606 17376
rect 28165 17370 28231 17373
rect 22050 17368 28231 17370
rect 22050 17312 28170 17368
rect 28226 17312 28231 17368
rect 22050 17310 28231 17312
rect 2405 17234 2471 17237
rect 22050 17234 22110 17310
rect 28165 17307 28231 17310
rect 30833 17370 30899 17373
rect 34513 17370 34579 17373
rect 30833 17368 34579 17370
rect 30833 17312 30838 17368
rect 30894 17312 34518 17368
rect 34574 17312 34579 17368
rect 30833 17310 34579 17312
rect 30833 17307 30899 17310
rect 34513 17307 34579 17310
rect 38653 17372 38719 17373
rect 38653 17368 38700 17372
rect 38764 17370 38770 17372
rect 38653 17312 38658 17368
rect 38653 17308 38700 17312
rect 38764 17310 38810 17370
rect 38764 17308 38770 17310
rect 38653 17307 38719 17308
rect 2405 17232 22110 17234
rect 2405 17176 2410 17232
rect 2466 17176 22110 17232
rect 2405 17174 22110 17176
rect 24393 17234 24459 17237
rect 25221 17234 25287 17237
rect 25446 17234 25452 17236
rect 24393 17232 25452 17234
rect 24393 17176 24398 17232
rect 24454 17176 25226 17232
rect 25282 17176 25452 17232
rect 24393 17174 25452 17176
rect 2405 17171 2471 17174
rect 24393 17171 24459 17174
rect 25221 17171 25287 17174
rect 25446 17172 25452 17174
rect 25516 17172 25522 17236
rect 29085 17234 29151 17237
rect 33041 17234 33107 17237
rect 29085 17232 33107 17234
rect 29085 17176 29090 17232
rect 29146 17176 33046 17232
rect 33102 17176 33107 17232
rect 29085 17174 33107 17176
rect 29085 17171 29151 17174
rect 33041 17171 33107 17174
rect 38745 17234 38811 17237
rect 41321 17234 41387 17237
rect 38745 17232 41387 17234
rect 38745 17176 38750 17232
rect 38806 17176 41326 17232
rect 41382 17176 41387 17232
rect 38745 17174 41387 17176
rect 38745 17171 38811 17174
rect 41321 17171 41387 17174
rect 51165 17234 51231 17237
rect 54293 17234 54359 17237
rect 51165 17232 54359 17234
rect 51165 17176 51170 17232
rect 51226 17176 54298 17232
rect 54354 17176 54359 17232
rect 51165 17174 54359 17176
rect 51165 17171 51231 17174
rect 54293 17171 54359 17174
rect 28717 17098 28783 17101
rect 38285 17098 38351 17101
rect 28717 17096 38351 17098
rect 28717 17040 28722 17096
rect 28778 17040 38290 17096
rect 38346 17040 38351 17096
rect 28717 17038 38351 17040
rect 28717 17035 28783 17038
rect 38285 17035 38351 17038
rect 38469 17098 38535 17101
rect 39757 17098 39823 17101
rect 38469 17096 39823 17098
rect 38469 17040 38474 17096
rect 38530 17040 39762 17096
rect 39818 17040 39823 17096
rect 38469 17038 39823 17040
rect 38469 17035 38535 17038
rect 39757 17035 39823 17038
rect 53925 17098 53991 17101
rect 55765 17098 55831 17101
rect 53925 17096 55831 17098
rect 53925 17040 53930 17096
rect 53986 17040 55770 17096
rect 55826 17040 55831 17096
rect 53925 17038 55831 17040
rect 53925 17035 53991 17038
rect 55765 17035 55831 17038
rect 0 16962 800 16992
rect 1761 16962 1827 16965
rect 0 16960 1827 16962
rect 0 16904 1766 16960
rect 1822 16904 1827 16960
rect 0 16902 1827 16904
rect 0 16872 800 16902
rect 1761 16899 1827 16902
rect 27521 16962 27587 16965
rect 28942 16962 28948 16964
rect 27521 16960 28948 16962
rect 27521 16904 27526 16960
rect 27582 16904 28948 16960
rect 27521 16902 28948 16904
rect 27521 16899 27587 16902
rect 28942 16900 28948 16902
rect 29012 16900 29018 16964
rect 38377 16962 38443 16965
rect 38837 16962 38903 16965
rect 38377 16960 38903 16962
rect 38377 16904 38382 16960
rect 38438 16904 38842 16960
rect 38898 16904 38903 16960
rect 38377 16902 38903 16904
rect 38377 16899 38443 16902
rect 38837 16899 38903 16902
rect 57329 16962 57395 16965
rect 59200 16962 60000 16992
rect 57329 16960 60000 16962
rect 57329 16904 57334 16960
rect 57390 16904 60000 16960
rect 57329 16902 60000 16904
rect 57329 16899 57395 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 59200 16872 60000 16902
rect 34930 16831 35246 16832
rect 31661 16826 31727 16829
rect 33593 16826 33659 16829
rect 31661 16824 33659 16826
rect 31661 16768 31666 16824
rect 31722 16768 33598 16824
rect 33654 16768 33659 16824
rect 31661 16766 33659 16768
rect 31661 16763 31727 16766
rect 33593 16763 33659 16766
rect 27889 16554 27955 16557
rect 42885 16556 42951 16557
rect 28022 16554 28028 16556
rect 27889 16552 28028 16554
rect 27889 16496 27894 16552
rect 27950 16496 28028 16552
rect 27889 16494 28028 16496
rect 27889 16491 27955 16494
rect 28022 16492 28028 16494
rect 28092 16492 28098 16556
rect 42885 16552 42932 16556
rect 42996 16554 43002 16556
rect 42885 16496 42890 16552
rect 42885 16492 42932 16496
rect 42996 16494 43042 16554
rect 42996 16492 43002 16494
rect 42885 16491 42951 16492
rect 24853 16418 24919 16421
rect 25221 16418 25287 16421
rect 25957 16418 26023 16421
rect 24853 16416 26023 16418
rect 24853 16360 24858 16416
rect 24914 16360 25226 16416
rect 25282 16360 25962 16416
rect 26018 16360 26023 16416
rect 24853 16358 26023 16360
rect 24853 16355 24919 16358
rect 25221 16355 25287 16358
rect 25957 16355 26023 16358
rect 57053 16418 57119 16421
rect 59200 16418 60000 16448
rect 57053 16416 60000 16418
rect 57053 16360 57058 16416
rect 57114 16360 60000 16416
rect 57053 16358 60000 16360
rect 57053 16355 57119 16358
rect 19570 16352 19886 16353
rect 0 16282 800 16312
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 59200 16328 60000 16358
rect 50290 16287 50606 16288
rect 1853 16282 1919 16285
rect 0 16280 1919 16282
rect 0 16224 1858 16280
rect 1914 16224 1919 16280
rect 0 16222 1919 16224
rect 0 16192 800 16222
rect 1853 16219 1919 16222
rect 29494 16220 29500 16284
rect 29564 16282 29570 16284
rect 38694 16282 38700 16284
rect 29564 16222 38700 16282
rect 29564 16220 29570 16222
rect 38694 16220 38700 16222
rect 38764 16282 38770 16284
rect 38837 16282 38903 16285
rect 38764 16280 38903 16282
rect 38764 16224 38842 16280
rect 38898 16224 38903 16280
rect 38764 16222 38903 16224
rect 38764 16220 38770 16222
rect 38837 16219 38903 16222
rect 15377 16146 15443 16149
rect 46565 16146 46631 16149
rect 15377 16144 46631 16146
rect 15377 16088 15382 16144
rect 15438 16088 46570 16144
rect 46626 16088 46631 16144
rect 15377 16086 46631 16088
rect 15377 16083 15443 16086
rect 46565 16083 46631 16086
rect 2405 16010 2471 16013
rect 20713 16010 20779 16013
rect 2405 16008 20779 16010
rect 2405 15952 2410 16008
rect 2466 15952 20718 16008
rect 20774 15952 20779 16008
rect 2405 15950 20779 15952
rect 2405 15947 2471 15950
rect 20713 15947 20779 15950
rect 22461 16010 22527 16013
rect 32397 16010 32463 16013
rect 22461 16008 32463 16010
rect 22461 15952 22466 16008
rect 22522 15952 32402 16008
rect 32458 15952 32463 16008
rect 22461 15950 32463 15952
rect 22461 15947 22527 15950
rect 32397 15947 32463 15950
rect 21541 15874 21607 15877
rect 21909 15874 21975 15877
rect 31845 15874 31911 15877
rect 32581 15874 32647 15877
rect 21541 15872 32647 15874
rect 21541 15816 21546 15872
rect 21602 15816 21914 15872
rect 21970 15816 31850 15872
rect 31906 15816 32586 15872
rect 32642 15816 32647 15872
rect 21541 15814 32647 15816
rect 21541 15811 21607 15814
rect 21909 15811 21975 15814
rect 31845 15811 31911 15814
rect 32581 15811 32647 15814
rect 40953 15874 41019 15877
rect 41086 15874 41092 15876
rect 40953 15872 41092 15874
rect 40953 15816 40958 15872
rect 41014 15816 41092 15872
rect 40953 15814 41092 15816
rect 40953 15811 41019 15814
rect 41086 15812 41092 15814
rect 41156 15812 41162 15876
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 59200 15784 60000 15904
rect 34930 15743 35246 15744
rect 20897 15738 20963 15741
rect 28441 15738 28507 15741
rect 20897 15736 28507 15738
rect 20897 15680 20902 15736
rect 20958 15680 28446 15736
rect 28502 15680 28507 15736
rect 20897 15678 28507 15680
rect 20897 15675 20963 15678
rect 28441 15675 28507 15678
rect 0 15602 800 15632
rect 1761 15602 1827 15605
rect 0 15600 1827 15602
rect 0 15544 1766 15600
rect 1822 15544 1827 15600
rect 0 15542 1827 15544
rect 0 15512 800 15542
rect 1761 15539 1827 15542
rect 25681 15602 25747 15605
rect 40033 15602 40099 15605
rect 41045 15602 41111 15605
rect 25681 15600 41111 15602
rect 25681 15544 25686 15600
rect 25742 15544 40038 15600
rect 40094 15544 41050 15600
rect 41106 15544 41111 15600
rect 25681 15542 41111 15544
rect 25681 15539 25747 15542
rect 40033 15539 40099 15542
rect 41045 15539 41111 15542
rect 23381 15466 23447 15469
rect 25313 15466 25379 15469
rect 23381 15464 25379 15466
rect 23381 15408 23386 15464
rect 23442 15408 25318 15464
rect 25374 15408 25379 15464
rect 23381 15406 25379 15408
rect 23381 15403 23447 15406
rect 25313 15403 25379 15406
rect 28441 15466 28507 15469
rect 57145 15466 57211 15469
rect 28441 15464 57211 15466
rect 28441 15408 28446 15464
rect 28502 15408 57150 15464
rect 57206 15408 57211 15464
rect 28441 15406 57211 15408
rect 28441 15403 28507 15406
rect 57145 15403 57211 15406
rect 26693 15330 26759 15333
rect 30465 15330 30531 15333
rect 26693 15328 30531 15330
rect 26693 15272 26698 15328
rect 26754 15272 30470 15328
rect 30526 15272 30531 15328
rect 26693 15270 30531 15272
rect 26693 15267 26759 15270
rect 30465 15267 30531 15270
rect 58157 15330 58223 15333
rect 59200 15330 60000 15360
rect 58157 15328 60000 15330
rect 58157 15272 58162 15328
rect 58218 15272 60000 15328
rect 58157 15270 60000 15272
rect 58157 15267 58223 15270
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 59200 15240 60000 15270
rect 50290 15199 50606 15200
rect 20437 15194 20503 15197
rect 24669 15194 24735 15197
rect 20437 15192 24735 15194
rect 20437 15136 20442 15192
rect 20498 15136 24674 15192
rect 24730 15136 24735 15192
rect 20437 15134 24735 15136
rect 20437 15131 20503 15134
rect 24669 15131 24735 15134
rect 29821 15058 29887 15061
rect 30465 15058 30531 15061
rect 29821 15056 30531 15058
rect 29821 15000 29826 15056
rect 29882 15000 30470 15056
rect 30526 15000 30531 15056
rect 29821 14998 30531 15000
rect 29821 14995 29887 14998
rect 30465 14995 30531 14998
rect 0 14922 800 14952
rect 1761 14922 1827 14925
rect 0 14920 1827 14922
rect 0 14864 1766 14920
rect 1822 14864 1827 14920
rect 0 14862 1827 14864
rect 0 14832 800 14862
rect 1761 14859 1827 14862
rect 57973 14786 58039 14789
rect 59200 14786 60000 14816
rect 57973 14784 60000 14786
rect 57973 14728 57978 14784
rect 58034 14728 60000 14784
rect 57973 14726 60000 14728
rect 57973 14723 58039 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 59200 14696 60000 14726
rect 34930 14655 35246 14656
rect 20713 14650 20779 14653
rect 30598 14650 30604 14652
rect 20713 14648 30604 14650
rect 20713 14592 20718 14648
rect 20774 14592 30604 14648
rect 20713 14590 30604 14592
rect 20713 14587 20779 14590
rect 30598 14588 30604 14590
rect 30668 14588 30674 14652
rect 2405 14514 2471 14517
rect 31886 14514 31892 14516
rect 2405 14512 31892 14514
rect 2405 14456 2410 14512
rect 2466 14456 31892 14512
rect 2405 14454 31892 14456
rect 2405 14451 2471 14454
rect 31886 14452 31892 14454
rect 31956 14452 31962 14516
rect 32857 14514 32923 14517
rect 42517 14514 42583 14517
rect 32857 14512 42583 14514
rect 32857 14456 32862 14512
rect 32918 14456 42522 14512
rect 42578 14456 42583 14512
rect 32857 14454 42583 14456
rect 32857 14451 32923 14454
rect 42517 14451 42583 14454
rect 19609 14378 19675 14381
rect 21449 14378 21515 14381
rect 19609 14376 21515 14378
rect 19609 14320 19614 14376
rect 19670 14320 21454 14376
rect 21510 14320 21515 14376
rect 19609 14318 21515 14320
rect 19609 14315 19675 14318
rect 21449 14315 21515 14318
rect 32029 14378 32095 14381
rect 35249 14378 35315 14381
rect 32029 14376 35315 14378
rect 32029 14320 32034 14376
rect 32090 14320 35254 14376
rect 35310 14320 35315 14376
rect 32029 14318 35315 14320
rect 32029 14315 32095 14318
rect 35249 14315 35315 14318
rect 0 14242 800 14272
rect 1853 14242 1919 14245
rect 0 14240 1919 14242
rect 0 14184 1858 14240
rect 1914 14184 1919 14240
rect 0 14182 1919 14184
rect 0 14152 800 14182
rect 1853 14179 1919 14182
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 59200 14152 60000 14272
rect 50290 14111 50606 14112
rect 26141 13970 26207 13973
rect 28993 13970 29059 13973
rect 26141 13968 29059 13970
rect 26141 13912 26146 13968
rect 26202 13912 28998 13968
rect 29054 13912 29059 13968
rect 26141 13910 29059 13912
rect 26141 13907 26207 13910
rect 28993 13907 29059 13910
rect 18689 13834 18755 13837
rect 22185 13834 22251 13837
rect 18689 13832 22251 13834
rect 18689 13776 18694 13832
rect 18750 13776 22190 13832
rect 22246 13776 22251 13832
rect 18689 13774 22251 13776
rect 18689 13771 18755 13774
rect 22185 13771 22251 13774
rect 24393 13834 24459 13837
rect 58065 13834 58131 13837
rect 24393 13832 58131 13834
rect 24393 13776 24398 13832
rect 24454 13776 58070 13832
rect 58126 13776 58131 13832
rect 24393 13774 58131 13776
rect 24393 13771 24459 13774
rect 58065 13771 58131 13774
rect 58157 13698 58223 13701
rect 59200 13698 60000 13728
rect 58157 13696 60000 13698
rect 58157 13640 58162 13696
rect 58218 13640 60000 13696
rect 58157 13638 60000 13640
rect 58157 13635 58223 13638
rect 4210 13632 4526 13633
rect 0 13562 800 13592
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 59200 13608 60000 13638
rect 34930 13567 35246 13568
rect 1761 13562 1827 13565
rect 0 13560 1827 13562
rect 0 13504 1766 13560
rect 1822 13504 1827 13560
rect 0 13502 1827 13504
rect 0 13472 800 13502
rect 1761 13499 1827 13502
rect 15101 13426 15167 13429
rect 18413 13426 18479 13429
rect 15101 13424 18479 13426
rect 15101 13368 15106 13424
rect 15162 13368 18418 13424
rect 18474 13368 18479 13424
rect 15101 13366 18479 13368
rect 15101 13363 15167 13366
rect 18413 13363 18479 13366
rect 31569 13426 31635 13429
rect 38561 13426 38627 13429
rect 31569 13424 38627 13426
rect 31569 13368 31574 13424
rect 31630 13368 38566 13424
rect 38622 13368 38627 13424
rect 31569 13366 38627 13368
rect 31569 13363 31635 13366
rect 38561 13363 38627 13366
rect 6913 13290 6979 13293
rect 32121 13290 32187 13293
rect 6913 13288 32187 13290
rect 6913 13232 6918 13288
rect 6974 13232 32126 13288
rect 32182 13232 32187 13288
rect 6913 13230 32187 13232
rect 6913 13227 6979 13230
rect 32121 13227 32187 13230
rect 36261 13290 36327 13293
rect 37273 13290 37339 13293
rect 36261 13288 37339 13290
rect 36261 13232 36266 13288
rect 36322 13232 37278 13288
rect 37334 13232 37339 13288
rect 36261 13230 37339 13232
rect 36261 13227 36327 13230
rect 37273 13227 37339 13230
rect 23841 13154 23907 13157
rect 27613 13154 27679 13157
rect 23841 13152 27679 13154
rect 23841 13096 23846 13152
rect 23902 13096 27618 13152
rect 27674 13096 27679 13152
rect 23841 13094 27679 13096
rect 23841 13091 23907 13094
rect 27613 13091 27679 13094
rect 32673 13154 32739 13157
rect 37457 13154 37523 13157
rect 32673 13152 37523 13154
rect 32673 13096 32678 13152
rect 32734 13096 37462 13152
rect 37518 13096 37523 13152
rect 32673 13094 37523 13096
rect 32673 13091 32739 13094
rect 37457 13091 37523 13094
rect 56961 13154 57027 13157
rect 59200 13154 60000 13184
rect 56961 13152 60000 13154
rect 56961 13096 56966 13152
rect 57022 13096 60000 13152
rect 56961 13094 60000 13096
rect 56961 13091 57027 13094
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 59200 13064 60000 13094
rect 50290 13023 50606 13024
rect 11881 13018 11947 13021
rect 17953 13018 18019 13021
rect 11881 13016 18019 13018
rect 11881 12960 11886 13016
rect 11942 12960 17958 13016
rect 18014 12960 18019 13016
rect 11881 12958 18019 12960
rect 11881 12955 11947 12958
rect 17953 12955 18019 12958
rect 28942 12956 28948 13020
rect 29012 13018 29018 13020
rect 45134 13018 45140 13020
rect 29012 12958 45140 13018
rect 29012 12956 29018 12958
rect 45134 12956 45140 12958
rect 45204 12956 45210 13020
rect 0 12882 800 12912
rect 1853 12882 1919 12885
rect 0 12880 1919 12882
rect 0 12824 1858 12880
rect 1914 12824 1919 12880
rect 0 12822 1919 12824
rect 0 12792 800 12822
rect 1853 12819 1919 12822
rect 31385 12882 31451 12885
rect 36445 12882 36511 12885
rect 31385 12880 36511 12882
rect 31385 12824 31390 12880
rect 31446 12824 36450 12880
rect 36506 12824 36511 12880
rect 31385 12822 36511 12824
rect 31385 12819 31451 12822
rect 36445 12819 36511 12822
rect 34237 12746 34303 12749
rect 39021 12746 39087 12749
rect 34237 12744 39087 12746
rect 34237 12688 34242 12744
rect 34298 12688 39026 12744
rect 39082 12688 39087 12744
rect 34237 12686 39087 12688
rect 34237 12683 34303 12686
rect 39021 12683 39087 12686
rect 19517 12610 19583 12613
rect 20161 12610 20227 12613
rect 19517 12608 20227 12610
rect 19517 12552 19522 12608
rect 19578 12552 20166 12608
rect 20222 12552 20227 12608
rect 19517 12550 20227 12552
rect 19517 12547 19583 12550
rect 20161 12547 20227 12550
rect 39062 12548 39068 12612
rect 39132 12610 39138 12612
rect 39205 12610 39271 12613
rect 39132 12608 39271 12610
rect 39132 12552 39210 12608
rect 39266 12552 39271 12608
rect 39132 12550 39271 12552
rect 39132 12548 39138 12550
rect 39205 12547 39271 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 59200 12520 60000 12640
rect 34930 12479 35246 12480
rect 21817 12474 21883 12477
rect 28165 12474 28231 12477
rect 21817 12472 28231 12474
rect 21817 12416 21822 12472
rect 21878 12416 28170 12472
rect 28226 12416 28231 12472
rect 21817 12414 28231 12416
rect 21817 12411 21883 12414
rect 28165 12411 28231 12414
rect 40718 12412 40724 12476
rect 40788 12474 40794 12476
rect 42149 12474 42215 12477
rect 40788 12472 42215 12474
rect 40788 12416 42154 12472
rect 42210 12416 42215 12472
rect 40788 12414 42215 12416
rect 40788 12412 40794 12414
rect 42149 12411 42215 12414
rect 26969 12338 27035 12341
rect 27337 12338 27403 12341
rect 26969 12336 27403 12338
rect 26969 12280 26974 12336
rect 27030 12280 27342 12336
rect 27398 12280 27403 12336
rect 26969 12278 27403 12280
rect 26969 12275 27035 12278
rect 27337 12275 27403 12278
rect 0 12202 800 12232
rect 1853 12202 1919 12205
rect 0 12200 1919 12202
rect 0 12144 1858 12200
rect 1914 12144 1919 12200
rect 0 12142 1919 12144
rect 0 12112 800 12142
rect 1853 12139 1919 12142
rect 12065 12202 12131 12205
rect 21265 12202 21331 12205
rect 12065 12200 21331 12202
rect 12065 12144 12070 12200
rect 12126 12144 21270 12200
rect 21326 12144 21331 12200
rect 12065 12142 21331 12144
rect 12065 12139 12131 12142
rect 21265 12139 21331 12142
rect 35341 12202 35407 12205
rect 36077 12202 36143 12205
rect 35341 12200 36143 12202
rect 35341 12144 35346 12200
rect 35402 12144 36082 12200
rect 36138 12144 36143 12200
rect 35341 12142 36143 12144
rect 35341 12139 35407 12142
rect 36077 12139 36143 12142
rect 24025 12066 24091 12069
rect 22050 12064 24091 12066
rect 22050 12008 24030 12064
rect 24086 12008 24091 12064
rect 22050 12006 24091 12008
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 19977 11930 20043 11933
rect 22050 11930 22110 12006
rect 24025 12003 24091 12006
rect 24301 12066 24367 12069
rect 28349 12066 28415 12069
rect 24301 12064 28415 12066
rect 24301 12008 24306 12064
rect 24362 12008 28354 12064
rect 28410 12008 28415 12064
rect 24301 12006 28415 12008
rect 24301 12003 24367 12006
rect 28349 12003 28415 12006
rect 32305 12066 32371 12069
rect 35801 12066 35867 12069
rect 38101 12066 38167 12069
rect 32305 12064 38167 12066
rect 32305 12008 32310 12064
rect 32366 12008 35806 12064
rect 35862 12008 38106 12064
rect 38162 12008 38167 12064
rect 32305 12006 38167 12008
rect 32305 12003 32371 12006
rect 35801 12003 35867 12006
rect 38101 12003 38167 12006
rect 58157 12066 58223 12069
rect 59200 12066 60000 12096
rect 58157 12064 60000 12066
rect 58157 12008 58162 12064
rect 58218 12008 60000 12064
rect 58157 12006 60000 12008
rect 58157 12003 58223 12006
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 59200 11976 60000 12006
rect 50290 11935 50606 11936
rect 19977 11928 22110 11930
rect 19977 11872 19982 11928
rect 20038 11872 22110 11928
rect 19977 11870 22110 11872
rect 23289 11930 23355 11933
rect 36721 11930 36787 11933
rect 23289 11928 36787 11930
rect 23289 11872 23294 11928
rect 23350 11872 36726 11928
rect 36782 11872 36787 11928
rect 23289 11870 36787 11872
rect 19977 11867 20043 11870
rect 23289 11867 23355 11870
rect 36721 11867 36787 11870
rect 11881 11794 11947 11797
rect 16113 11794 16179 11797
rect 11881 11792 16179 11794
rect 11881 11736 11886 11792
rect 11942 11736 16118 11792
rect 16174 11736 16179 11792
rect 11881 11734 16179 11736
rect 11881 11731 11947 11734
rect 16113 11731 16179 11734
rect 17033 11794 17099 11797
rect 27337 11794 27403 11797
rect 17033 11792 27403 11794
rect 17033 11736 17038 11792
rect 17094 11736 27342 11792
rect 27398 11736 27403 11792
rect 17033 11734 27403 11736
rect 17033 11731 17099 11734
rect 27337 11731 27403 11734
rect 40125 11794 40191 11797
rect 41689 11794 41755 11797
rect 40125 11792 41755 11794
rect 40125 11736 40130 11792
rect 40186 11736 41694 11792
rect 41750 11736 41755 11792
rect 40125 11734 41755 11736
rect 40125 11731 40191 11734
rect 41689 11731 41755 11734
rect 14733 11658 14799 11661
rect 15285 11658 15351 11661
rect 16665 11658 16731 11661
rect 19241 11658 19307 11661
rect 14733 11656 19307 11658
rect 14733 11600 14738 11656
rect 14794 11600 15290 11656
rect 15346 11600 16670 11656
rect 16726 11600 19246 11656
rect 19302 11600 19307 11656
rect 14733 11598 19307 11600
rect 14733 11595 14799 11598
rect 15285 11595 15351 11598
rect 16665 11595 16731 11598
rect 19241 11595 19307 11598
rect 19793 11658 19859 11661
rect 22185 11658 22251 11661
rect 19793 11656 22251 11658
rect 19793 11600 19798 11656
rect 19854 11600 22190 11656
rect 22246 11600 22251 11656
rect 19793 11598 22251 11600
rect 19793 11595 19859 11598
rect 22185 11595 22251 11598
rect 23013 11658 23079 11661
rect 24485 11658 24551 11661
rect 23013 11656 24551 11658
rect 23013 11600 23018 11656
rect 23074 11600 24490 11656
rect 24546 11600 24551 11656
rect 23013 11598 24551 11600
rect 23013 11595 23079 11598
rect 24485 11595 24551 11598
rect 0 11522 800 11552
rect 1761 11522 1827 11525
rect 0 11520 1827 11522
rect 0 11464 1766 11520
rect 1822 11464 1827 11520
rect 0 11462 1827 11464
rect 0 11432 800 11462
rect 1761 11459 1827 11462
rect 14825 11522 14891 11525
rect 17401 11522 17467 11525
rect 14825 11520 17467 11522
rect 14825 11464 14830 11520
rect 14886 11464 17406 11520
rect 17462 11464 17467 11520
rect 14825 11462 17467 11464
rect 14825 11459 14891 11462
rect 17401 11459 17467 11462
rect 20069 11522 20135 11525
rect 26049 11522 26115 11525
rect 20069 11520 26115 11522
rect 20069 11464 20074 11520
rect 20130 11464 26054 11520
rect 26110 11464 26115 11520
rect 20069 11462 26115 11464
rect 20069 11459 20135 11462
rect 26049 11459 26115 11462
rect 57145 11522 57211 11525
rect 59200 11522 60000 11552
rect 57145 11520 60000 11522
rect 57145 11464 57150 11520
rect 57206 11464 60000 11520
rect 57145 11462 60000 11464
rect 57145 11459 57211 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 59200 11432 60000 11462
rect 34930 11391 35246 11392
rect 19701 11386 19767 11389
rect 21449 11386 21515 11389
rect 19701 11384 21515 11386
rect 19701 11328 19706 11384
rect 19762 11328 21454 11384
rect 21510 11328 21515 11384
rect 19701 11326 21515 11328
rect 19701 11323 19767 11326
rect 21449 11323 21515 11326
rect 40033 11386 40099 11389
rect 42425 11386 42491 11389
rect 40033 11384 42491 11386
rect 40033 11328 40038 11384
rect 40094 11328 42430 11384
rect 42486 11328 42491 11384
rect 40033 11326 42491 11328
rect 40033 11323 40099 11326
rect 42425 11323 42491 11326
rect 14825 11250 14891 11253
rect 17861 11250 17927 11253
rect 14825 11248 17927 11250
rect 14825 11192 14830 11248
rect 14886 11192 17866 11248
rect 17922 11192 17927 11248
rect 14825 11190 17927 11192
rect 14825 11187 14891 11190
rect 17861 11187 17927 11190
rect 24393 11250 24459 11253
rect 29177 11250 29243 11253
rect 24393 11248 29243 11250
rect 24393 11192 24398 11248
rect 24454 11192 29182 11248
rect 29238 11192 29243 11248
rect 24393 11190 29243 11192
rect 24393 11187 24459 11190
rect 29177 11187 29243 11190
rect 31753 11250 31819 11253
rect 41413 11250 41479 11253
rect 31753 11248 41479 11250
rect 31753 11192 31758 11248
rect 31814 11192 41418 11248
rect 41474 11192 41479 11248
rect 31753 11190 41479 11192
rect 31753 11187 31819 11190
rect 41413 11187 41479 11190
rect 16849 11114 16915 11117
rect 21725 11114 21791 11117
rect 23933 11114 23999 11117
rect 16849 11112 23999 11114
rect 16849 11056 16854 11112
rect 16910 11056 21730 11112
rect 21786 11056 23938 11112
rect 23994 11056 23999 11112
rect 16849 11054 23999 11056
rect 16849 11051 16915 11054
rect 21725 11051 21791 11054
rect 23933 11051 23999 11054
rect 24485 11114 24551 11117
rect 27337 11114 27403 11117
rect 27797 11114 27863 11117
rect 24485 11112 27863 11114
rect 24485 11056 24490 11112
rect 24546 11056 27342 11112
rect 27398 11056 27802 11112
rect 27858 11056 27863 11112
rect 24485 11054 27863 11056
rect 24485 11051 24551 11054
rect 27337 11051 27403 11054
rect 27797 11051 27863 11054
rect 28165 11114 28231 11117
rect 31385 11114 31451 11117
rect 28165 11112 31451 11114
rect 28165 11056 28170 11112
rect 28226 11056 31390 11112
rect 31446 11056 31451 11112
rect 28165 11054 31451 11056
rect 28165 11051 28231 11054
rect 31385 11051 31451 11054
rect 37825 11114 37891 11117
rect 39246 11114 39252 11116
rect 37825 11112 39252 11114
rect 37825 11056 37830 11112
rect 37886 11056 39252 11112
rect 37825 11054 39252 11056
rect 37825 11051 37891 11054
rect 39246 11052 39252 11054
rect 39316 11052 39322 11116
rect 23657 10978 23723 10981
rect 24669 10978 24735 10981
rect 23657 10976 24735 10978
rect 23657 10920 23662 10976
rect 23718 10920 24674 10976
rect 24730 10920 24735 10976
rect 23657 10918 24735 10920
rect 23657 10915 23723 10918
rect 24669 10915 24735 10918
rect 30005 10980 30071 10981
rect 30005 10976 30052 10980
rect 30116 10978 30122 10980
rect 30005 10920 30010 10976
rect 30005 10916 30052 10920
rect 30116 10918 30162 10978
rect 30116 10916 30122 10918
rect 30005 10915 30071 10916
rect 19570 10912 19886 10913
rect 0 10842 800 10872
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 59200 10888 60000 11008
rect 50290 10847 50606 10848
rect 1853 10842 1919 10845
rect 0 10840 1919 10842
rect 0 10784 1858 10840
rect 1914 10784 1919 10840
rect 0 10782 1919 10784
rect 0 10752 800 10782
rect 1853 10779 1919 10782
rect 24945 10842 25011 10845
rect 25589 10842 25655 10845
rect 30189 10842 30255 10845
rect 32029 10842 32095 10845
rect 35249 10842 35315 10845
rect 24945 10840 30255 10842
rect 24945 10784 24950 10840
rect 25006 10784 25594 10840
rect 25650 10784 30194 10840
rect 30250 10784 30255 10840
rect 24945 10782 30255 10784
rect 24945 10779 25011 10782
rect 25589 10779 25655 10782
rect 30189 10779 30255 10782
rect 31572 10840 35315 10842
rect 31572 10784 32034 10840
rect 32090 10784 35254 10840
rect 35310 10784 35315 10840
rect 31572 10782 35315 10784
rect 19609 10706 19675 10709
rect 28993 10706 29059 10709
rect 19609 10704 29059 10706
rect 19609 10648 19614 10704
rect 19670 10648 28998 10704
rect 29054 10648 29059 10704
rect 19609 10646 29059 10648
rect 19609 10643 19675 10646
rect 28993 10643 29059 10646
rect 29177 10706 29243 10709
rect 31572 10706 31632 10782
rect 32029 10779 32095 10782
rect 35249 10779 35315 10782
rect 29177 10704 31632 10706
rect 29177 10648 29182 10704
rect 29238 10648 31632 10704
rect 29177 10646 31632 10648
rect 31753 10706 31819 10709
rect 32121 10706 32187 10709
rect 31753 10704 32187 10706
rect 31753 10648 31758 10704
rect 31814 10648 32126 10704
rect 32182 10648 32187 10704
rect 31753 10646 32187 10648
rect 29177 10643 29243 10646
rect 31753 10643 31819 10646
rect 32121 10643 32187 10646
rect 33409 10706 33475 10709
rect 36077 10706 36143 10709
rect 33409 10704 36143 10706
rect 33409 10648 33414 10704
rect 33470 10648 36082 10704
rect 36138 10648 36143 10704
rect 33409 10646 36143 10648
rect 33409 10643 33475 10646
rect 36077 10643 36143 10646
rect 9489 10570 9555 10573
rect 36537 10570 36603 10573
rect 9489 10568 36603 10570
rect 9489 10512 9494 10568
rect 9550 10512 36542 10568
rect 36598 10512 36603 10568
rect 9489 10510 36603 10512
rect 9489 10507 9555 10510
rect 36537 10507 36603 10510
rect 17769 10434 17835 10437
rect 23105 10434 23171 10437
rect 26049 10436 26115 10437
rect 25998 10434 26004 10436
rect 17769 10432 23171 10434
rect 17769 10376 17774 10432
rect 17830 10376 23110 10432
rect 23166 10376 23171 10432
rect 17769 10374 23171 10376
rect 25958 10374 26004 10434
rect 26068 10432 26115 10436
rect 26110 10376 26115 10432
rect 17769 10371 17835 10374
rect 23105 10371 23171 10374
rect 25998 10372 26004 10374
rect 26068 10372 26115 10376
rect 26049 10371 26115 10372
rect 27245 10434 27311 10437
rect 31569 10434 31635 10437
rect 34421 10434 34487 10437
rect 27245 10432 34487 10434
rect 27245 10376 27250 10432
rect 27306 10376 31574 10432
rect 31630 10376 34426 10432
rect 34482 10376 34487 10432
rect 27245 10374 34487 10376
rect 27245 10371 27311 10374
rect 31569 10371 31635 10374
rect 34421 10371 34487 10374
rect 58157 10434 58223 10437
rect 59200 10434 60000 10464
rect 58157 10432 60000 10434
rect 58157 10376 58162 10432
rect 58218 10376 60000 10432
rect 58157 10374 60000 10376
rect 58157 10371 58223 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 59200 10344 60000 10374
rect 34930 10303 35246 10304
rect 6821 10298 6887 10301
rect 17677 10298 17743 10301
rect 6821 10296 17743 10298
rect 6821 10240 6826 10296
rect 6882 10240 17682 10296
rect 17738 10240 17743 10296
rect 6821 10238 17743 10240
rect 6821 10235 6887 10238
rect 17677 10235 17743 10238
rect 19793 10298 19859 10301
rect 28901 10298 28967 10301
rect 19793 10296 28967 10298
rect 19793 10240 19798 10296
rect 19854 10240 28906 10296
rect 28962 10240 28967 10296
rect 19793 10238 28967 10240
rect 19793 10235 19859 10238
rect 28901 10235 28967 10238
rect 38745 10298 38811 10301
rect 44541 10298 44607 10301
rect 38745 10296 44607 10298
rect 38745 10240 38750 10296
rect 38806 10240 44546 10296
rect 44602 10240 44607 10296
rect 38745 10238 44607 10240
rect 38745 10235 38811 10238
rect 44541 10235 44607 10238
rect 0 10162 800 10192
rect 1761 10162 1827 10165
rect 0 10160 1827 10162
rect 0 10104 1766 10160
rect 1822 10104 1827 10160
rect 0 10102 1827 10104
rect 0 10072 800 10102
rect 1761 10099 1827 10102
rect 21909 10162 21975 10165
rect 22093 10162 22159 10165
rect 21909 10160 22159 10162
rect 21909 10104 21914 10160
rect 21970 10104 22098 10160
rect 22154 10104 22159 10160
rect 21909 10102 22159 10104
rect 21909 10099 21975 10102
rect 22093 10099 22159 10102
rect 23013 10162 23079 10165
rect 27889 10162 27955 10165
rect 23013 10160 27955 10162
rect 23013 10104 23018 10160
rect 23074 10104 27894 10160
rect 27950 10104 27955 10160
rect 23013 10102 27955 10104
rect 23013 10099 23079 10102
rect 27889 10099 27955 10102
rect 29453 10162 29519 10165
rect 35525 10162 35591 10165
rect 29453 10160 35591 10162
rect 29453 10104 29458 10160
rect 29514 10104 35530 10160
rect 35586 10104 35591 10160
rect 29453 10102 35591 10104
rect 29453 10099 29519 10102
rect 35525 10099 35591 10102
rect 38653 10162 38719 10165
rect 42885 10162 42951 10165
rect 38653 10160 42951 10162
rect 38653 10104 38658 10160
rect 38714 10104 42890 10160
rect 42946 10104 42951 10160
rect 38653 10102 42951 10104
rect 38653 10099 38719 10102
rect 42885 10099 42951 10102
rect 1577 10026 1643 10029
rect 27613 10026 27679 10029
rect 1577 10024 27679 10026
rect 1577 9968 1582 10024
rect 1638 9968 27618 10024
rect 27674 9968 27679 10024
rect 1577 9966 27679 9968
rect 1577 9963 1643 9966
rect 27613 9963 27679 9966
rect 28717 10026 28783 10029
rect 32213 10026 32279 10029
rect 28717 10024 32279 10026
rect 28717 9968 28722 10024
rect 28778 9968 32218 10024
rect 32274 9968 32279 10024
rect 28717 9966 32279 9968
rect 28717 9963 28783 9966
rect 32213 9963 32279 9966
rect 36169 10026 36235 10029
rect 38837 10026 38903 10029
rect 36169 10024 38903 10026
rect 36169 9968 36174 10024
rect 36230 9968 38842 10024
rect 38898 9968 38903 10024
rect 36169 9966 38903 9968
rect 36169 9963 36235 9966
rect 38837 9963 38903 9966
rect 23381 9890 23447 9893
rect 25773 9890 25839 9893
rect 23381 9888 25839 9890
rect 23381 9832 23386 9888
rect 23442 9832 25778 9888
rect 25834 9832 25839 9888
rect 23381 9830 25839 9832
rect 23381 9827 23447 9830
rect 25773 9827 25839 9830
rect 28533 9890 28599 9893
rect 38653 9890 38719 9893
rect 28533 9888 38719 9890
rect 28533 9832 28538 9888
rect 28594 9832 38658 9888
rect 38714 9832 38719 9888
rect 28533 9830 38719 9832
rect 28533 9827 28599 9830
rect 38653 9827 38719 9830
rect 57053 9890 57119 9893
rect 59200 9890 60000 9920
rect 57053 9888 60000 9890
rect 57053 9832 57058 9888
rect 57114 9832 60000 9888
rect 57053 9830 60000 9832
rect 57053 9827 57119 9830
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 59200 9800 60000 9830
rect 50290 9759 50606 9760
rect 23381 9754 23447 9757
rect 25589 9754 25655 9757
rect 23381 9752 25655 9754
rect 23381 9696 23386 9752
rect 23442 9696 25594 9752
rect 25650 9696 25655 9752
rect 23381 9694 25655 9696
rect 23381 9691 23447 9694
rect 25589 9691 25655 9694
rect 29545 9754 29611 9757
rect 30005 9754 30071 9757
rect 29545 9752 30071 9754
rect 29545 9696 29550 9752
rect 29606 9696 30010 9752
rect 30066 9696 30071 9752
rect 29545 9694 30071 9696
rect 29545 9691 29611 9694
rect 30005 9691 30071 9694
rect 38745 9754 38811 9757
rect 39113 9754 39179 9757
rect 38745 9752 39179 9754
rect 38745 9696 38750 9752
rect 38806 9696 39118 9752
rect 39174 9696 39179 9752
rect 38745 9694 39179 9696
rect 38745 9691 38811 9694
rect 39113 9691 39179 9694
rect 15929 9618 15995 9621
rect 26417 9618 26483 9621
rect 15929 9616 26483 9618
rect 15929 9560 15934 9616
rect 15990 9560 26422 9616
rect 26478 9560 26483 9616
rect 15929 9558 26483 9560
rect 15929 9555 15995 9558
rect 26417 9555 26483 9558
rect 26601 9618 26667 9621
rect 27797 9618 27863 9621
rect 26601 9616 27863 9618
rect 26601 9560 26606 9616
rect 26662 9560 27802 9616
rect 27858 9560 27863 9616
rect 26601 9558 27863 9560
rect 26601 9555 26667 9558
rect 27797 9555 27863 9558
rect 28441 9618 28507 9621
rect 28809 9620 28875 9621
rect 28574 9618 28580 9620
rect 28441 9616 28580 9618
rect 28441 9560 28446 9616
rect 28502 9560 28580 9616
rect 28441 9558 28580 9560
rect 28441 9555 28507 9558
rect 28574 9556 28580 9558
rect 28644 9556 28650 9620
rect 28758 9618 28764 9620
rect 28718 9558 28764 9618
rect 28828 9616 28875 9620
rect 28870 9560 28875 9616
rect 28758 9556 28764 9558
rect 28828 9556 28875 9560
rect 28809 9555 28875 9556
rect 29729 9618 29795 9621
rect 29862 9618 29868 9620
rect 29729 9616 29868 9618
rect 29729 9560 29734 9616
rect 29790 9560 29868 9616
rect 29729 9558 29868 9560
rect 29729 9555 29795 9558
rect 29862 9556 29868 9558
rect 29932 9556 29938 9620
rect 30189 9618 30255 9621
rect 30649 9618 30715 9621
rect 33409 9618 33475 9621
rect 30189 9616 33475 9618
rect 30189 9560 30194 9616
rect 30250 9560 30654 9616
rect 30710 9560 33414 9616
rect 33470 9560 33475 9616
rect 30189 9558 33475 9560
rect 30189 9555 30255 9558
rect 30649 9555 30715 9558
rect 33409 9555 33475 9558
rect 38745 9618 38811 9621
rect 38745 9616 38946 9618
rect 38745 9560 38750 9616
rect 38806 9560 38946 9616
rect 38745 9558 38946 9560
rect 38745 9555 38811 9558
rect 0 9482 800 9512
rect 1761 9482 1827 9485
rect 0 9480 1827 9482
rect 0 9424 1766 9480
rect 1822 9424 1827 9480
rect 0 9422 1827 9424
rect 0 9392 800 9422
rect 1761 9419 1827 9422
rect 15285 9482 15351 9485
rect 15837 9482 15903 9485
rect 28942 9482 28948 9484
rect 15285 9480 28948 9482
rect 15285 9424 15290 9480
rect 15346 9424 15842 9480
rect 15898 9424 28948 9480
rect 15285 9422 28948 9424
rect 15285 9419 15351 9422
rect 15837 9419 15903 9422
rect 28942 9420 28948 9422
rect 29012 9420 29018 9484
rect 29545 9482 29611 9485
rect 29678 9482 29684 9484
rect 29545 9480 29684 9482
rect 29545 9424 29550 9480
rect 29606 9424 29684 9480
rect 29545 9422 29684 9424
rect 29545 9419 29611 9422
rect 29678 9420 29684 9422
rect 29748 9420 29754 9484
rect 38886 9482 38946 9558
rect 46933 9482 46999 9485
rect 38886 9480 46999 9482
rect 38886 9424 46938 9480
rect 46994 9424 46999 9480
rect 38886 9422 46999 9424
rect 46933 9419 46999 9422
rect 19241 9348 19307 9349
rect 19190 9346 19196 9348
rect 19114 9286 19196 9346
rect 19260 9346 19307 9348
rect 23381 9346 23447 9349
rect 19260 9344 23447 9346
rect 19302 9288 23386 9344
rect 23442 9288 23447 9344
rect 19190 9284 19196 9286
rect 19260 9286 23447 9288
rect 19260 9284 19307 9286
rect 19241 9283 19307 9284
rect 23381 9283 23447 9286
rect 23565 9346 23631 9349
rect 23841 9346 23907 9349
rect 23565 9344 23907 9346
rect 23565 9288 23570 9344
rect 23626 9288 23846 9344
rect 23902 9288 23907 9344
rect 23565 9286 23907 9288
rect 23565 9283 23631 9286
rect 23841 9283 23907 9286
rect 24301 9346 24367 9349
rect 25497 9346 25563 9349
rect 24301 9344 25563 9346
rect 24301 9288 24306 9344
rect 24362 9288 25502 9344
rect 25558 9288 25563 9344
rect 24301 9286 25563 9288
rect 24301 9283 24367 9286
rect 25497 9283 25563 9286
rect 27153 9346 27219 9349
rect 27286 9346 27292 9348
rect 27153 9344 27292 9346
rect 27153 9288 27158 9344
rect 27214 9288 27292 9344
rect 27153 9286 27292 9288
rect 27153 9283 27219 9286
rect 27286 9284 27292 9286
rect 27356 9284 27362 9348
rect 27521 9346 27587 9349
rect 35525 9346 35591 9349
rect 41873 9346 41939 9349
rect 27521 9344 27630 9346
rect 27521 9288 27526 9344
rect 27582 9288 27630 9344
rect 27521 9283 27630 9288
rect 35525 9344 41939 9346
rect 35525 9288 35530 9344
rect 35586 9288 41878 9344
rect 41934 9288 41939 9344
rect 35525 9286 41939 9288
rect 35525 9283 35591 9286
rect 41873 9283 41939 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 19190 9148 19196 9212
rect 19260 9210 19266 9212
rect 24393 9210 24459 9213
rect 25313 9212 25379 9213
rect 19260 9208 24459 9210
rect 19260 9152 24398 9208
rect 24454 9152 24459 9208
rect 19260 9150 24459 9152
rect 19260 9148 19266 9150
rect 24393 9147 24459 9150
rect 25262 9148 25268 9212
rect 25332 9210 25379 9212
rect 25332 9208 25424 9210
rect 25374 9152 25424 9208
rect 25332 9150 25424 9152
rect 25332 9148 25379 9150
rect 25313 9147 25379 9148
rect 19006 9012 19012 9076
rect 19076 9074 19082 9076
rect 19149 9074 19215 9077
rect 19076 9072 19215 9074
rect 19076 9016 19154 9072
rect 19210 9016 19215 9072
rect 19076 9014 19215 9016
rect 19076 9012 19082 9014
rect 19149 9011 19215 9014
rect 19374 9012 19380 9076
rect 19444 9074 19450 9076
rect 24669 9074 24735 9077
rect 19444 9072 24735 9074
rect 19444 9016 24674 9072
rect 24730 9016 24735 9072
rect 19444 9014 24735 9016
rect 27570 9074 27630 9283
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 59200 9256 60000 9376
rect 34930 9215 35246 9216
rect 31845 9210 31911 9213
rect 33225 9210 33291 9213
rect 31845 9208 33291 9210
rect 31845 9152 31850 9208
rect 31906 9152 33230 9208
rect 33286 9152 33291 9208
rect 31845 9150 33291 9152
rect 31845 9147 31911 9150
rect 33225 9147 33291 9150
rect 38377 9210 38443 9213
rect 46013 9210 46079 9213
rect 38377 9208 46079 9210
rect 38377 9152 38382 9208
rect 38438 9152 46018 9208
rect 46074 9152 46079 9208
rect 38377 9150 46079 9152
rect 38377 9147 38443 9150
rect 46013 9147 46079 9150
rect 32305 9074 32371 9077
rect 27570 9072 32371 9074
rect 27570 9016 32310 9072
rect 32366 9016 32371 9072
rect 27570 9014 32371 9016
rect 19444 9012 19450 9014
rect 24669 9011 24735 9014
rect 32305 9011 32371 9014
rect 36445 9074 36511 9077
rect 38561 9074 38627 9077
rect 36445 9072 38627 9074
rect 36445 9016 36450 9072
rect 36506 9016 38566 9072
rect 38622 9016 38627 9072
rect 36445 9014 38627 9016
rect 36445 9011 36511 9014
rect 38561 9011 38627 9014
rect 8293 8938 8359 8941
rect 22461 8938 22527 8941
rect 8293 8936 22527 8938
rect 8293 8880 8298 8936
rect 8354 8880 22466 8936
rect 22522 8880 22527 8936
rect 8293 8878 22527 8880
rect 8293 8875 8359 8878
rect 22461 8875 22527 8878
rect 22645 8938 22711 8941
rect 27981 8938 28047 8941
rect 34329 8938 34395 8941
rect 22645 8936 28047 8938
rect 22645 8880 22650 8936
rect 22706 8880 27986 8936
rect 28042 8880 28047 8936
rect 22645 8878 28047 8880
rect 22645 8875 22711 8878
rect 27981 8875 28047 8878
rect 30238 8936 34395 8938
rect 30238 8880 34334 8936
rect 34390 8880 34395 8936
rect 30238 8878 34395 8880
rect 0 8802 800 8832
rect 1853 8802 1919 8805
rect 0 8800 1919 8802
rect 0 8744 1858 8800
rect 1914 8744 1919 8800
rect 0 8742 1919 8744
rect 0 8712 800 8742
rect 1853 8739 1919 8742
rect 12893 8802 12959 8805
rect 19149 8802 19215 8805
rect 12893 8800 19215 8802
rect 12893 8744 12898 8800
rect 12954 8744 19154 8800
rect 19210 8744 19215 8800
rect 12893 8742 19215 8744
rect 12893 8739 12959 8742
rect 19149 8739 19215 8742
rect 22737 8802 22803 8805
rect 24117 8802 24183 8805
rect 22737 8800 24183 8802
rect 22737 8744 22742 8800
rect 22798 8744 24122 8800
rect 24178 8744 24183 8800
rect 22737 8742 24183 8744
rect 22737 8739 22803 8742
rect 24117 8739 24183 8742
rect 28942 8740 28948 8804
rect 29012 8802 29018 8804
rect 30238 8802 30298 8878
rect 34329 8875 34395 8878
rect 37089 8938 37155 8941
rect 39389 8938 39455 8941
rect 40217 8938 40283 8941
rect 37089 8936 40283 8938
rect 37089 8880 37094 8936
rect 37150 8880 39394 8936
rect 39450 8880 40222 8936
rect 40278 8880 40283 8936
rect 37089 8878 40283 8880
rect 37089 8875 37155 8878
rect 39389 8875 39455 8878
rect 40217 8875 40283 8878
rect 29012 8742 30298 8802
rect 31569 8802 31635 8805
rect 32949 8802 33015 8805
rect 36629 8802 36695 8805
rect 31569 8800 36695 8802
rect 31569 8744 31574 8800
rect 31630 8744 32954 8800
rect 33010 8744 36634 8800
rect 36690 8744 36695 8800
rect 31569 8742 36695 8744
rect 29012 8740 29018 8742
rect 31569 8739 31635 8742
rect 32949 8739 33015 8742
rect 36629 8739 36695 8742
rect 57329 8802 57395 8805
rect 59200 8802 60000 8832
rect 57329 8800 60000 8802
rect 57329 8744 57334 8800
rect 57390 8744 60000 8800
rect 57329 8742 60000 8744
rect 57329 8739 57395 8742
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 59200 8712 60000 8742
rect 50290 8671 50606 8672
rect 17033 8666 17099 8669
rect 19374 8666 19380 8668
rect 17033 8664 19380 8666
rect 17033 8608 17038 8664
rect 17094 8608 19380 8664
rect 17033 8606 19380 8608
rect 17033 8603 17099 8606
rect 19374 8604 19380 8606
rect 19444 8604 19450 8668
rect 20345 8666 20411 8669
rect 24301 8666 24367 8669
rect 20345 8664 24367 8666
rect 20345 8608 20350 8664
rect 20406 8608 24306 8664
rect 24362 8608 24367 8664
rect 20345 8606 24367 8608
rect 20345 8603 20411 8606
rect 24301 8603 24367 8606
rect 28758 8604 28764 8668
rect 28828 8666 28834 8668
rect 31661 8666 31727 8669
rect 37457 8666 37523 8669
rect 38285 8666 38351 8669
rect 28828 8664 31727 8666
rect 28828 8608 31666 8664
rect 31722 8608 31727 8664
rect 28828 8606 31727 8608
rect 28828 8604 28834 8606
rect 31661 8603 31727 8606
rect 31848 8664 38351 8666
rect 31848 8608 37462 8664
rect 37518 8608 38290 8664
rect 38346 8608 38351 8664
rect 31848 8606 38351 8608
rect 17493 8530 17559 8533
rect 26141 8530 26207 8533
rect 28165 8530 28231 8533
rect 17493 8528 28231 8530
rect 17493 8472 17498 8528
rect 17554 8472 26146 8528
rect 26202 8472 28170 8528
rect 28226 8472 28231 8528
rect 17493 8470 28231 8472
rect 17493 8467 17559 8470
rect 26141 8467 26207 8470
rect 28165 8467 28231 8470
rect 29545 8530 29611 8533
rect 31848 8530 31908 8606
rect 37457 8603 37523 8606
rect 38285 8603 38351 8606
rect 29545 8528 31908 8530
rect 29545 8472 29550 8528
rect 29606 8472 31908 8528
rect 29545 8470 31908 8472
rect 32765 8530 32831 8533
rect 33869 8530 33935 8533
rect 38469 8530 38535 8533
rect 32765 8528 38535 8530
rect 32765 8472 32770 8528
rect 32826 8472 33874 8528
rect 33930 8472 38474 8528
rect 38530 8472 38535 8528
rect 32765 8470 38535 8472
rect 29545 8467 29611 8470
rect 32765 8467 32831 8470
rect 33869 8467 33935 8470
rect 38469 8467 38535 8470
rect 18505 8394 18571 8397
rect 21081 8394 21147 8397
rect 18505 8392 21147 8394
rect 18505 8336 18510 8392
rect 18566 8336 21086 8392
rect 21142 8336 21147 8392
rect 18505 8334 21147 8336
rect 18505 8331 18571 8334
rect 21081 8331 21147 8334
rect 24669 8394 24735 8397
rect 26693 8394 26759 8397
rect 31293 8394 31359 8397
rect 24669 8392 31359 8394
rect 24669 8336 24674 8392
rect 24730 8336 26698 8392
rect 26754 8336 31298 8392
rect 31354 8336 31359 8392
rect 24669 8334 31359 8336
rect 24669 8331 24735 8334
rect 26693 8331 26759 8334
rect 31293 8331 31359 8334
rect 31661 8394 31727 8397
rect 37457 8394 37523 8397
rect 31661 8392 37523 8394
rect 31661 8336 31666 8392
rect 31722 8336 37462 8392
rect 37518 8336 37523 8392
rect 31661 8334 37523 8336
rect 31661 8331 31727 8334
rect 37457 8331 37523 8334
rect 15101 8258 15167 8261
rect 15745 8258 15811 8261
rect 24945 8258 25011 8261
rect 15101 8256 25011 8258
rect 15101 8200 15106 8256
rect 15162 8200 15750 8256
rect 15806 8200 24950 8256
rect 25006 8200 25011 8256
rect 15101 8198 25011 8200
rect 15101 8195 15167 8198
rect 15745 8195 15811 8198
rect 24945 8195 25011 8198
rect 30925 8260 30991 8261
rect 30925 8256 30972 8260
rect 31036 8258 31042 8260
rect 30925 8200 30930 8256
rect 30925 8196 30972 8200
rect 31036 8198 31082 8258
rect 31036 8196 31042 8198
rect 31886 8196 31892 8260
rect 31956 8258 31962 8260
rect 32489 8258 32555 8261
rect 31956 8256 32555 8258
rect 31956 8200 32494 8256
rect 32550 8200 32555 8256
rect 31956 8198 32555 8200
rect 31956 8196 31962 8198
rect 30925 8195 30991 8196
rect 32489 8195 32555 8198
rect 56225 8258 56291 8261
rect 59200 8258 60000 8288
rect 56225 8256 60000 8258
rect 56225 8200 56230 8256
rect 56286 8200 60000 8256
rect 56225 8198 60000 8200
rect 56225 8195 56291 8198
rect 4210 8192 4526 8193
rect 0 8122 800 8152
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 59200 8168 60000 8198
rect 34930 8127 35246 8128
rect 1761 8122 1827 8125
rect 0 8120 1827 8122
rect 0 8064 1766 8120
rect 1822 8064 1827 8120
rect 0 8062 1827 8064
rect 0 8032 800 8062
rect 1761 8059 1827 8062
rect 15285 8122 15351 8125
rect 19977 8122 20043 8125
rect 15285 8120 20043 8122
rect 15285 8064 15290 8120
rect 15346 8064 19982 8120
rect 20038 8064 20043 8120
rect 15285 8062 20043 8064
rect 15285 8059 15351 8062
rect 19977 8059 20043 8062
rect 38653 8122 38719 8125
rect 47853 8122 47919 8125
rect 38653 8120 47919 8122
rect 38653 8064 38658 8120
rect 38714 8064 47858 8120
rect 47914 8064 47919 8120
rect 38653 8062 47919 8064
rect 38653 8059 38719 8062
rect 47853 8059 47919 8062
rect 7925 7986 7991 7989
rect 36537 7986 36603 7989
rect 7925 7984 36603 7986
rect 7925 7928 7930 7984
rect 7986 7928 36542 7984
rect 36598 7928 36603 7984
rect 7925 7926 36603 7928
rect 7925 7923 7991 7926
rect 36537 7923 36603 7926
rect 38653 7986 38719 7989
rect 39205 7986 39271 7989
rect 38653 7984 39271 7986
rect 38653 7928 38658 7984
rect 38714 7928 39210 7984
rect 39266 7928 39271 7984
rect 38653 7926 39271 7928
rect 38653 7923 38719 7926
rect 39205 7923 39271 7926
rect 16297 7850 16363 7853
rect 25681 7850 25747 7853
rect 16297 7848 25747 7850
rect 16297 7792 16302 7848
rect 16358 7792 25686 7848
rect 25742 7792 25747 7848
rect 16297 7790 25747 7792
rect 16297 7787 16363 7790
rect 25681 7787 25747 7790
rect 19006 7652 19012 7716
rect 19076 7714 19082 7716
rect 19149 7714 19215 7717
rect 19076 7712 19215 7714
rect 19076 7656 19154 7712
rect 19210 7656 19215 7712
rect 19076 7654 19215 7656
rect 19076 7652 19082 7654
rect 19149 7651 19215 7654
rect 30557 7714 30623 7717
rect 31201 7714 31267 7717
rect 30557 7712 31267 7714
rect 30557 7656 30562 7712
rect 30618 7656 31206 7712
rect 31262 7656 31267 7712
rect 30557 7654 31267 7656
rect 30557 7651 30623 7654
rect 31201 7651 31267 7654
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 59200 7624 60000 7744
rect 50290 7583 50606 7584
rect 12525 7578 12591 7581
rect 18965 7578 19031 7581
rect 12525 7576 19031 7578
rect 12525 7520 12530 7576
rect 12586 7520 18970 7576
rect 19026 7520 19031 7576
rect 12525 7518 19031 7520
rect 12525 7515 12591 7518
rect 18965 7515 19031 7518
rect 31477 7578 31543 7581
rect 35433 7578 35499 7581
rect 31477 7576 35499 7578
rect 31477 7520 31482 7576
rect 31538 7520 35438 7576
rect 35494 7520 35499 7576
rect 31477 7518 35499 7520
rect 31477 7515 31543 7518
rect 35433 7515 35499 7518
rect 0 7442 800 7472
rect 1853 7442 1919 7445
rect 0 7440 1919 7442
rect 0 7384 1858 7440
rect 1914 7384 1919 7440
rect 0 7382 1919 7384
rect 0 7352 800 7382
rect 1853 7379 1919 7382
rect 18597 7442 18663 7445
rect 19517 7442 19583 7445
rect 18597 7440 19583 7442
rect 18597 7384 18602 7440
rect 18658 7384 19522 7440
rect 19578 7384 19583 7440
rect 18597 7382 19583 7384
rect 18597 7379 18663 7382
rect 19517 7379 19583 7382
rect 15193 7306 15259 7309
rect 19149 7306 19215 7309
rect 15193 7304 19215 7306
rect 15193 7248 15198 7304
rect 15254 7248 19154 7304
rect 19210 7248 19215 7304
rect 15193 7246 19215 7248
rect 15193 7243 15259 7246
rect 19149 7243 19215 7246
rect 19885 7306 19951 7309
rect 21541 7306 21607 7309
rect 19885 7304 21607 7306
rect 19885 7248 19890 7304
rect 19946 7248 21546 7304
rect 21602 7248 21607 7304
rect 19885 7246 21607 7248
rect 19885 7243 19951 7246
rect 21541 7243 21607 7246
rect 9765 7170 9831 7173
rect 19057 7170 19123 7173
rect 9765 7168 19123 7170
rect 9765 7112 9770 7168
rect 9826 7112 19062 7168
rect 19118 7112 19123 7168
rect 9765 7110 19123 7112
rect 9765 7107 9831 7110
rect 19057 7107 19123 7110
rect 22369 7170 22435 7173
rect 23841 7170 23907 7173
rect 22369 7168 23907 7170
rect 22369 7112 22374 7168
rect 22430 7112 23846 7168
rect 23902 7112 23907 7168
rect 22369 7110 23907 7112
rect 22369 7107 22435 7110
rect 23841 7107 23907 7110
rect 27521 7170 27587 7173
rect 29913 7170 29979 7173
rect 33685 7170 33751 7173
rect 27521 7168 33751 7170
rect 27521 7112 27526 7168
rect 27582 7112 29918 7168
rect 29974 7112 33690 7168
rect 33746 7112 33751 7168
rect 27521 7110 33751 7112
rect 27521 7107 27587 7110
rect 29913 7107 29979 7110
rect 33685 7107 33751 7110
rect 58157 7170 58223 7173
rect 59200 7170 60000 7200
rect 58157 7168 60000 7170
rect 58157 7112 58162 7168
rect 58218 7112 60000 7168
rect 58157 7110 60000 7112
rect 58157 7107 58223 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 59200 7080 60000 7110
rect 34930 7039 35246 7040
rect 17217 7034 17283 7037
rect 30373 7034 30439 7037
rect 30833 7036 30899 7037
rect 17217 7032 30439 7034
rect 17217 6976 17222 7032
rect 17278 6976 30378 7032
rect 30434 6976 30439 7032
rect 17217 6974 30439 6976
rect 17217 6971 17283 6974
rect 30373 6971 30439 6974
rect 30782 6972 30788 7036
rect 30852 7034 30899 7036
rect 30852 7032 30944 7034
rect 30894 6976 30944 7032
rect 30852 6974 30944 6976
rect 30852 6972 30899 6974
rect 30833 6971 30899 6972
rect 39573 6898 39639 6901
rect 39982 6898 39988 6900
rect 39573 6896 39988 6898
rect 39573 6840 39578 6896
rect 39634 6840 39988 6896
rect 39573 6838 39988 6840
rect 39573 6835 39639 6838
rect 39982 6836 39988 6838
rect 40052 6836 40058 6900
rect 0 6762 800 6792
rect 1853 6762 1919 6765
rect 0 6760 1919 6762
rect 0 6704 1858 6760
rect 1914 6704 1919 6760
rect 0 6702 1919 6704
rect 0 6672 800 6702
rect 1853 6699 1919 6702
rect 31477 6762 31543 6765
rect 35801 6762 35867 6765
rect 31477 6760 35867 6762
rect 31477 6704 31482 6760
rect 31538 6704 35806 6760
rect 35862 6704 35867 6760
rect 31477 6702 35867 6704
rect 31477 6699 31543 6702
rect 35801 6699 35867 6702
rect 57145 6626 57211 6629
rect 59200 6626 60000 6656
rect 57145 6624 60000 6626
rect 57145 6568 57150 6624
rect 57206 6568 60000 6624
rect 57145 6566 60000 6568
rect 57145 6563 57211 6566
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 59200 6536 60000 6566
rect 50290 6495 50606 6496
rect 38377 6490 38443 6493
rect 29686 6488 38443 6490
rect 29686 6432 38382 6488
rect 38438 6432 38443 6488
rect 29686 6430 38443 6432
rect 29686 6357 29746 6430
rect 38377 6427 38443 6430
rect 15377 6354 15443 6357
rect 16113 6354 16179 6357
rect 28165 6354 28231 6357
rect 29637 6356 29746 6357
rect 29637 6354 29684 6356
rect 15377 6352 28231 6354
rect 15377 6296 15382 6352
rect 15438 6296 16118 6352
rect 16174 6296 28170 6352
rect 28226 6296 28231 6352
rect 15377 6294 28231 6296
rect 29592 6352 29684 6354
rect 29592 6296 29642 6352
rect 29592 6294 29684 6296
rect 15377 6291 15443 6294
rect 16113 6291 16179 6294
rect 28165 6291 28231 6294
rect 29637 6292 29684 6294
rect 29748 6292 29754 6356
rect 32581 6354 32647 6357
rect 45001 6354 45067 6357
rect 32581 6352 45067 6354
rect 32581 6296 32586 6352
rect 32642 6296 45006 6352
rect 45062 6296 45067 6352
rect 32581 6294 45067 6296
rect 29637 6291 29703 6292
rect 32581 6291 32647 6294
rect 45001 6291 45067 6294
rect 19057 6218 19123 6221
rect 20621 6218 20687 6221
rect 38101 6218 38167 6221
rect 57053 6218 57119 6221
rect 19057 6216 57119 6218
rect 19057 6160 19062 6216
rect 19118 6160 20626 6216
rect 20682 6160 38106 6216
rect 38162 6160 57058 6216
rect 57114 6160 57119 6216
rect 19057 6158 57119 6160
rect 19057 6155 19123 6158
rect 20621 6155 20687 6158
rect 38101 6155 38167 6158
rect 57053 6155 57119 6158
rect 0 6082 800 6112
rect 1761 6082 1827 6085
rect 0 6080 1827 6082
rect 0 6024 1766 6080
rect 1822 6024 1827 6080
rect 0 6022 1827 6024
rect 0 5992 800 6022
rect 1761 6019 1827 6022
rect 14825 6082 14891 6085
rect 29862 6082 29868 6084
rect 14825 6080 29868 6082
rect 14825 6024 14830 6080
rect 14886 6024 29868 6080
rect 14825 6022 29868 6024
rect 14825 6019 14891 6022
rect 29862 6020 29868 6022
rect 29932 6020 29938 6084
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 59200 5992 60000 6112
rect 34930 5951 35246 5952
rect 14457 5946 14523 5949
rect 27153 5946 27219 5949
rect 32857 5946 32923 5949
rect 14457 5944 32923 5946
rect 14457 5888 14462 5944
rect 14518 5888 27158 5944
rect 27214 5888 32862 5944
rect 32918 5888 32923 5944
rect 14457 5886 32923 5888
rect 14457 5883 14523 5886
rect 27153 5883 27219 5886
rect 32857 5883 32923 5886
rect 19517 5810 19583 5813
rect 26233 5810 26299 5813
rect 19517 5808 26299 5810
rect 19517 5752 19522 5808
rect 19578 5752 26238 5808
rect 26294 5752 26299 5808
rect 19517 5750 26299 5752
rect 19517 5747 19583 5750
rect 26233 5747 26299 5750
rect 27797 5810 27863 5813
rect 29729 5810 29795 5813
rect 27797 5808 29795 5810
rect 27797 5752 27802 5808
rect 27858 5752 29734 5808
rect 29790 5752 29795 5808
rect 27797 5750 29795 5752
rect 27797 5747 27863 5750
rect 29729 5747 29795 5750
rect 37406 5748 37412 5812
rect 37476 5810 37482 5812
rect 41965 5810 42031 5813
rect 37476 5808 42031 5810
rect 37476 5752 41970 5808
rect 42026 5752 42031 5808
rect 37476 5750 42031 5752
rect 37476 5748 37482 5750
rect 41965 5747 42031 5750
rect 18873 5674 18939 5677
rect 21817 5674 21883 5677
rect 32213 5674 32279 5677
rect 32581 5674 32647 5677
rect 18873 5672 32647 5674
rect 18873 5616 18878 5672
rect 18934 5616 21822 5672
rect 21878 5616 32218 5672
rect 32274 5616 32586 5672
rect 32642 5616 32647 5672
rect 18873 5614 32647 5616
rect 18873 5611 18939 5614
rect 21817 5611 21883 5614
rect 32213 5611 32279 5614
rect 32581 5611 32647 5614
rect 22369 5538 22435 5541
rect 22870 5538 22876 5540
rect 22369 5536 22876 5538
rect 22369 5480 22374 5536
rect 22430 5480 22876 5536
rect 22369 5478 22876 5480
rect 22369 5475 22435 5478
rect 22870 5476 22876 5478
rect 22940 5476 22946 5540
rect 33501 5538 33567 5541
rect 23062 5536 33567 5538
rect 23062 5480 33506 5536
rect 33562 5480 33567 5536
rect 23062 5478 33567 5480
rect 19570 5472 19886 5473
rect 0 5402 800 5432
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 1853 5402 1919 5405
rect 23062 5402 23122 5478
rect 33501 5475 33567 5478
rect 57237 5538 57303 5541
rect 59200 5538 60000 5568
rect 57237 5536 60000 5538
rect 57237 5480 57242 5536
rect 57298 5480 60000 5536
rect 57237 5478 60000 5480
rect 57237 5475 57303 5478
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 59200 5448 60000 5478
rect 50290 5407 50606 5408
rect 0 5400 1919 5402
rect 0 5344 1858 5400
rect 1914 5344 1919 5400
rect 0 5342 1919 5344
rect 0 5312 800 5342
rect 1853 5339 1919 5342
rect 19980 5342 23122 5402
rect 23381 5402 23447 5405
rect 29494 5402 29500 5404
rect 23381 5400 29500 5402
rect 23381 5344 23386 5400
rect 23442 5344 29500 5400
rect 23381 5342 29500 5344
rect 19425 5266 19491 5269
rect 19980 5266 20040 5342
rect 23381 5339 23447 5342
rect 29494 5340 29500 5342
rect 29564 5340 29570 5404
rect 30598 5340 30604 5404
rect 30668 5402 30674 5404
rect 30833 5402 30899 5405
rect 30668 5400 30899 5402
rect 30668 5344 30838 5400
rect 30894 5344 30899 5400
rect 30668 5342 30899 5344
rect 30668 5340 30674 5342
rect 30833 5339 30899 5342
rect 32581 5402 32647 5405
rect 34145 5402 34211 5405
rect 36353 5402 36419 5405
rect 32581 5400 36419 5402
rect 32581 5344 32586 5400
rect 32642 5344 34150 5400
rect 34206 5344 36358 5400
rect 36414 5344 36419 5400
rect 32581 5342 36419 5344
rect 32581 5339 32647 5342
rect 34145 5339 34211 5342
rect 36353 5339 36419 5342
rect 19425 5264 20040 5266
rect 19425 5208 19430 5264
rect 19486 5208 20040 5264
rect 19425 5206 20040 5208
rect 20897 5266 20963 5269
rect 28809 5266 28875 5269
rect 20897 5264 28875 5266
rect 20897 5208 20902 5264
rect 20958 5208 28814 5264
rect 28870 5208 28875 5264
rect 20897 5206 28875 5208
rect 19425 5203 19491 5206
rect 20897 5203 20963 5206
rect 28809 5203 28875 5206
rect 30189 5266 30255 5269
rect 31293 5266 31359 5269
rect 30189 5264 31359 5266
rect 30189 5208 30194 5264
rect 30250 5208 31298 5264
rect 31354 5208 31359 5264
rect 30189 5206 31359 5208
rect 30189 5203 30255 5206
rect 31293 5203 31359 5206
rect 21449 5130 21515 5133
rect 23565 5130 23631 5133
rect 27613 5130 27679 5133
rect 21449 5128 27679 5130
rect 21449 5072 21454 5128
rect 21510 5072 23570 5128
rect 23626 5072 27618 5128
rect 27674 5072 27679 5128
rect 21449 5070 27679 5072
rect 21449 5067 21515 5070
rect 23565 5067 23631 5070
rect 27613 5067 27679 5070
rect 38142 5068 38148 5132
rect 38212 5130 38218 5132
rect 40677 5130 40743 5133
rect 38212 5128 40743 5130
rect 38212 5072 40682 5128
rect 40738 5072 40743 5128
rect 38212 5070 40743 5072
rect 38212 5068 38218 5070
rect 40677 5067 40743 5070
rect 17769 4994 17835 4997
rect 23657 4994 23723 4997
rect 17769 4992 23723 4994
rect 17769 4936 17774 4992
rect 17830 4936 23662 4992
rect 23718 4936 23723 4992
rect 17769 4934 23723 4936
rect 17769 4931 17835 4934
rect 23657 4931 23723 4934
rect 58065 4994 58131 4997
rect 59200 4994 60000 5024
rect 58065 4992 60000 4994
rect 58065 4936 58070 4992
rect 58126 4936 60000 4992
rect 58065 4934 60000 4936
rect 58065 4931 58131 4934
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 59200 4904 60000 4934
rect 34930 4863 35246 4864
rect 16941 4858 17007 4861
rect 33409 4858 33475 4861
rect 16941 4856 33475 4858
rect 16941 4800 16946 4856
rect 17002 4800 33414 4856
rect 33470 4800 33475 4856
rect 16941 4798 33475 4800
rect 16941 4795 17007 4798
rect 33409 4795 33475 4798
rect 0 4722 800 4752
rect 1761 4722 1827 4725
rect 0 4720 1827 4722
rect 0 4664 1766 4720
rect 1822 4664 1827 4720
rect 0 4662 1827 4664
rect 0 4632 800 4662
rect 1761 4659 1827 4662
rect 9857 4722 9923 4725
rect 18965 4722 19031 4725
rect 9857 4720 19031 4722
rect 9857 4664 9862 4720
rect 9918 4664 18970 4720
rect 19026 4664 19031 4720
rect 9857 4662 19031 4664
rect 9857 4659 9923 4662
rect 18965 4659 19031 4662
rect 27153 4722 27219 4725
rect 28717 4722 28783 4725
rect 27153 4720 28783 4722
rect 27153 4664 27158 4720
rect 27214 4664 28722 4720
rect 28778 4664 28783 4720
rect 27153 4662 28783 4664
rect 27153 4659 27219 4662
rect 28717 4659 28783 4662
rect 31937 4722 32003 4725
rect 34605 4722 34671 4725
rect 31937 4720 34671 4722
rect 31937 4664 31942 4720
rect 31998 4664 34610 4720
rect 34666 4664 34671 4720
rect 31937 4662 34671 4664
rect 31937 4659 32003 4662
rect 34605 4659 34671 4662
rect 19425 4588 19491 4589
rect 19374 4586 19380 4588
rect 19334 4526 19380 4586
rect 19444 4584 19491 4588
rect 19486 4528 19491 4584
rect 19374 4524 19380 4526
rect 19444 4524 19491 4528
rect 19425 4523 19491 4524
rect 19885 4586 19951 4589
rect 20805 4586 20871 4589
rect 19885 4584 20871 4586
rect 19885 4528 19890 4584
rect 19946 4528 20810 4584
rect 20866 4528 20871 4584
rect 19885 4526 20871 4528
rect 19885 4523 19951 4526
rect 20805 4523 20871 4526
rect 24393 4586 24459 4589
rect 31477 4586 31543 4589
rect 24393 4584 31543 4586
rect 24393 4528 24398 4584
rect 24454 4528 31482 4584
rect 31538 4528 31543 4584
rect 24393 4526 31543 4528
rect 24393 4523 24459 4526
rect 31477 4523 31543 4526
rect 43345 4586 43411 4589
rect 43989 4586 44055 4589
rect 43345 4584 44055 4586
rect 43345 4528 43350 4584
rect 43406 4528 43994 4584
rect 44050 4528 44055 4584
rect 43345 4526 44055 4528
rect 43345 4523 43411 4526
rect 43989 4523 44055 4526
rect 19333 4450 19399 4453
rect 19290 4448 19399 4450
rect 19290 4392 19338 4448
rect 19394 4392 19399 4448
rect 19290 4387 19399 4392
rect 32213 4450 32279 4453
rect 33133 4450 33199 4453
rect 32213 4448 33199 4450
rect 32213 4392 32218 4448
rect 32274 4392 33138 4448
rect 33194 4392 33199 4448
rect 32213 4390 33199 4392
rect 32213 4387 32279 4390
rect 33133 4387 33199 4390
rect 19290 4317 19350 4387
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 59200 4360 60000 4480
rect 50290 4319 50606 4320
rect 19290 4312 19399 4317
rect 19290 4256 19338 4312
rect 19394 4256 19399 4312
rect 19290 4254 19399 4256
rect 19333 4251 19399 4254
rect 19517 4178 19583 4181
rect 21081 4178 21147 4181
rect 45001 4178 45067 4181
rect 19517 4176 21147 4178
rect 19517 4120 19522 4176
rect 19578 4120 21086 4176
rect 21142 4120 21147 4176
rect 19517 4118 21147 4120
rect 19517 4115 19583 4118
rect 21081 4115 21147 4118
rect 43348 4176 45067 4178
rect 43348 4120 45006 4176
rect 45062 4120 45067 4176
rect 43348 4118 45067 4120
rect 0 4042 800 4072
rect 43348 4045 43408 4118
rect 45001 4115 45067 4118
rect 1761 4042 1827 4045
rect 0 4040 1827 4042
rect 0 3984 1766 4040
rect 1822 3984 1827 4040
rect 0 3982 1827 3984
rect 0 3952 800 3982
rect 1761 3979 1827 3982
rect 5901 4042 5967 4045
rect 8569 4042 8635 4045
rect 5901 4040 8635 4042
rect 5901 3984 5906 4040
rect 5962 3984 8574 4040
rect 8630 3984 8635 4040
rect 5901 3982 8635 3984
rect 5901 3979 5967 3982
rect 8569 3979 8635 3982
rect 19425 4042 19491 4045
rect 21173 4042 21239 4045
rect 19425 4040 21239 4042
rect 19425 3984 19430 4040
rect 19486 3984 21178 4040
rect 21234 3984 21239 4040
rect 19425 3982 21239 3984
rect 19425 3979 19491 3982
rect 21173 3979 21239 3982
rect 32765 4042 32831 4045
rect 35985 4042 36051 4045
rect 32765 4040 36051 4042
rect 32765 3984 32770 4040
rect 32826 3984 35990 4040
rect 36046 3984 36051 4040
rect 32765 3982 36051 3984
rect 32765 3979 32831 3982
rect 35985 3979 36051 3982
rect 36261 4044 36327 4045
rect 36261 4040 36308 4044
rect 36372 4042 36378 4044
rect 36261 3984 36266 4040
rect 36261 3980 36308 3984
rect 36372 3982 36418 4042
rect 36372 3980 36378 3982
rect 39982 3980 39988 4044
rect 40052 4042 40058 4044
rect 40125 4042 40191 4045
rect 40052 4040 40191 4042
rect 40052 3984 40130 4040
rect 40186 3984 40191 4040
rect 40052 3982 40191 3984
rect 40052 3980 40058 3982
rect 36261 3979 36327 3980
rect 40125 3979 40191 3982
rect 40534 3980 40540 4044
rect 40604 4042 40610 4044
rect 42609 4042 42675 4045
rect 40604 4040 42675 4042
rect 40604 3984 42614 4040
rect 42670 3984 42675 4040
rect 40604 3982 42675 3984
rect 40604 3980 40610 3982
rect 42609 3979 42675 3982
rect 43345 4040 43411 4045
rect 45185 4044 45251 4045
rect 45134 4042 45140 4044
rect 43345 3984 43350 4040
rect 43406 3984 43411 4040
rect 43345 3979 43411 3984
rect 45094 3982 45140 4042
rect 45204 4040 45251 4044
rect 45246 3984 45251 4040
rect 45134 3980 45140 3982
rect 45204 3980 45251 3984
rect 45185 3979 45251 3980
rect 7649 3906 7715 3909
rect 9397 3906 9463 3909
rect 7649 3904 9463 3906
rect 7649 3848 7654 3904
rect 7710 3848 9402 3904
rect 9458 3848 9463 3904
rect 7649 3846 9463 3848
rect 7649 3843 7715 3846
rect 9397 3843 9463 3846
rect 12525 3906 12591 3909
rect 12985 3906 13051 3909
rect 12525 3904 13051 3906
rect 12525 3848 12530 3904
rect 12586 3848 12990 3904
rect 13046 3848 13051 3904
rect 12525 3846 13051 3848
rect 12525 3843 12591 3846
rect 12985 3843 13051 3846
rect 17953 3906 18019 3909
rect 30373 3906 30439 3909
rect 17953 3904 30439 3906
rect 17953 3848 17958 3904
rect 18014 3848 30378 3904
rect 30434 3848 30439 3904
rect 17953 3846 30439 3848
rect 17953 3843 18019 3846
rect 30373 3843 30439 3846
rect 37365 3906 37431 3909
rect 39941 3906 40007 3909
rect 37365 3904 40007 3906
rect 37365 3848 37370 3904
rect 37426 3848 39946 3904
rect 40002 3848 40007 3904
rect 37365 3846 40007 3848
rect 37365 3843 37431 3846
rect 39941 3843 40007 3846
rect 42701 3906 42767 3909
rect 45461 3906 45527 3909
rect 42701 3904 45527 3906
rect 42701 3848 42706 3904
rect 42762 3848 45466 3904
rect 45522 3848 45527 3904
rect 42701 3846 45527 3848
rect 42701 3843 42767 3846
rect 45461 3843 45527 3846
rect 57881 3906 57947 3909
rect 59200 3906 60000 3936
rect 57881 3904 60000 3906
rect 57881 3848 57886 3904
rect 57942 3848 60000 3904
rect 57881 3846 60000 3848
rect 57881 3843 57947 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 59200 3816 60000 3846
rect 34930 3775 35246 3776
rect 7005 3770 7071 3773
rect 20713 3770 20779 3773
rect 7005 3768 20779 3770
rect 7005 3712 7010 3768
rect 7066 3712 20718 3768
rect 20774 3712 20779 3768
rect 7005 3710 20779 3712
rect 7005 3707 7071 3710
rect 20713 3707 20779 3710
rect 27061 3770 27127 3773
rect 27705 3770 27771 3773
rect 27061 3768 27771 3770
rect 27061 3712 27066 3768
rect 27122 3712 27710 3768
rect 27766 3712 27771 3768
rect 27061 3710 27771 3712
rect 27061 3707 27127 3710
rect 27705 3707 27771 3710
rect 43437 3770 43503 3773
rect 46841 3770 46907 3773
rect 43437 3768 46907 3770
rect 43437 3712 43442 3768
rect 43498 3712 46846 3768
rect 46902 3712 46907 3768
rect 43437 3710 46907 3712
rect 43437 3707 43503 3710
rect 46841 3707 46907 3710
rect 18413 3634 18479 3637
rect 19190 3634 19196 3636
rect 18413 3632 19196 3634
rect 18413 3576 18418 3632
rect 18474 3576 19196 3632
rect 18413 3574 19196 3576
rect 18413 3571 18479 3574
rect 19190 3572 19196 3574
rect 19260 3572 19266 3636
rect 19517 3634 19583 3637
rect 20897 3634 20963 3637
rect 19517 3632 20963 3634
rect 19517 3576 19522 3632
rect 19578 3576 20902 3632
rect 20958 3576 20963 3632
rect 19517 3574 20963 3576
rect 19517 3571 19583 3574
rect 20897 3571 20963 3574
rect 24853 3634 24919 3637
rect 28073 3634 28139 3637
rect 24853 3632 28139 3634
rect 24853 3576 24858 3632
rect 24914 3576 28078 3632
rect 28134 3576 28139 3632
rect 24853 3574 28139 3576
rect 24853 3571 24919 3574
rect 28073 3571 28139 3574
rect 43662 3572 43668 3636
rect 43732 3634 43738 3636
rect 43805 3634 43871 3637
rect 43732 3632 43871 3634
rect 43732 3576 43810 3632
rect 43866 3576 43871 3632
rect 43732 3574 43871 3576
rect 43732 3572 43738 3574
rect 43805 3571 43871 3574
rect 44173 3634 44239 3637
rect 47485 3634 47551 3637
rect 44173 3632 47551 3634
rect 44173 3576 44178 3632
rect 44234 3576 47490 3632
rect 47546 3576 47551 3632
rect 44173 3574 47551 3576
rect 44173 3571 44239 3574
rect 47485 3571 47551 3574
rect 12893 3498 12959 3501
rect 27245 3498 27311 3501
rect 12893 3496 27311 3498
rect 12893 3440 12898 3496
rect 12954 3440 27250 3496
rect 27306 3440 27311 3496
rect 12893 3438 27311 3440
rect 12893 3435 12959 3438
rect 27245 3435 27311 3438
rect 0 3362 800 3392
rect 1853 3362 1919 3365
rect 0 3360 1919 3362
rect 0 3304 1858 3360
rect 1914 3304 1919 3360
rect 0 3302 1919 3304
rect 0 3272 800 3302
rect 1853 3299 1919 3302
rect 36353 3362 36419 3365
rect 38561 3362 38627 3365
rect 36353 3360 38627 3362
rect 36353 3304 36358 3360
rect 36414 3304 38566 3360
rect 38622 3304 38627 3360
rect 36353 3302 38627 3304
rect 36353 3299 36419 3302
rect 38561 3299 38627 3302
rect 58157 3362 58223 3365
rect 59200 3362 60000 3392
rect 58157 3360 60000 3362
rect 58157 3304 58162 3360
rect 58218 3304 60000 3360
rect 58157 3302 60000 3304
rect 58157 3299 58223 3302
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 59200 3272 60000 3302
rect 50290 3231 50606 3232
rect 22277 3226 22343 3229
rect 32438 3226 32444 3228
rect 22277 3224 32444 3226
rect 22277 3168 22282 3224
rect 22338 3168 32444 3224
rect 22277 3166 32444 3168
rect 22277 3163 22343 3166
rect 32438 3164 32444 3166
rect 32508 3164 32514 3228
rect 9581 3090 9647 3093
rect 27153 3090 27219 3093
rect 27521 3090 27587 3093
rect 9581 3088 27587 3090
rect 9581 3032 9586 3088
rect 9642 3032 27158 3088
rect 27214 3032 27526 3088
rect 27582 3032 27587 3088
rect 9581 3030 27587 3032
rect 9581 3027 9647 3030
rect 27153 3027 27219 3030
rect 27521 3027 27587 3030
rect 28073 3090 28139 3093
rect 29085 3090 29151 3093
rect 28073 3088 29151 3090
rect 28073 3032 28078 3088
rect 28134 3032 29090 3088
rect 29146 3032 29151 3088
rect 28073 3030 29151 3032
rect 28073 3027 28139 3030
rect 29085 3027 29151 3030
rect 37365 3090 37431 3093
rect 38285 3090 38351 3093
rect 37365 3088 38351 3090
rect 37365 3032 37370 3088
rect 37426 3032 38290 3088
rect 38346 3032 38351 3088
rect 37365 3030 38351 3032
rect 37365 3027 37431 3030
rect 38285 3027 38351 3030
rect 8201 2954 8267 2957
rect 10317 2954 10383 2957
rect 8201 2952 10383 2954
rect 8201 2896 8206 2952
rect 8262 2896 10322 2952
rect 10378 2896 10383 2952
rect 8201 2894 10383 2896
rect 8201 2891 8267 2894
rect 10317 2891 10383 2894
rect 16757 2954 16823 2957
rect 21725 2954 21791 2957
rect 16757 2952 21791 2954
rect 16757 2896 16762 2952
rect 16818 2896 21730 2952
rect 21786 2896 21791 2952
rect 16757 2894 21791 2896
rect 16757 2891 16823 2894
rect 21725 2891 21791 2894
rect 23565 2954 23631 2957
rect 32765 2954 32831 2957
rect 23565 2952 32831 2954
rect 23565 2896 23570 2952
rect 23626 2896 32770 2952
rect 32826 2896 32831 2952
rect 23565 2894 32831 2896
rect 23565 2891 23631 2894
rect 32765 2891 32831 2894
rect 36537 2954 36603 2957
rect 37273 2954 37339 2957
rect 36537 2952 37339 2954
rect 36537 2896 36542 2952
rect 36598 2896 37278 2952
rect 37334 2896 37339 2952
rect 36537 2894 37339 2896
rect 36537 2891 36603 2894
rect 37273 2891 37339 2894
rect 6637 2818 6703 2821
rect 24209 2818 24275 2821
rect 6637 2816 24275 2818
rect 6637 2760 6642 2816
rect 6698 2760 24214 2816
rect 24270 2760 24275 2816
rect 6637 2758 24275 2760
rect 6637 2755 6703 2758
rect 24209 2755 24275 2758
rect 49601 2818 49667 2821
rect 50521 2818 50587 2821
rect 49601 2816 50587 2818
rect 49601 2760 49606 2816
rect 49662 2760 50526 2816
rect 50582 2760 50587 2816
rect 49601 2758 50587 2760
rect 49601 2755 49667 2758
rect 50521 2755 50587 2758
rect 58157 2818 58223 2821
rect 59200 2818 60000 2848
rect 58157 2816 60000 2818
rect 58157 2760 58162 2816
rect 58218 2760 60000 2816
rect 58157 2758 60000 2760
rect 58157 2755 58223 2758
rect 4210 2752 4526 2753
rect 0 2682 800 2712
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 59200 2728 60000 2758
rect 34930 2687 35246 2688
rect 1761 2682 1827 2685
rect 0 2680 1827 2682
rect 0 2624 1766 2680
rect 1822 2624 1827 2680
rect 0 2622 1827 2624
rect 0 2592 800 2622
rect 1761 2619 1827 2622
rect 17493 2684 17559 2685
rect 17493 2680 17540 2684
rect 17604 2682 17610 2684
rect 19885 2682 19951 2685
rect 42609 2684 42675 2685
rect 25446 2682 25452 2684
rect 17493 2624 17498 2680
rect 17493 2620 17540 2624
rect 17604 2622 17650 2682
rect 19885 2680 25452 2682
rect 19885 2624 19890 2680
rect 19946 2624 25452 2680
rect 19885 2622 25452 2624
rect 17604 2620 17610 2622
rect 17493 2619 17559 2620
rect 19885 2619 19951 2622
rect 25446 2620 25452 2622
rect 25516 2620 25522 2684
rect 42558 2682 42564 2684
rect 42518 2622 42564 2682
rect 42628 2680 42675 2684
rect 42670 2624 42675 2680
rect 42558 2620 42564 2622
rect 42628 2620 42675 2624
rect 42609 2619 42675 2620
rect 43345 2682 43411 2685
rect 43621 2682 43687 2685
rect 45369 2684 45435 2685
rect 43345 2680 43687 2682
rect 43345 2624 43350 2680
rect 43406 2624 43626 2680
rect 43682 2624 43687 2680
rect 43345 2622 43687 2624
rect 43345 2619 43411 2622
rect 43621 2619 43687 2622
rect 45318 2620 45324 2684
rect 45388 2682 45435 2684
rect 45388 2680 45480 2682
rect 45430 2624 45480 2680
rect 45388 2622 45480 2624
rect 45388 2620 45435 2622
rect 45369 2619 45435 2620
rect 8937 2546 9003 2549
rect 27889 2546 27955 2549
rect 8937 2544 27955 2546
rect 8937 2488 8942 2544
rect 8998 2488 27894 2544
rect 27950 2488 27955 2544
rect 8937 2486 27955 2488
rect 8937 2483 9003 2486
rect 27889 2483 27955 2486
rect 20989 2410 21055 2413
rect 41086 2410 41092 2412
rect 20989 2408 41092 2410
rect 20989 2352 20994 2408
rect 21050 2352 41092 2408
rect 20989 2350 41092 2352
rect 20989 2347 21055 2350
rect 41086 2348 41092 2350
rect 41156 2348 41162 2412
rect 57329 2274 57395 2277
rect 59200 2274 60000 2304
rect 57329 2272 60000 2274
rect 57329 2216 57334 2272
rect 57390 2216 60000 2272
rect 57329 2214 60000 2216
rect 57329 2211 57395 2214
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 59200 2184 60000 2214
rect 50290 2143 50606 2144
rect 0 2002 800 2032
rect 1853 2002 1919 2005
rect 0 2000 1919 2002
rect 0 1944 1858 2000
rect 1914 1944 1919 2000
rect 0 1942 1919 1944
rect 0 1912 800 1942
rect 1853 1939 1919 1942
rect 19374 1940 19380 2004
rect 19444 2002 19450 2004
rect 19701 2002 19767 2005
rect 19444 2000 19767 2002
rect 19444 1944 19706 2000
rect 19762 1944 19767 2000
rect 19444 1942 19767 1944
rect 19444 1940 19450 1942
rect 19701 1939 19767 1942
rect 57789 1730 57855 1733
rect 59200 1730 60000 1760
rect 57789 1728 60000 1730
rect 57789 1672 57794 1728
rect 57850 1672 60000 1728
rect 57789 1670 60000 1672
rect 57789 1667 57855 1670
rect 59200 1640 60000 1670
rect 55949 1186 56015 1189
rect 59200 1186 60000 1216
rect 55949 1184 60000 1186
rect 55949 1128 55954 1184
rect 56010 1128 60000 1184
rect 55949 1126 60000 1128
rect 55949 1123 56015 1126
rect 59200 1096 60000 1126
<< via3 >>
rect 4216 61500 4280 61504
rect 4216 61444 4220 61500
rect 4220 61444 4276 61500
rect 4276 61444 4280 61500
rect 4216 61440 4280 61444
rect 4296 61500 4360 61504
rect 4296 61444 4300 61500
rect 4300 61444 4356 61500
rect 4356 61444 4360 61500
rect 4296 61440 4360 61444
rect 4376 61500 4440 61504
rect 4376 61444 4380 61500
rect 4380 61444 4436 61500
rect 4436 61444 4440 61500
rect 4376 61440 4440 61444
rect 4456 61500 4520 61504
rect 4456 61444 4460 61500
rect 4460 61444 4516 61500
rect 4516 61444 4520 61500
rect 4456 61440 4520 61444
rect 34936 61500 35000 61504
rect 34936 61444 34940 61500
rect 34940 61444 34996 61500
rect 34996 61444 35000 61500
rect 34936 61440 35000 61444
rect 35016 61500 35080 61504
rect 35016 61444 35020 61500
rect 35020 61444 35076 61500
rect 35076 61444 35080 61500
rect 35016 61440 35080 61444
rect 35096 61500 35160 61504
rect 35096 61444 35100 61500
rect 35100 61444 35156 61500
rect 35156 61444 35160 61500
rect 35096 61440 35160 61444
rect 35176 61500 35240 61504
rect 35176 61444 35180 61500
rect 35180 61444 35236 61500
rect 35236 61444 35240 61500
rect 35176 61440 35240 61444
rect 28580 61100 28644 61164
rect 30052 61100 30116 61164
rect 19576 60956 19640 60960
rect 19576 60900 19580 60956
rect 19580 60900 19636 60956
rect 19636 60900 19640 60956
rect 19576 60896 19640 60900
rect 19656 60956 19720 60960
rect 19656 60900 19660 60956
rect 19660 60900 19716 60956
rect 19716 60900 19720 60956
rect 19656 60896 19720 60900
rect 19736 60956 19800 60960
rect 19736 60900 19740 60956
rect 19740 60900 19796 60956
rect 19796 60900 19800 60956
rect 19736 60896 19800 60900
rect 19816 60956 19880 60960
rect 19816 60900 19820 60956
rect 19820 60900 19876 60956
rect 19876 60900 19880 60956
rect 19816 60896 19880 60900
rect 50296 60956 50360 60960
rect 50296 60900 50300 60956
rect 50300 60900 50356 60956
rect 50356 60900 50360 60956
rect 50296 60896 50360 60900
rect 50376 60956 50440 60960
rect 50376 60900 50380 60956
rect 50380 60900 50436 60956
rect 50436 60900 50440 60956
rect 50376 60896 50440 60900
rect 50456 60956 50520 60960
rect 50456 60900 50460 60956
rect 50460 60900 50516 60956
rect 50516 60900 50520 60956
rect 50456 60896 50520 60900
rect 50536 60956 50600 60960
rect 50536 60900 50540 60956
rect 50540 60900 50596 60956
rect 50596 60900 50600 60956
rect 50536 60896 50600 60900
rect 28764 60692 28828 60756
rect 4216 60412 4280 60416
rect 4216 60356 4220 60412
rect 4220 60356 4276 60412
rect 4276 60356 4280 60412
rect 4216 60352 4280 60356
rect 4296 60412 4360 60416
rect 4296 60356 4300 60412
rect 4300 60356 4356 60412
rect 4356 60356 4360 60412
rect 4296 60352 4360 60356
rect 4376 60412 4440 60416
rect 4376 60356 4380 60412
rect 4380 60356 4436 60412
rect 4436 60356 4440 60412
rect 4376 60352 4440 60356
rect 4456 60412 4520 60416
rect 4456 60356 4460 60412
rect 4460 60356 4516 60412
rect 4516 60356 4520 60412
rect 4456 60352 4520 60356
rect 34936 60412 35000 60416
rect 34936 60356 34940 60412
rect 34940 60356 34996 60412
rect 34996 60356 35000 60412
rect 34936 60352 35000 60356
rect 35016 60412 35080 60416
rect 35016 60356 35020 60412
rect 35020 60356 35076 60412
rect 35076 60356 35080 60412
rect 35016 60352 35080 60356
rect 35096 60412 35160 60416
rect 35096 60356 35100 60412
rect 35100 60356 35156 60412
rect 35156 60356 35160 60412
rect 35096 60352 35160 60356
rect 35176 60412 35240 60416
rect 35176 60356 35180 60412
rect 35180 60356 35236 60412
rect 35236 60356 35240 60412
rect 35176 60352 35240 60356
rect 22508 60344 22572 60348
rect 22508 60288 22558 60344
rect 22558 60288 22572 60344
rect 22508 60284 22572 60288
rect 40540 60012 40604 60076
rect 19576 59868 19640 59872
rect 19576 59812 19580 59868
rect 19580 59812 19636 59868
rect 19636 59812 19640 59868
rect 19576 59808 19640 59812
rect 19656 59868 19720 59872
rect 19656 59812 19660 59868
rect 19660 59812 19716 59868
rect 19716 59812 19720 59868
rect 19656 59808 19720 59812
rect 19736 59868 19800 59872
rect 19736 59812 19740 59868
rect 19740 59812 19796 59868
rect 19796 59812 19800 59868
rect 19736 59808 19800 59812
rect 19816 59868 19880 59872
rect 19816 59812 19820 59868
rect 19820 59812 19876 59868
rect 19876 59812 19880 59868
rect 19816 59808 19880 59812
rect 50296 59868 50360 59872
rect 50296 59812 50300 59868
rect 50300 59812 50356 59868
rect 50356 59812 50360 59868
rect 50296 59808 50360 59812
rect 50376 59868 50440 59872
rect 50376 59812 50380 59868
rect 50380 59812 50436 59868
rect 50436 59812 50440 59868
rect 50376 59808 50440 59812
rect 50456 59868 50520 59872
rect 50456 59812 50460 59868
rect 50460 59812 50516 59868
rect 50516 59812 50520 59868
rect 50456 59808 50520 59812
rect 50536 59868 50600 59872
rect 50536 59812 50540 59868
rect 50540 59812 50596 59868
rect 50596 59812 50600 59868
rect 50536 59808 50600 59812
rect 19196 59332 19260 59396
rect 42564 59332 42628 59396
rect 4216 59324 4280 59328
rect 4216 59268 4220 59324
rect 4220 59268 4276 59324
rect 4276 59268 4280 59324
rect 4216 59264 4280 59268
rect 4296 59324 4360 59328
rect 4296 59268 4300 59324
rect 4300 59268 4356 59324
rect 4356 59268 4360 59324
rect 4296 59264 4360 59268
rect 4376 59324 4440 59328
rect 4376 59268 4380 59324
rect 4380 59268 4436 59324
rect 4436 59268 4440 59324
rect 4376 59264 4440 59268
rect 4456 59324 4520 59328
rect 4456 59268 4460 59324
rect 4460 59268 4516 59324
rect 4516 59268 4520 59324
rect 4456 59264 4520 59268
rect 34936 59324 35000 59328
rect 34936 59268 34940 59324
rect 34940 59268 34996 59324
rect 34996 59268 35000 59324
rect 34936 59264 35000 59268
rect 35016 59324 35080 59328
rect 35016 59268 35020 59324
rect 35020 59268 35076 59324
rect 35076 59268 35080 59324
rect 35016 59264 35080 59268
rect 35096 59324 35160 59328
rect 35096 59268 35100 59324
rect 35100 59268 35156 59324
rect 35156 59268 35160 59324
rect 35096 59264 35160 59268
rect 35176 59324 35240 59328
rect 35176 59268 35180 59324
rect 35180 59268 35236 59324
rect 35236 59268 35240 59324
rect 35176 59264 35240 59268
rect 39252 58924 39316 58988
rect 19576 58780 19640 58784
rect 19576 58724 19580 58780
rect 19580 58724 19636 58780
rect 19636 58724 19640 58780
rect 19576 58720 19640 58724
rect 19656 58780 19720 58784
rect 19656 58724 19660 58780
rect 19660 58724 19716 58780
rect 19716 58724 19720 58780
rect 19656 58720 19720 58724
rect 19736 58780 19800 58784
rect 19736 58724 19740 58780
rect 19740 58724 19796 58780
rect 19796 58724 19800 58780
rect 19736 58720 19800 58724
rect 19816 58780 19880 58784
rect 19816 58724 19820 58780
rect 19820 58724 19876 58780
rect 19876 58724 19880 58780
rect 19816 58720 19880 58724
rect 50296 58780 50360 58784
rect 50296 58724 50300 58780
rect 50300 58724 50356 58780
rect 50356 58724 50360 58780
rect 50296 58720 50360 58724
rect 50376 58780 50440 58784
rect 50376 58724 50380 58780
rect 50380 58724 50436 58780
rect 50436 58724 50440 58780
rect 50376 58720 50440 58724
rect 50456 58780 50520 58784
rect 50456 58724 50460 58780
rect 50460 58724 50516 58780
rect 50516 58724 50520 58780
rect 50456 58720 50520 58724
rect 50536 58780 50600 58784
rect 50536 58724 50540 58780
rect 50540 58724 50596 58780
rect 50596 58724 50600 58780
rect 50536 58720 50600 58724
rect 4216 58236 4280 58240
rect 4216 58180 4220 58236
rect 4220 58180 4276 58236
rect 4276 58180 4280 58236
rect 4216 58176 4280 58180
rect 4296 58236 4360 58240
rect 4296 58180 4300 58236
rect 4300 58180 4356 58236
rect 4356 58180 4360 58236
rect 4296 58176 4360 58180
rect 4376 58236 4440 58240
rect 4376 58180 4380 58236
rect 4380 58180 4436 58236
rect 4436 58180 4440 58236
rect 4376 58176 4440 58180
rect 4456 58236 4520 58240
rect 4456 58180 4460 58236
rect 4460 58180 4516 58236
rect 4516 58180 4520 58236
rect 4456 58176 4520 58180
rect 34936 58236 35000 58240
rect 34936 58180 34940 58236
rect 34940 58180 34996 58236
rect 34996 58180 35000 58236
rect 34936 58176 35000 58180
rect 35016 58236 35080 58240
rect 35016 58180 35020 58236
rect 35020 58180 35076 58236
rect 35076 58180 35080 58236
rect 35016 58176 35080 58180
rect 35096 58236 35160 58240
rect 35096 58180 35100 58236
rect 35100 58180 35156 58236
rect 35156 58180 35160 58236
rect 35096 58176 35160 58180
rect 35176 58236 35240 58240
rect 35176 58180 35180 58236
rect 35180 58180 35236 58236
rect 35236 58180 35240 58236
rect 35176 58176 35240 58180
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 43668 57292 43732 57356
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 22876 53952 22940 53956
rect 22876 53896 22890 53952
rect 22890 53896 22940 53952
rect 22876 53892 22940 53896
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 36308 50220 36372 50284
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 42932 48860 42996 48924
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 38148 45324 38212 45388
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 27292 43148 27356 43212
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 37412 42604 37476 42668
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 39068 42060 39132 42124
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 57284 41576 57348 41580
rect 57284 41520 57334 41576
rect 57334 41520 57348 41576
rect 57284 41516 57348 41520
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 40724 37708 40788 37772
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 25268 34580 25332 34644
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 26004 33356 26068 33420
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 45324 29548 45388 29612
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 32444 27508 32508 27572
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 22508 25528 22572 25532
rect 22508 25472 22558 25528
rect 22558 25472 22572 25528
rect 22508 25468 22572 25472
rect 17540 25196 17604 25260
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 57284 19892 57348 19956
rect 22876 19756 22940 19820
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 30788 18804 30852 18868
rect 30972 18668 31036 18732
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 28028 17988 28092 18052
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 28764 17852 28828 17916
rect 32444 17776 32508 17780
rect 32444 17720 32458 17776
rect 32458 17720 32508 17776
rect 32444 17716 32508 17720
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 38700 17368 38764 17372
rect 38700 17312 38714 17368
rect 38714 17312 38764 17368
rect 38700 17308 38764 17312
rect 25452 17172 25516 17236
rect 28948 16900 29012 16964
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 28028 16492 28092 16556
rect 42932 16552 42996 16556
rect 42932 16496 42946 16552
rect 42946 16496 42996 16552
rect 42932 16492 42996 16496
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 29500 16220 29564 16284
rect 38700 16220 38764 16284
rect 41092 15812 41156 15876
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 30604 14588 30668 14652
rect 31892 14452 31956 14516
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 28948 12956 29012 13020
rect 45140 12956 45204 13020
rect 39068 12548 39132 12612
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 40724 12412 40788 12476
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 39252 11052 39316 11116
rect 30052 10976 30116 10980
rect 30052 10920 30066 10976
rect 30066 10920 30116 10976
rect 30052 10916 30116 10920
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 26004 10432 26068 10436
rect 26004 10376 26054 10432
rect 26054 10376 26068 10432
rect 26004 10372 26068 10376
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 28580 9556 28644 9620
rect 28764 9616 28828 9620
rect 28764 9560 28814 9616
rect 28814 9560 28828 9616
rect 28764 9556 28828 9560
rect 29868 9556 29932 9620
rect 28948 9420 29012 9484
rect 29684 9420 29748 9484
rect 19196 9344 19260 9348
rect 19196 9288 19246 9344
rect 19246 9288 19260 9344
rect 19196 9284 19260 9288
rect 27292 9284 27356 9348
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 19196 9148 19260 9212
rect 25268 9208 25332 9212
rect 25268 9152 25318 9208
rect 25318 9152 25332 9208
rect 25268 9148 25332 9152
rect 19012 9012 19076 9076
rect 19380 9012 19444 9076
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 28948 8740 29012 8804
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 19380 8604 19444 8668
rect 28764 8604 28828 8668
rect 30972 8256 31036 8260
rect 30972 8200 30986 8256
rect 30986 8200 31036 8256
rect 30972 8196 31036 8200
rect 31892 8196 31956 8260
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19012 7652 19076 7716
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 30788 7032 30852 7036
rect 30788 6976 30838 7032
rect 30838 6976 30852 7032
rect 30788 6972 30852 6976
rect 39988 6836 40052 6900
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 29684 6352 29748 6356
rect 29684 6296 29698 6352
rect 29698 6296 29748 6352
rect 29684 6292 29748 6296
rect 29868 6020 29932 6084
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 37412 5748 37476 5812
rect 22876 5476 22940 5540
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 29500 5340 29564 5404
rect 30604 5340 30668 5404
rect 38148 5068 38212 5132
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19380 4584 19444 4588
rect 19380 4528 19430 4584
rect 19430 4528 19444 4584
rect 19380 4524 19444 4528
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 36308 4040 36372 4044
rect 36308 3984 36322 4040
rect 36322 3984 36372 4040
rect 36308 3980 36372 3984
rect 39988 3980 40052 4044
rect 40540 3980 40604 4044
rect 45140 4040 45204 4044
rect 45140 3984 45190 4040
rect 45190 3984 45204 4040
rect 45140 3980 45204 3984
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19196 3572 19260 3636
rect 43668 3572 43732 3636
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 32444 3164 32508 3228
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 17540 2680 17604 2684
rect 17540 2624 17554 2680
rect 17554 2624 17604 2680
rect 17540 2620 17604 2624
rect 25452 2620 25516 2684
rect 42564 2680 42628 2684
rect 42564 2624 42614 2680
rect 42614 2624 42628 2680
rect 42564 2620 42628 2624
rect 45324 2680 45388 2684
rect 45324 2624 45374 2680
rect 45374 2624 45388 2680
rect 45324 2620 45388 2624
rect 41092 2348 41156 2412
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
rect 19380 1940 19444 2004
<< metal4 >>
rect 4208 61504 4528 61520
rect 4208 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4528 61504
rect 4208 60416 4528 61440
rect 4208 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4528 60416
rect 4208 59328 4528 60352
rect 19568 60960 19888 61520
rect 34928 61504 35248 61520
rect 34928 61440 34936 61504
rect 35000 61440 35016 61504
rect 35080 61440 35096 61504
rect 35160 61440 35176 61504
rect 35240 61440 35248 61504
rect 28579 61164 28645 61165
rect 28579 61100 28580 61164
rect 28644 61100 28645 61164
rect 28579 61099 28645 61100
rect 30051 61164 30117 61165
rect 30051 61100 30052 61164
rect 30116 61100 30117 61164
rect 30051 61099 30117 61100
rect 19568 60896 19576 60960
rect 19640 60896 19656 60960
rect 19720 60896 19736 60960
rect 19800 60896 19816 60960
rect 19880 60896 19888 60960
rect 19568 59872 19888 60896
rect 22507 60348 22573 60349
rect 22507 60284 22508 60348
rect 22572 60284 22573 60348
rect 22507 60283 22573 60284
rect 19568 59808 19576 59872
rect 19640 59808 19656 59872
rect 19720 59808 19736 59872
rect 19800 59808 19816 59872
rect 19880 59808 19888 59872
rect 19195 59396 19261 59397
rect 19195 59332 19196 59396
rect 19260 59332 19261 59396
rect 19195 59331 19261 59332
rect 4208 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4528 59328
rect 4208 58240 4528 59264
rect 4208 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4528 58240
rect 4208 57152 4528 58176
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 17539 25260 17605 25261
rect 17539 25196 17540 25260
rect 17604 25196 17605 25260
rect 17539 25195 17605 25196
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 17542 2685 17602 25195
rect 19198 9349 19258 59331
rect 19568 58784 19888 59808
rect 19568 58720 19576 58784
rect 19640 58720 19656 58784
rect 19720 58720 19736 58784
rect 19800 58720 19816 58784
rect 19880 58720 19888 58784
rect 19568 57696 19888 58720
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 22510 25533 22570 60283
rect 22875 53956 22941 53957
rect 22875 53892 22876 53956
rect 22940 53892 22941 53956
rect 22875 53891 22941 53892
rect 22507 25532 22573 25533
rect 22507 25468 22508 25532
rect 22572 25468 22573 25532
rect 22507 25467 22573 25468
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 22878 19821 22938 53891
rect 27291 43212 27357 43213
rect 27291 43148 27292 43212
rect 27356 43148 27357 43212
rect 27291 43147 27357 43148
rect 25267 34644 25333 34645
rect 25267 34580 25268 34644
rect 25332 34580 25333 34644
rect 25267 34579 25333 34580
rect 22875 19820 22941 19821
rect 22875 19756 22876 19820
rect 22940 19756 22941 19820
rect 22875 19755 22941 19756
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19195 9348 19261 9349
rect 19195 9284 19196 9348
rect 19260 9284 19261 9348
rect 19195 9283 19261 9284
rect 19195 9212 19261 9213
rect 19195 9148 19196 9212
rect 19260 9148 19261 9212
rect 19195 9147 19261 9148
rect 19011 9076 19077 9077
rect 19011 9012 19012 9076
rect 19076 9012 19077 9076
rect 19011 9011 19077 9012
rect 19014 7717 19074 9011
rect 19011 7716 19077 7717
rect 19011 7652 19012 7716
rect 19076 7652 19077 7716
rect 19011 7651 19077 7652
rect 19198 3637 19258 9147
rect 19379 9076 19445 9077
rect 19379 9012 19380 9076
rect 19444 9012 19445 9076
rect 19379 9011 19445 9012
rect 19382 8669 19442 9011
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19379 8668 19445 8669
rect 19379 8604 19380 8668
rect 19444 8604 19445 8668
rect 19379 8603 19445 8604
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 22878 5541 22938 19755
rect 25270 9213 25330 34579
rect 26003 33420 26069 33421
rect 26003 33356 26004 33420
rect 26068 33356 26069 33420
rect 26003 33355 26069 33356
rect 25451 17236 25517 17237
rect 25451 17172 25452 17236
rect 25516 17172 25517 17236
rect 25451 17171 25517 17172
rect 25267 9212 25333 9213
rect 25267 9148 25268 9212
rect 25332 9148 25333 9212
rect 25267 9147 25333 9148
rect 22875 5540 22941 5541
rect 22875 5476 22876 5540
rect 22940 5476 22941 5540
rect 22875 5475 22941 5476
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19379 4588 19445 4589
rect 19379 4524 19380 4588
rect 19444 4524 19445 4588
rect 19379 4523 19445 4524
rect 19195 3636 19261 3637
rect 19195 3572 19196 3636
rect 19260 3572 19261 3636
rect 19195 3571 19261 3572
rect 17539 2684 17605 2685
rect 17539 2620 17540 2684
rect 17604 2620 17605 2684
rect 17539 2619 17605 2620
rect 19382 2005 19442 4523
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 25454 2685 25514 17171
rect 26006 10437 26066 33355
rect 26003 10436 26069 10437
rect 26003 10372 26004 10436
rect 26068 10372 26069 10436
rect 26003 10371 26069 10372
rect 27294 9349 27354 43147
rect 28027 18052 28093 18053
rect 28027 17988 28028 18052
rect 28092 17988 28093 18052
rect 28027 17987 28093 17988
rect 28030 16557 28090 17987
rect 28027 16556 28093 16557
rect 28027 16492 28028 16556
rect 28092 16492 28093 16556
rect 28027 16491 28093 16492
rect 28582 9621 28642 61099
rect 28763 60756 28829 60757
rect 28763 60692 28764 60756
rect 28828 60692 28829 60756
rect 28763 60691 28829 60692
rect 28766 17917 28826 60691
rect 28763 17916 28829 17917
rect 28763 17852 28764 17916
rect 28828 17852 28829 17916
rect 28763 17851 28829 17852
rect 28947 16964 29013 16965
rect 28947 16900 28948 16964
rect 29012 16900 29013 16964
rect 28947 16899 29013 16900
rect 28950 13021 29010 16899
rect 29499 16284 29565 16285
rect 29499 16220 29500 16284
rect 29564 16220 29565 16284
rect 29499 16219 29565 16220
rect 28947 13020 29013 13021
rect 28947 12956 28948 13020
rect 29012 12956 29013 13020
rect 28947 12955 29013 12956
rect 28579 9620 28645 9621
rect 28579 9556 28580 9620
rect 28644 9556 28645 9620
rect 28579 9555 28645 9556
rect 28763 9620 28829 9621
rect 28763 9556 28764 9620
rect 28828 9556 28829 9620
rect 28763 9555 28829 9556
rect 27291 9348 27357 9349
rect 27291 9284 27292 9348
rect 27356 9284 27357 9348
rect 27291 9283 27357 9284
rect 28766 8669 28826 9555
rect 28947 9484 29013 9485
rect 28947 9420 28948 9484
rect 29012 9420 29013 9484
rect 28947 9419 29013 9420
rect 28950 8805 29010 9419
rect 28947 8804 29013 8805
rect 28947 8740 28948 8804
rect 29012 8740 29013 8804
rect 28947 8739 29013 8740
rect 28763 8668 28829 8669
rect 28763 8604 28764 8668
rect 28828 8604 28829 8668
rect 28763 8603 28829 8604
rect 29502 5405 29562 16219
rect 30054 10981 30114 61099
rect 34928 60416 35248 61440
rect 34928 60352 34936 60416
rect 35000 60352 35016 60416
rect 35080 60352 35096 60416
rect 35160 60352 35176 60416
rect 35240 60352 35248 60416
rect 34928 59328 35248 60352
rect 50288 60960 50608 61520
rect 50288 60896 50296 60960
rect 50360 60896 50376 60960
rect 50440 60896 50456 60960
rect 50520 60896 50536 60960
rect 50600 60896 50608 60960
rect 40539 60076 40605 60077
rect 40539 60012 40540 60076
rect 40604 60012 40605 60076
rect 40539 60011 40605 60012
rect 34928 59264 34936 59328
rect 35000 59264 35016 59328
rect 35080 59264 35096 59328
rect 35160 59264 35176 59328
rect 35240 59264 35248 59328
rect 34928 58240 35248 59264
rect 39251 58988 39317 58989
rect 39251 58924 39252 58988
rect 39316 58924 39317 58988
rect 39251 58923 39317 58924
rect 34928 58176 34936 58240
rect 35000 58176 35016 58240
rect 35080 58176 35096 58240
rect 35160 58176 35176 58240
rect 35240 58176 35248 58240
rect 34928 57152 35248 58176
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 36307 50284 36373 50285
rect 36307 50220 36308 50284
rect 36372 50220 36373 50284
rect 36307 50219 36373 50220
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 32443 27572 32509 27573
rect 32443 27508 32444 27572
rect 32508 27508 32509 27572
rect 32443 27507 32509 27508
rect 30787 18868 30853 18869
rect 30787 18804 30788 18868
rect 30852 18804 30853 18868
rect 30787 18803 30853 18804
rect 30603 14652 30669 14653
rect 30603 14588 30604 14652
rect 30668 14588 30669 14652
rect 30603 14587 30669 14588
rect 30051 10980 30117 10981
rect 30051 10916 30052 10980
rect 30116 10916 30117 10980
rect 30051 10915 30117 10916
rect 29867 9620 29933 9621
rect 29867 9556 29868 9620
rect 29932 9556 29933 9620
rect 29867 9555 29933 9556
rect 29683 9484 29749 9485
rect 29683 9420 29684 9484
rect 29748 9420 29749 9484
rect 29683 9419 29749 9420
rect 29686 6357 29746 9419
rect 29683 6356 29749 6357
rect 29683 6292 29684 6356
rect 29748 6292 29749 6356
rect 29683 6291 29749 6292
rect 29870 6085 29930 9555
rect 29867 6084 29933 6085
rect 29867 6020 29868 6084
rect 29932 6020 29933 6084
rect 29867 6019 29933 6020
rect 30606 5405 30666 14587
rect 30790 7037 30850 18803
rect 30971 18732 31037 18733
rect 30971 18668 30972 18732
rect 31036 18668 31037 18732
rect 30971 18667 31037 18668
rect 30974 8261 31034 18667
rect 32446 17781 32506 27507
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 32443 17780 32509 17781
rect 32443 17716 32444 17780
rect 32508 17716 32509 17780
rect 32443 17715 32509 17716
rect 31891 14516 31957 14517
rect 31891 14452 31892 14516
rect 31956 14452 31957 14516
rect 31891 14451 31957 14452
rect 31894 8261 31954 14451
rect 30971 8260 31037 8261
rect 30971 8196 30972 8260
rect 31036 8196 31037 8260
rect 30971 8195 31037 8196
rect 31891 8260 31957 8261
rect 31891 8196 31892 8260
rect 31956 8196 31957 8260
rect 31891 8195 31957 8196
rect 30787 7036 30853 7037
rect 30787 6972 30788 7036
rect 30852 6972 30853 7036
rect 30787 6971 30853 6972
rect 29499 5404 29565 5405
rect 29499 5340 29500 5404
rect 29564 5340 29565 5404
rect 29499 5339 29565 5340
rect 30603 5404 30669 5405
rect 30603 5340 30604 5404
rect 30668 5340 30669 5404
rect 30603 5339 30669 5340
rect 32446 3229 32506 17715
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 36310 4045 36370 50219
rect 38147 45388 38213 45389
rect 38147 45324 38148 45388
rect 38212 45324 38213 45388
rect 38147 45323 38213 45324
rect 37411 42668 37477 42669
rect 37411 42604 37412 42668
rect 37476 42604 37477 42668
rect 37411 42603 37477 42604
rect 37414 5813 37474 42603
rect 37411 5812 37477 5813
rect 37411 5748 37412 5812
rect 37476 5748 37477 5812
rect 37411 5747 37477 5748
rect 38150 5133 38210 45323
rect 39067 42124 39133 42125
rect 39067 42060 39068 42124
rect 39132 42060 39133 42124
rect 39067 42059 39133 42060
rect 38699 17372 38765 17373
rect 38699 17308 38700 17372
rect 38764 17308 38765 17372
rect 38699 17307 38765 17308
rect 38702 16285 38762 17307
rect 38699 16284 38765 16285
rect 38699 16220 38700 16284
rect 38764 16220 38765 16284
rect 38699 16219 38765 16220
rect 39070 12613 39130 42059
rect 39067 12612 39133 12613
rect 39067 12548 39068 12612
rect 39132 12548 39133 12612
rect 39067 12547 39133 12548
rect 39254 11117 39314 58923
rect 39251 11116 39317 11117
rect 39251 11052 39252 11116
rect 39316 11052 39317 11116
rect 39251 11051 39317 11052
rect 39987 6900 40053 6901
rect 39987 6836 39988 6900
rect 40052 6836 40053 6900
rect 39987 6835 40053 6836
rect 38147 5132 38213 5133
rect 38147 5068 38148 5132
rect 38212 5068 38213 5132
rect 38147 5067 38213 5068
rect 39990 4045 40050 6835
rect 40542 4045 40602 60011
rect 50288 59872 50608 60896
rect 50288 59808 50296 59872
rect 50360 59808 50376 59872
rect 50440 59808 50456 59872
rect 50520 59808 50536 59872
rect 50600 59808 50608 59872
rect 42563 59396 42629 59397
rect 42563 59332 42564 59396
rect 42628 59332 42629 59396
rect 42563 59331 42629 59332
rect 40723 37772 40789 37773
rect 40723 37708 40724 37772
rect 40788 37708 40789 37772
rect 40723 37707 40789 37708
rect 40726 12477 40786 37707
rect 41091 15876 41157 15877
rect 41091 15812 41092 15876
rect 41156 15812 41157 15876
rect 41091 15811 41157 15812
rect 40723 12476 40789 12477
rect 40723 12412 40724 12476
rect 40788 12412 40789 12476
rect 40723 12411 40789 12412
rect 36307 4044 36373 4045
rect 36307 3980 36308 4044
rect 36372 3980 36373 4044
rect 36307 3979 36373 3980
rect 39987 4044 40053 4045
rect 39987 3980 39988 4044
rect 40052 3980 40053 4044
rect 39987 3979 40053 3980
rect 40539 4044 40605 4045
rect 40539 3980 40540 4044
rect 40604 3980 40605 4044
rect 40539 3979 40605 3980
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 32443 3228 32509 3229
rect 32443 3164 32444 3228
rect 32508 3164 32509 3228
rect 32443 3163 32509 3164
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 25451 2684 25517 2685
rect 25451 2620 25452 2684
rect 25516 2620 25517 2684
rect 25451 2619 25517 2620
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2128 35248 2688
rect 41094 2413 41154 15811
rect 42566 2685 42626 59331
rect 50288 58784 50608 59808
rect 50288 58720 50296 58784
rect 50360 58720 50376 58784
rect 50440 58720 50456 58784
rect 50520 58720 50536 58784
rect 50600 58720 50608 58784
rect 50288 57696 50608 58720
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 43667 57356 43733 57357
rect 43667 57292 43668 57356
rect 43732 57292 43733 57356
rect 43667 57291 43733 57292
rect 42931 48924 42997 48925
rect 42931 48860 42932 48924
rect 42996 48860 42997 48924
rect 42931 48859 42997 48860
rect 42934 16557 42994 48859
rect 42931 16556 42997 16557
rect 42931 16492 42932 16556
rect 42996 16492 42997 16556
rect 42931 16491 42997 16492
rect 43670 3637 43730 57291
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 57283 41580 57349 41581
rect 57283 41516 57284 41580
rect 57348 41516 57349 41580
rect 57283 41515 57349 41516
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 45323 29612 45389 29613
rect 45323 29548 45324 29612
rect 45388 29548 45389 29612
rect 45323 29547 45389 29548
rect 45139 13020 45205 13021
rect 45139 12956 45140 13020
rect 45204 12956 45205 13020
rect 45139 12955 45205 12956
rect 45142 4045 45202 12955
rect 45139 4044 45205 4045
rect 45139 3980 45140 4044
rect 45204 3980 45205 4044
rect 45139 3979 45205 3980
rect 43667 3636 43733 3637
rect 43667 3572 43668 3636
rect 43732 3572 43733 3636
rect 43667 3571 43733 3572
rect 45326 2685 45386 29547
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 57286 19957 57346 41515
rect 57283 19956 57349 19957
rect 57283 19892 57284 19956
rect 57348 19892 57349 19956
rect 57283 19891 57349 19892
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 42563 2684 42629 2685
rect 42563 2620 42564 2684
rect 42628 2620 42629 2684
rect 42563 2619 42629 2620
rect 45323 2684 45389 2685
rect 45323 2620 45324 2684
rect 45388 2620 45389 2684
rect 45323 2619 45389 2620
rect 41091 2412 41157 2413
rect 41091 2348 41092 2412
rect 41156 2348 41157 2412
rect 41091 2347 41157 2348
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
rect 19379 2004 19445 2005
rect 19379 1940 19380 2004
rect 19444 1940 19445 2004
rect 19379 1939 19445 1940
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20240 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform 1 0 21068 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1676037725
transform 1 0 29992 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1676037725
transform 1 0 29348 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1676037725
transform 1 0 30636 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1676037725
transform 1 0 8832 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1676037725
transform 1 0 22356 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1676037725
transform 1 0 22448 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1676037725
transform 1 0 20516 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1676037725
transform 1 0 22356 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1676037725
transform 1 0 41216 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1676037725
transform 1 0 20240 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1676037725
transform 1 0 37904 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1676037725
transform 1 0 26956 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1676037725
transform 1 0 28428 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1676037725
transform 1 0 35236 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1676037725
transform 1 0 32936 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1676037725
transform 1 0 35604 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1676037725
transform 1 0 38364 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1676037725
transform 1 0 17756 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1676037725
transform 1 0 22632 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1676037725
transform 1 0 23460 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1676037725
transform 1 0 2300 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1676037725
transform 1 0 2300 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1676037725
transform 1 0 2300 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1676037725
transform 1 0 2300 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1676037725
transform 1 0 28060 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1676037725
transform 1 0 54004 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1676037725
transform 1 0 23368 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1676037725
transform 1 0 27140 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1676037725
transform 1 0 37628 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1676037725
transform 1 0 36340 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1676037725
transform 1 0 35788 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp 1676037725
transform 1 0 20332 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp 1676037725
transform 1 0 2300 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp 1676037725
transform 1 0 20608 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_37
timestamp 1676037725
transform 1 0 35972 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_38
timestamp 1676037725
transform 1 0 34224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_39
timestamp 1676037725
transform 1 0 34684 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_40
timestamp 1676037725
transform 1 0 35604 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_41
timestamp 1676037725
transform 1 0 35604 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2116 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1676037725
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4140 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38
timestamp 1676037725
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46
timestamp 1676037725
transform 1 0 5336 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1676037725
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1676037725
transform 1 0 6716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66
timestamp 1676037725
transform 1 0 7176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74
timestamp 1676037725
transform 1 0 7912 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1676037725
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89
timestamp 1676037725
transform 1 0 9292 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_94
timestamp 1676037725
transform 1 0 9752 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_102
timestamp 1676037725
transform 1 0 10488 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1676037725
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_118
timestamp 1676037725
transform 1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_128
timestamp 1676037725
transform 1 0 12880 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1676037725
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1676037725
transform 1 0 14536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1676037725
transform 1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1676037725
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_174
timestamp 1676037725
transform 1 0 17112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_184
timestamp 1676037725
transform 1 0 18032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1676037725
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_202
timestamp 1676037725
transform 1 0 19688 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_210
timestamp 1676037725
transform 1 0 20424 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_214
timestamp 1676037725
transform 1 0 20792 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1676037725
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_230
timestamp 1676037725
transform 1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_240
timestamp 1676037725
transform 1 0 23184 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1676037725
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_258
timestamp 1676037725
transform 1 0 24840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_268
timestamp 1676037725
transform 1 0 25760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1676037725
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_286
timestamp 1676037725
transform 1 0 27416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_296
timestamp 1676037725
transform 1 0 28336 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1676037725
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_309 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_315
timestamp 1676037725
transform 1 0 30084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_322
timestamp 1676037725
transform 1 0 30728 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_332
timestamp 1676037725
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_345
timestamp 1676037725
transform 1 0 32844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_355
timestamp 1676037725
transform 1 0 33764 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1676037725
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_373
timestamp 1676037725
transform 1 0 35420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_383
timestamp 1676037725
transform 1 0 36340 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1676037725
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1676037725
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_401
timestamp 1676037725
transform 1 0 37996 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_411
timestamp 1676037725
transform 1 0 38916 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1676037725
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 1676037725
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_429
timestamp 1676037725
transform 1 0 40572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_439
timestamp 1676037725
transform 1 0 41492 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_447
timestamp 1676037725
transform 1 0 42228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_449
timestamp 1676037725
transform 1 0 42412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_460
timestamp 1676037725
transform 1 0 43424 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_468
timestamp 1676037725
transform 1 0 44160 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_477
timestamp 1676037725
transform 1 0 44988 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_483
timestamp 1676037725
transform 1 0 45540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_487
timestamp 1676037725
transform 1 0 45908 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_494
timestamp 1676037725
transform 1 0 46552 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_502
timestamp 1676037725
transform 1 0 47288 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_505
timestamp 1676037725
transform 1 0 47564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_513
timestamp 1676037725
transform 1 0 48300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_523
timestamp 1676037725
transform 1 0 49220 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_531
timestamp 1676037725
transform 1 0 49956 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_533
timestamp 1676037725
transform 1 0 50140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_539
timestamp 1676037725
transform 1 0 50692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_547
timestamp 1676037725
transform 1 0 51428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_555
timestamp 1676037725
transform 1 0 52164 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_559
timestamp 1676037725
transform 1 0 52532 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_561
timestamp 1676037725
transform 1 0 52716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_569
timestamp 1676037725
transform 1 0 53452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_579
timestamp 1676037725
transform 1 0 54372 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_587
timestamp 1676037725
transform 1 0 55108 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_589
timestamp 1676037725
transform 1 0 55292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_597
timestamp 1676037725
transform 1 0 56028 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_605
timestamp 1676037725
transform 1 0 56764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_614
timestamp 1676037725
transform 1 0 57592 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_617
timestamp 1676037725
transform 1 0 57868 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_623
timestamp 1676037725
transform 1 0 58420 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_23
timestamp 1676037725
transform 1 0 3220 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_31
timestamp 1676037725
transform 1 0 3956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_38
timestamp 1676037725
transform 1 0 4600 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_46
timestamp 1676037725
transform 1 0 5336 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1676037725
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_63
timestamp 1676037725
transform 1 0 6900 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_68
timestamp 1676037725
transform 1 0 7360 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_76
timestamp 1676037725
transform 1 0 8096 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_86
timestamp 1676037725
transform 1 0 9016 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_97
timestamp 1676037725
transform 1 0 10028 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_107
timestamp 1676037725
transform 1 0 10948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_123
timestamp 1676037725
transform 1 0 12420 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_131
timestamp 1676037725
transform 1 0 13156 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_141
timestamp 1676037725
transform 1 0 14076 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_151
timestamp 1676037725
transform 1 0 14996 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_162
timestamp 1676037725
transform 1 0 16008 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_177
timestamp 1676037725
transform 1 0 17388 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_187
timestamp 1676037725
transform 1 0 18308 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_197
timestamp 1676037725
transform 1 0 19228 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1676037725
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1676037725
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_229
timestamp 1676037725
transform 1 0 22172 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_236
timestamp 1676037725
transform 1 0 22816 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_249
timestamp 1676037725
transform 1 0 24012 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_258
timestamp 1676037725
transform 1 0 24840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_268
timestamp 1676037725
transform 1 0 25760 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1676037725
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_293
timestamp 1676037725
transform 1 0 28060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_316
timestamp 1676037725
transform 1 0 30176 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_322
timestamp 1676037725
transform 1 0 30728 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1676037725
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1676037725
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_345
timestamp 1676037725
transform 1 0 32844 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_368
timestamp 1676037725
transform 1 0 34960 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_378
timestamp 1676037725
transform 1 0 35880 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1676037725
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_408
timestamp 1676037725
transform 1 0 38640 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_418
timestamp 1676037725
transform 1 0 39560 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_428
timestamp 1676037725
transform 1 0 40480 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_436
timestamp 1676037725
transform 1 0 41216 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_446
timestamp 1676037725
transform 1 0 42136 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_449
timestamp 1676037725
transform 1 0 42412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_465
timestamp 1676037725
transform 1 0 43884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_473
timestamp 1676037725
transform 1 0 44620 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_481
timestamp 1676037725
transform 1 0 45356 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_489
timestamp 1676037725
transform 1 0 46092 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1676037725
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1676037725
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_505
timestamp 1676037725
transform 1 0 47564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_513
timestamp 1676037725
transform 1 0 48300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_523
timestamp 1676037725
transform 1 0 49220 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_533
timestamp 1676037725
transform 1 0 50140 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_541
timestamp 1676037725
transform 1 0 50876 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_549
timestamp 1676037725
transform 1 0 51612 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_557
timestamp 1676037725
transform 1 0 52348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_561
timestamp 1676037725
transform 1 0 52716 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_567
timestamp 1676037725
transform 1 0 53268 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_581
timestamp 1676037725
transform 1 0 54556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_591
timestamp 1676037725
transform 1 0 55476 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_601
timestamp 1676037725
transform 1 0 56396 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_607
timestamp 1676037725
transform 1 0 56948 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_614
timestamp 1676037725
transform 1 0 57592 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_617
timestamp 1676037725
transform 1 0 57868 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_623
timestamp 1676037725
transform 1 0 58420 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_11
timestamp 1676037725
transform 1 0 2116 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_23
timestamp 1676037725
transform 1 0 3220 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_46
timestamp 1676037725
transform 1 0 5336 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_54
timestamp 1676037725
transform 1 0 6072 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_62
timestamp 1676037725
transform 1 0 6808 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_72
timestamp 1676037725
transform 1 0 7728 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1676037725
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_89
timestamp 1676037725
transform 1 0 9292 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_107
timestamp 1676037725
transform 1 0 10948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_113
timestamp 1676037725
transform 1 0 11500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_118
timestamp 1676037725
transform 1 0 11960 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_128
timestamp 1676037725
transform 1 0 12880 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1676037725
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_147
timestamp 1676037725
transform 1 0 14628 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_154
timestamp 1676037725
transform 1 0 15272 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_174
timestamp 1676037725
transform 1 0 17112 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_184
timestamp 1676037725
transform 1 0 18032 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1676037725
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_217
timestamp 1676037725
transform 1 0 21068 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_230
timestamp 1676037725
transform 1 0 22264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1676037725
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_264
timestamp 1676037725
transform 1 0 25392 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_274
timestamp 1676037725
transform 1 0 26312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_285
timestamp 1676037725
transform 1 0 27324 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_298
timestamp 1676037725
transform 1 0 28520 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_306
timestamp 1676037725
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_323
timestamp 1676037725
transform 1 0 30820 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_329
timestamp 1676037725
transform 1 0 31372 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_335
timestamp 1676037725
transform 1 0 31924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_358
timestamp 1676037725
transform 1 0 34040 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_373
timestamp 1676037725
transform 1 0 35420 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_379
timestamp 1676037725
transform 1 0 35972 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_389
timestamp 1676037725
transform 1 0 36892 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_412
timestamp 1676037725
transform 1 0 39008 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_421
timestamp 1676037725
transform 1 0 39836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_438
timestamp 1676037725
transform 1 0 41400 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_446
timestamp 1676037725
transform 1 0 42136 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_452
timestamp 1676037725
transform 1 0 42688 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_470
timestamp 1676037725
transform 1 0 44344 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_477
timestamp 1676037725
transform 1 0 44988 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_483
timestamp 1676037725
transform 1 0 45540 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_491
timestamp 1676037725
transform 1 0 46276 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_503
timestamp 1676037725
transform 1 0 47380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_511
timestamp 1676037725
transform 1 0 48116 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_519
timestamp 1676037725
transform 1 0 48852 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_527
timestamp 1676037725
transform 1 0 49588 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1676037725
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_533
timestamp 1676037725
transform 1 0 50140 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_539
timestamp 1676037725
transform 1 0 50692 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_547
timestamp 1676037725
transform 1 0 51428 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_555
timestamp 1676037725
transform 1 0 52164 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_563
timestamp 1676037725
transform 1 0 52900 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_571
timestamp 1676037725
transform 1 0 53636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_579
timestamp 1676037725
transform 1 0 54372 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1676037725
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_589
timestamp 1676037725
transform 1 0 55292 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_595
timestamp 1676037725
transform 1 0 55844 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_603
timestamp 1676037725
transform 1 0 56580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_622
timestamp 1676037725
transform 1 0 58328 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_11
timestamp 1676037725
transform 1 0 2116 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_23
timestamp 1676037725
transform 1 0 3220 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_35
timestamp 1676037725
transform 1 0 4324 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_47
timestamp 1676037725
transform 1 0 5428 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1676037725
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_63
timestamp 1676037725
transform 1 0 6900 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_71
timestamp 1676037725
transform 1 0 7636 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_92
timestamp 1676037725
transform 1 0 9568 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_102
timestamp 1676037725
transform 1 0 10488 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1676037725
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_119
timestamp 1676037725
transform 1 0 12052 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_129
timestamp 1676037725
transform 1 0 12972 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_139
timestamp 1676037725
transform 1 0 13892 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_157
timestamp 1676037725
transform 1 0 15548 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1676037725
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_178
timestamp 1676037725
transform 1 0 17480 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_188
timestamp 1676037725
transform 1 0 18400 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_201
timestamp 1676037725
transform 1 0 19596 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_221
timestamp 1676037725
transform 1 0 21436 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_237
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_257
timestamp 1676037725
transform 1 0 24748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_267
timestamp 1676037725
transform 1 0 25668 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1676037725
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_301
timestamp 1676037725
transform 1 0 28796 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_309
timestamp 1676037725
transform 1 0 29532 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_317
timestamp 1676037725
transform 1 0 30268 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_325
timestamp 1676037725
transform 1 0 31004 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_329
timestamp 1676037725
transform 1 0 31372 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_334
timestamp 1676037725
transform 1 0 31832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_348
timestamp 1676037725
transform 1 0 33120 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_358
timestamp 1676037725
transform 1 0 34040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_368
timestamp 1676037725
transform 1 0 34960 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_378
timestamp 1676037725
transform 1 0 35880 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_388
timestamp 1676037725
transform 1 0 36800 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_401
timestamp 1676037725
transform 1 0 37996 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_424
timestamp 1676037725
transform 1 0 40112 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_432
timestamp 1676037725
transform 1 0 40848 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_440
timestamp 1676037725
transform 1 0 41584 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_449
timestamp 1676037725
transform 1 0 42412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_466
timestamp 1676037725
transform 1 0 43976 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_474
timestamp 1676037725
transform 1 0 44712 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_482
timestamp 1676037725
transform 1 0 45448 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_490
timestamp 1676037725
transform 1 0 46184 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_498
timestamp 1676037725
transform 1 0 46920 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_505
timestamp 1676037725
transform 1 0 47564 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_511
timestamp 1676037725
transform 1 0 48116 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_516
timestamp 1676037725
transform 1 0 48576 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_528
timestamp 1676037725
transform 1 0 49680 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_540
timestamp 1676037725
transform 1 0 50784 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_552
timestamp 1676037725
transform 1 0 51888 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_558
timestamp 1676037725
transform 1 0 52440 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_561
timestamp 1676037725
transform 1 0 52716 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_567
timestamp 1676037725
transform 1 0 53268 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_575
timestamp 1676037725
transform 1 0 54004 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1676037725
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1676037725
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1676037725
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1676037725
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_617
timestamp 1676037725
transform 1 0 57868 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_623
timestamp 1676037725
transform 1 0 58420 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_61
timestamp 1676037725
transform 1 0 6716 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_66
timestamp 1676037725
transform 1 0 7176 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_74
timestamp 1676037725
transform 1 0 7912 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1676037725
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1676037725
transform 1 0 9476 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_99
timestamp 1676037725
transform 1 0 10212 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_115
timestamp 1676037725
transform 1 0 11684 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_120
timestamp 1676037725
transform 1 0 12144 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_128
timestamp 1676037725
transform 1 0 12880 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1676037725
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_149
timestamp 1676037725
transform 1 0 14812 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_157
timestamp 1676037725
transform 1 0 15548 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_164
timestamp 1676037725
transform 1 0 16192 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_174
timestamp 1676037725
transform 1 0 17112 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_184
timestamp 1676037725
transform 1 0 18032 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1676037725
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_207
timestamp 1676037725
transform 1 0 20148 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_220
timestamp 1676037725
transform 1 0 21344 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_227
timestamp 1676037725
transform 1 0 21988 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_237
timestamp 1676037725
transform 1 0 22908 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1676037725
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_264
timestamp 1676037725
transform 1 0 25392 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_272
timestamp 1676037725
transform 1 0 26128 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_279
timestamp 1676037725
transform 1 0 26772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_290
timestamp 1676037725
transform 1 0 27784 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_296
timestamp 1676037725
transform 1 0 28336 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_306
timestamp 1676037725
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_315
timestamp 1676037725
transform 1 0 30084 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_322
timestamp 1676037725
transform 1 0 30728 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_334
timestamp 1676037725
transform 1 0 31832 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_346
timestamp 1676037725
transform 1 0 32936 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_355
timestamp 1676037725
transform 1 0 33764 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1676037725
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_373
timestamp 1676037725
transform 1 0 35420 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_391
timestamp 1676037725
transform 1 0 37076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_399
timestamp 1676037725
transform 1 0 37812 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_412
timestamp 1676037725
transform 1 0 39008 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_421
timestamp 1676037725
transform 1 0 39836 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_427
timestamp 1676037725
transform 1 0 40388 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_435
timestamp 1676037725
transform 1 0 41124 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_455
timestamp 1676037725
transform 1 0 42964 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_461
timestamp 1676037725
transform 1 0 43516 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_470
timestamp 1676037725
transform 1 0 44344 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_477
timestamp 1676037725
transform 1 0 44988 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_483
timestamp 1676037725
transform 1 0 45540 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_491
timestamp 1676037725
transform 1 0 46276 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_503
timestamp 1676037725
transform 1 0 47380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_515
timestamp 1676037725
transform 1 0 48484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_527
timestamp 1676037725
transform 1 0 49588 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1676037725
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1676037725
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_550
timestamp 1676037725
transform 1 0 51704 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_562
timestamp 1676037725
transform 1 0 52808 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_574
timestamp 1676037725
transform 1 0 53912 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_586
timestamp 1676037725
transform 1 0 55016 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1676037725
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1676037725
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_613
timestamp 1676037725
transform 1 0 57500 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_623
timestamp 1676037725
transform 1 0 58420 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_11
timestamp 1676037725
transform 1 0 2116 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_23
timestamp 1676037725
transform 1 0 3220 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_35
timestamp 1676037725
transform 1 0 4324 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_47
timestamp 1676037725
transform 1 0 5428 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_91
timestamp 1676037725
transform 1 0 9476 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_97
timestamp 1676037725
transform 1 0 10028 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_123
timestamp 1676037725
transform 1 0 12420 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_127
timestamp 1676037725
transform 1 0 12788 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_134
timestamp 1676037725
transform 1 0 13432 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_144
timestamp 1676037725
transform 1 0 14352 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_156
timestamp 1676037725
transform 1 0 15456 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_162
timestamp 1676037725
transform 1 0 16008 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1676037725
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_179
timestamp 1676037725
transform 1 0 17572 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_192
timestamp 1676037725
transform 1 0 18768 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_196
timestamp 1676037725
transform 1 0 19136 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_206
timestamp 1676037725
transform 1 0 20056 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_210
timestamp 1676037725
transform 1 0 20424 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_221
timestamp 1676037725
transform 1 0 21436 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_239
timestamp 1676037725
transform 1 0 23092 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_250
timestamp 1676037725
transform 1 0 24104 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_257
timestamp 1676037725
transform 1 0 24748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_265
timestamp 1676037725
transform 1 0 25484 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_278
timestamp 1676037725
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_289
timestamp 1676037725
transform 1 0 27692 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_302
timestamp 1676037725
transform 1 0 28888 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_310
timestamp 1676037725
transform 1 0 29624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_319
timestamp 1676037725
transform 1 0 30452 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_330
timestamp 1676037725
transform 1 0 31464 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_343
timestamp 1676037725
transform 1 0 32660 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_348
timestamp 1676037725
transform 1 0 33120 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_356
timestamp 1676037725
transform 1 0 33856 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_364
timestamp 1676037725
transform 1 0 34592 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_374
timestamp 1676037725
transform 1 0 35512 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_384
timestamp 1676037725
transform 1 0 36432 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_393
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_400
timestamp 1676037725
transform 1 0 37904 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_408
timestamp 1676037725
transform 1 0 38640 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_414
timestamp 1676037725
transform 1 0 39192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_422
timestamp 1676037725
transform 1 0 39928 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_430
timestamp 1676037725
transform 1 0 40664 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_438
timestamp 1676037725
transform 1 0 41400 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_446
timestamp 1676037725
transform 1 0 42136 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_449
timestamp 1676037725
transform 1 0 42412 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_455
timestamp 1676037725
transform 1 0 42964 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_463
timestamp 1676037725
transform 1 0 43700 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_471
timestamp 1676037725
transform 1 0 44436 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_479
timestamp 1676037725
transform 1 0 45172 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_489
timestamp 1676037725
transform 1 0 46092 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_501
timestamp 1676037725
transform 1 0 47196 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1676037725
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_517
timestamp 1676037725
transform 1 0 48668 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_534
timestamp 1676037725
transform 1 0 50232 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_546
timestamp 1676037725
transform 1 0 51336 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_558
timestamp 1676037725
transform 1 0 52440 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1676037725
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1676037725
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1676037725
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1676037725
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1676037725
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1676037725
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_617
timestamp 1676037725
transform 1 0 57868 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_623
timestamp 1676037725
transform 1 0 58420 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_11
timestamp 1676037725
transform 1 0 2116 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1676037725
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_94
timestamp 1676037725
transform 1 0 9752 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_100
timestamp 1676037725
transform 1 0 10304 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_107
timestamp 1676037725
transform 1 0 10948 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_119
timestamp 1676037725
transform 1 0 12052 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_131
timestamp 1676037725
transform 1 0 13156 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1676037725
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_149
timestamp 1676037725
transform 1 0 14812 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_168
timestamp 1676037725
transform 1 0 16560 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_191
timestamp 1676037725
transform 1 0 18676 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_217
timestamp 1676037725
transform 1 0 21068 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_227
timestamp 1676037725
transform 1 0 21988 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_234
timestamp 1676037725
transform 1 0 22632 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_247
timestamp 1676037725
transform 1 0 23828 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1676037725
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_285
timestamp 1676037725
transform 1 0 27324 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_292
timestamp 1676037725
transform 1 0 27968 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_296
timestamp 1676037725
transform 1 0 28336 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp 1676037725
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_320
timestamp 1676037725
transform 1 0 30544 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_326
timestamp 1676037725
transform 1 0 31096 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_343
timestamp 1676037725
transform 1 0 32660 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_349
timestamp 1676037725
transform 1 0 33212 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_354
timestamp 1676037725
transform 1 0 33672 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_362
timestamp 1676037725
transform 1 0 34408 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_371
timestamp 1676037725
transform 1 0 35236 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_377
timestamp 1676037725
transform 1 0 35788 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_388
timestamp 1676037725
transform 1 0 36800 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_394
timestamp 1676037725
transform 1 0 37352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_400
timestamp 1676037725
transform 1 0 37904 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_404
timestamp 1676037725
transform 1 0 38272 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_407
timestamp 1676037725
transform 1 0 38548 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_418
timestamp 1676037725
transform 1 0 39560 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_421
timestamp 1676037725
transform 1 0 39836 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_427
timestamp 1676037725
transform 1 0 40388 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_435
timestamp 1676037725
transform 1 0 41124 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_441
timestamp 1676037725
transform 1 0 41676 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_453
timestamp 1676037725
transform 1 0 42780 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_465
timestamp 1676037725
transform 1 0 43884 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_473
timestamp 1676037725
transform 1 0 44620 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1676037725
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1676037725
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1676037725
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1676037725
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1676037725
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1676037725
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1676037725
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1676037725
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1676037725
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1676037725
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1676037725
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1676037725
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1676037725
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_601
timestamp 1676037725
transform 1 0 56396 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_613
timestamp 1676037725
transform 1 0 57500 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_623
timestamp 1676037725
transform 1 0 58420 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_11
timestamp 1676037725
transform 1 0 2116 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_23
timestamp 1676037725
transform 1 0 3220 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_35
timestamp 1676037725
transform 1 0 4324 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_47
timestamp 1676037725
transform 1 0 5428 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_94
timestamp 1676037725
transform 1 0 9752 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_106
timestamp 1676037725
transform 1 0 10856 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_133
timestamp 1676037725
transform 1 0 13340 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_138
timestamp 1676037725
transform 1 0 13800 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_148
timestamp 1676037725
transform 1 0 14720 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_152
timestamp 1676037725
transform 1 0 15088 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1676037725
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_177
timestamp 1676037725
transform 1 0 17388 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_189
timestamp 1676037725
transform 1 0 18492 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_197
timestamp 1676037725
transform 1 0 19228 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_216
timestamp 1676037725
transform 1 0 20976 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_235
timestamp 1676037725
transform 1 0 22724 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_241
timestamp 1676037725
transform 1 0 23276 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_262
timestamp 1676037725
transform 1 0 25208 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_275
timestamp 1676037725
transform 1 0 26404 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1676037725
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_290
timestamp 1676037725
transform 1 0 27784 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_302
timestamp 1676037725
transform 1 0 28888 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_330
timestamp 1676037725
transform 1 0 31464 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_349
timestamp 1676037725
transform 1 0 33212 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_359
timestamp 1676037725
transform 1 0 34132 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_369
timestamp 1676037725
transform 1 0 35052 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_379
timestamp 1676037725
transform 1 0 35972 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_387
timestamp 1676037725
transform 1 0 36708 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1676037725
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_399
timestamp 1676037725
transform 1 0 37812 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_411
timestamp 1676037725
transform 1 0 38916 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_423
timestamp 1676037725
transform 1 0 40020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_435
timestamp 1676037725
transform 1 0 41124 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1676037725
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1676037725
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1676037725
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1676037725
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_485
timestamp 1676037725
transform 1 0 45724 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_491
timestamp 1676037725
transform 1 0 46276 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1676037725
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1676037725
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1676037725
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1676037725
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1676037725
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1676037725
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1676037725
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1676037725
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1676037725
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1676037725
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1676037725
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_597
timestamp 1676037725
transform 1 0 56028 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_605
timestamp 1676037725
transform 1 0 56764 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_614
timestamp 1676037725
transform 1 0 57592 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_617
timestamp 1676037725
transform 1 0 57868 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_11
timestamp 1676037725
transform 1 0 2116 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_23
timestamp 1676037725
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1676037725
transform 1 0 9476 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_96
timestamp 1676037725
transform 1 0 9936 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_104
timestamp 1676037725
transform 1 0 10672 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_112
timestamp 1676037725
transform 1 0 11408 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_124
timestamp 1676037725
transform 1 0 12512 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_136
timestamp 1676037725
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_179
timestamp 1676037725
transform 1 0 17572 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_183
timestamp 1676037725
transform 1 0 17940 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1676037725
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_208
timestamp 1676037725
transform 1 0 20240 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_216
timestamp 1676037725
transform 1 0 20976 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_227
timestamp 1676037725
transform 1 0 21988 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_231
timestamp 1676037725
transform 1 0 22356 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_248
timestamp 1676037725
transform 1 0 23920 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_272
timestamp 1676037725
transform 1 0 26128 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_290
timestamp 1676037725
transform 1 0 27784 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_306
timestamp 1676037725
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_325
timestamp 1676037725
transform 1 0 31004 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_338
timestamp 1676037725
transform 1 0 32200 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_347
timestamp 1676037725
transform 1 0 33028 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_355
timestamp 1676037725
transform 1 0 33764 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_362
timestamp 1676037725
transform 1 0 34408 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_376
timestamp 1676037725
transform 1 0 35696 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_387
timestamp 1676037725
transform 1 0 36708 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_399
timestamp 1676037725
transform 1 0 37812 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_411
timestamp 1676037725
transform 1 0 38916 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1676037725
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1676037725
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1676037725
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1676037725
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1676037725
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1676037725
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1676037725
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_477
timestamp 1676037725
transform 1 0 44988 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_482
timestamp 1676037725
transform 1 0 45448 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_495
timestamp 1676037725
transform 1 0 46644 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_507
timestamp 1676037725
transform 1 0 47748 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_519
timestamp 1676037725
transform 1 0 48852 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1676037725
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1676037725
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1676037725
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1676037725
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1676037725
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1676037725
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1676037725
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1676037725
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_601
timestamp 1676037725
transform 1 0 56396 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_605
timestamp 1676037725
transform 1 0 56764 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_622
timestamp 1676037725
transform 1 0 58328 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1676037725
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_89
timestamp 1676037725
transform 1 0 9292 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_95
timestamp 1676037725
transform 1 0 9844 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1676037725
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_119
timestamp 1676037725
transform 1 0 12052 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_129
timestamp 1676037725
transform 1 0 12972 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_141
timestamp 1676037725
transform 1 0 14076 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1676037725
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_184
timestamp 1676037725
transform 1 0 18032 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_198
timestamp 1676037725
transform 1 0 19320 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1676037725
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_237
timestamp 1676037725
transform 1 0 22908 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_248
timestamp 1676037725
transform 1 0 23920 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1676037725
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_285
timestamp 1676037725
transform 1 0 27324 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_295
timestamp 1676037725
transform 1 0 28244 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_319
timestamp 1676037725
transform 1 0 30452 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1676037725
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1676037725
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_346
timestamp 1676037725
transform 1 0 32936 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_375
timestamp 1676037725
transform 1 0 35604 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_379
timestamp 1676037725
transform 1 0 35972 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_390
timestamp 1676037725
transform 1 0 36984 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1676037725
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1676037725
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1676037725
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1676037725
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1676037725
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1676037725
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_461
timestamp 1676037725
transform 1 0 43516 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_469
timestamp 1676037725
transform 1 0 44252 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_473
timestamp 1676037725
transform 1 0 44620 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_493
timestamp 1676037725
transform 1 0 46460 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_501
timestamp 1676037725
transform 1 0 47196 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1676037725
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1676037725
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1676037725
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1676037725
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1676037725
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1676037725
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1676037725
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1676037725
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_585
timestamp 1676037725
transform 1 0 54924 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_597
timestamp 1676037725
transform 1 0 56028 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_610
timestamp 1676037725
transform 1 0 57224 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_617
timestamp 1676037725
transform 1 0 57868 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_622
timestamp 1676037725
transform 1 0 58328 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_11
timestamp 1676037725
transform 1 0 2116 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_23
timestamp 1676037725
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_69
timestamp 1676037725
transform 1 0 7452 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1676037725
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_100
timestamp 1676037725
transform 1 0 10304 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_120
timestamp 1676037725
transform 1 0 12144 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_130
timestamp 1676037725
transform 1 0 13064 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1676037725
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_162
timestamp 1676037725
transform 1 0 16008 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_185
timestamp 1676037725
transform 1 0 18124 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp 1676037725
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_215
timestamp 1676037725
transform 1 0 20884 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_227
timestamp 1676037725
transform 1 0 21988 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_233
timestamp 1676037725
transform 1 0 22540 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_243
timestamp 1676037725
transform 1 0 23460 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1676037725
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_285
timestamp 1676037725
transform 1 0 27324 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_293
timestamp 1676037725
transform 1 0 28060 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_304
timestamp 1676037725
transform 1 0 29072 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_325
timestamp 1676037725
transform 1 0 31004 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_338
timestamp 1676037725
transform 1 0 32200 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_349
timestamp 1676037725
transform 1 0 33212 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_357
timestamp 1676037725
transform 1 0 33948 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_362
timestamp 1676037725
transform 1 0 34408 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_365
timestamp 1676037725
transform 1 0 34684 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_373
timestamp 1676037725
transform 1 0 35420 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_381
timestamp 1676037725
transform 1 0 36156 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_399
timestamp 1676037725
transform 1 0 37812 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_407
timestamp 1676037725
transform 1 0 38548 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_416
timestamp 1676037725
transform 1 0 39376 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1676037725
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1676037725
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_445
timestamp 1676037725
transform 1 0 42044 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_456
timestamp 1676037725
transform 1 0 43056 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_462
timestamp 1676037725
transform 1 0 43608 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_472
timestamp 1676037725
transform 1 0 44528 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_477
timestamp 1676037725
transform 1 0 44988 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_484
timestamp 1676037725
transform 1 0 45632 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_499
timestamp 1676037725
transform 1 0 47012 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_511
timestamp 1676037725
transform 1 0 48116 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_523
timestamp 1676037725
transform 1 0 49220 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1676037725
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1676037725
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1676037725
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1676037725
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1676037725
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1676037725
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1676037725
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_589
timestamp 1676037725
transform 1 0 55292 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_594
timestamp 1676037725
transform 1 0 55752 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_602
timestamp 1676037725
transform 1 0 56488 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_622
timestamp 1676037725
transform 1 0 58328 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_11
timestamp 1676037725
transform 1 0 2116 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_23
timestamp 1676037725
transform 1 0 3220 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_35
timestamp 1676037725
transform 1 0 4324 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_47
timestamp 1676037725
transform 1 0 5428 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_137
timestamp 1676037725
transform 1 0 13708 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_143
timestamp 1676037725
transform 1 0 14260 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_151
timestamp 1676037725
transform 1 0 14996 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_159
timestamp 1676037725
transform 1 0 15732 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1676037725
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_182
timestamp 1676037725
transform 1 0 17848 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1676037725
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1676037725
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1676037725
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_235
timestamp 1676037725
transform 1 0 22724 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_246
timestamp 1676037725
transform 1 0 23736 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_276
timestamp 1676037725
transform 1 0 26496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_299
timestamp 1676037725
transform 1 0 28612 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_307
timestamp 1676037725
transform 1 0 29348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_320
timestamp 1676037725
transform 1 0 30544 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_333
timestamp 1676037725
transform 1 0 31740 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_337
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_343
timestamp 1676037725
transform 1 0 32660 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_352
timestamp 1676037725
transform 1 0 33488 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_364
timestamp 1676037725
transform 1 0 34592 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_381
timestamp 1676037725
transform 1 0 36156 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_390
timestamp 1676037725
transform 1 0 36984 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_393
timestamp 1676037725
transform 1 0 37260 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_404
timestamp 1676037725
transform 1 0 38272 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_412
timestamp 1676037725
transform 1 0 39008 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_430
timestamp 1676037725
transform 1 0 40664 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_442
timestamp 1676037725
transform 1 0 41768 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_449
timestamp 1676037725
transform 1 0 42412 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_462
timestamp 1676037725
transform 1 0 43608 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_468
timestamp 1676037725
transform 1 0 44160 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_476
timestamp 1676037725
transform 1 0 44896 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_486
timestamp 1676037725
transform 1 0 45816 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_498
timestamp 1676037725
transform 1 0 46920 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1676037725
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1676037725
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1676037725
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1676037725
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1676037725
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1676037725
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1676037725
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_573
timestamp 1676037725
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_585
timestamp 1676037725
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_597
timestamp 1676037725
transform 1 0 56028 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_604
timestamp 1676037725
transform 1 0 56672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_614
timestamp 1676037725
transform 1 0 57592 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_617
timestamp 1676037725
transform 1 0 57868 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_11
timestamp 1676037725
transform 1 0 2116 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_23
timestamp 1676037725
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_127
timestamp 1676037725
transform 1 0 12788 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_134
timestamp 1676037725
transform 1 0 13432 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_147
timestamp 1676037725
transform 1 0 14628 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_155
timestamp 1676037725
transform 1 0 15364 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_179
timestamp 1676037725
transform 1 0 17572 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp 1676037725
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_203
timestamp 1676037725
transform 1 0 19780 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_230
timestamp 1676037725
transform 1 0 22264 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_242
timestamp 1676037725
transform 1 0 23368 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1676037725
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_263
timestamp 1676037725
transform 1 0 25300 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_284
timestamp 1676037725
transform 1 0 27232 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_293
timestamp 1676037725
transform 1 0 28060 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_306
timestamp 1676037725
transform 1 0 29256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_313
timestamp 1676037725
transform 1 0 29900 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_325
timestamp 1676037725
transform 1 0 31004 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_336
timestamp 1676037725
transform 1 0 32016 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_344
timestamp 1676037725
transform 1 0 32752 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_351
timestamp 1676037725
transform 1 0 33396 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_361
timestamp 1676037725
transform 1 0 34316 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1676037725
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_386
timestamp 1676037725
transform 1 0 36616 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_406
timestamp 1676037725
transform 1 0 38456 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_414
timestamp 1676037725
transform 1 0 39192 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_421
timestamp 1676037725
transform 1 0 39836 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_427
timestamp 1676037725
transform 1 0 40388 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_434
timestamp 1676037725
transform 1 0 41032 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_446
timestamp 1676037725
transform 1 0 42136 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_458
timestamp 1676037725
transform 1 0 43240 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_462
timestamp 1676037725
transform 1 0 43608 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_474
timestamp 1676037725
transform 1 0 44712 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_477
timestamp 1676037725
transform 1 0 44988 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_485
timestamp 1676037725
transform 1 0 45724 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_492
timestamp 1676037725
transform 1 0 46368 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_504
timestamp 1676037725
transform 1 0 47472 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_516
timestamp 1676037725
transform 1 0 48576 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_528
timestamp 1676037725
transform 1 0 49680 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1676037725
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_545
timestamp 1676037725
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_557
timestamp 1676037725
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_569
timestamp 1676037725
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1676037725
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1676037725
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_589
timestamp 1676037725
transform 1 0 55292 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_597
timestamp 1676037725
transform 1 0 56028 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_602
timestamp 1676037725
transform 1 0 56488 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_622
timestamp 1676037725
transform 1 0 58328 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_11
timestamp 1676037725
transform 1 0 2116 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_23
timestamp 1676037725
transform 1 0 3220 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_35
timestamp 1676037725
transform 1 0 4324 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_47
timestamp 1676037725
transform 1 0 5428 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_89
timestamp 1676037725
transform 1 0 9292 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_101
timestamp 1676037725
transform 1 0 10396 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_109
timestamp 1676037725
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_125
timestamp 1676037725
transform 1 0 12604 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_129
timestamp 1676037725
transform 1 0 12972 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_138
timestamp 1676037725
transform 1 0 13800 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_145
timestamp 1676037725
transform 1 0 14444 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1676037725
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_187
timestamp 1676037725
transform 1 0 18308 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_199
timestamp 1676037725
transform 1 0 19412 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_219
timestamp 1676037725
transform 1 0 21252 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1676037725
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_236
timestamp 1676037725
transform 1 0 22816 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_242
timestamp 1676037725
transform 1 0 23368 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_253
timestamp 1676037725
transform 1 0 24380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_274
timestamp 1676037725
transform 1 0 26312 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_290
timestamp 1676037725
transform 1 0 27784 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_301
timestamp 1676037725
transform 1 0 28796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_312
timestamp 1676037725
transform 1 0 29808 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_320
timestamp 1676037725
transform 1 0 30544 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_330
timestamp 1676037725
transform 1 0 31464 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_337
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_345
timestamp 1676037725
transform 1 0 32844 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_353
timestamp 1676037725
transform 1 0 33580 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_365
timestamp 1676037725
transform 1 0 34684 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_377
timestamp 1676037725
transform 1 0 35788 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_382
timestamp 1676037725
transform 1 0 36248 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_390
timestamp 1676037725
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_393
timestamp 1676037725
transform 1 0 37260 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_403
timestamp 1676037725
transform 1 0 38180 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_415
timestamp 1676037725
transform 1 0 39284 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_427
timestamp 1676037725
transform 1 0 40388 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_439
timestamp 1676037725
transform 1 0 41492 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1676037725
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1676037725
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_461
timestamp 1676037725
transform 1 0 43516 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_471
timestamp 1676037725
transform 1 0 44436 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_495
timestamp 1676037725
transform 1 0 46644 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1676037725
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1676037725
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1676037725
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_529
timestamp 1676037725
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1676037725
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1676037725
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1676037725
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1676037725
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_573
timestamp 1676037725
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_585
timestamp 1676037725
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_597
timestamp 1676037725
transform 1 0 56028 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_605
timestamp 1676037725
transform 1 0 56764 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_610
timestamp 1676037725
transform 1 0 57224 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_617
timestamp 1676037725
transform 1 0 57868 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_11
timestamp 1676037725
transform 1 0 2116 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_23
timestamp 1676037725
transform 1 0 3220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_105
timestamp 1676037725
transform 1 0 10764 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_114
timestamp 1676037725
transform 1 0 11592 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_126
timestamp 1676037725
transform 1 0 12696 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_136
timestamp 1676037725
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_152
timestamp 1676037725
transform 1 0 15088 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_177
timestamp 1676037725
transform 1 0 17388 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1676037725
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_219
timestamp 1676037725
transform 1 0 21252 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_232
timestamp 1676037725
transform 1 0 22448 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_240
timestamp 1676037725
transform 1 0 23184 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1676037725
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_262
timestamp 1676037725
transform 1 0 25208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_286
timestamp 1676037725
transform 1 0 27416 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_295
timestamp 1676037725
transform 1 0 28244 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_306
timestamp 1676037725
transform 1 0 29256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1676037725
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_318
timestamp 1676037725
transform 1 0 30360 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_328
timestamp 1676037725
transform 1 0 31280 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_341
timestamp 1676037725
transform 1 0 32476 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_349
timestamp 1676037725
transform 1 0 33212 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_358
timestamp 1676037725
transform 1 0 34040 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_14_365
timestamp 1676037725
transform 1 0 34684 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_373
timestamp 1676037725
transform 1 0 35420 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_385
timestamp 1676037725
transform 1 0 36524 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_398
timestamp 1676037725
transform 1 0 37720 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_409
timestamp 1676037725
transform 1 0 38732 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_417
timestamp 1676037725
transform 1 0 39468 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1676037725
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1676037725
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1676037725
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_457
timestamp 1676037725
transform 1 0 43148 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_463
timestamp 1676037725
transform 1 0 43700 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_472
timestamp 1676037725
transform 1 0 44528 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_477
timestamp 1676037725
transform 1 0 44988 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_491
timestamp 1676037725
transform 1 0 46276 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_517
timestamp 1676037725
transform 1 0 48668 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_529
timestamp 1676037725
transform 1 0 49772 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1676037725
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_545
timestamp 1676037725
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_557
timestamp 1676037725
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_569
timestamp 1676037725
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1676037725
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1676037725
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_589
timestamp 1676037725
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_601
timestamp 1676037725
transform 1 0 56396 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_613
timestamp 1676037725
transform 1 0 57500 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_623
timestamp 1676037725
transform 1 0 58420 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_11
timestamp 1676037725
transform 1 0 2116 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_23
timestamp 1676037725
transform 1 0 3220 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_35
timestamp 1676037725
transform 1 0 4324 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_47
timestamp 1676037725
transform 1 0 5428 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_81
timestamp 1676037725
transform 1 0 8556 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_86
timestamp 1676037725
transform 1 0 9016 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_95
timestamp 1676037725
transform 1 0 9844 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_107
timestamp 1676037725
transform 1 0 10948 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_121
timestamp 1676037725
transform 1 0 12236 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_127
timestamp 1676037725
transform 1 0 12788 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1676037725
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_149
timestamp 1676037725
transform 1 0 14812 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1676037725
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_184
timestamp 1676037725
transform 1 0 18032 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_188
timestamp 1676037725
transform 1 0 18400 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_198
timestamp 1676037725
transform 1 0 19320 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_218
timestamp 1676037725
transform 1 0 21160 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_237
timestamp 1676037725
transform 1 0 22908 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_245
timestamp 1676037725
transform 1 0 23644 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_256
timestamp 1676037725
transform 1 0 24656 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_272
timestamp 1676037725
transform 1 0 26128 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_292
timestamp 1676037725
transform 1 0 27968 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_319
timestamp 1676037725
transform 1 0 30452 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_325
timestamp 1676037725
transform 1 0 31004 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_334
timestamp 1676037725
transform 1 0 31832 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1676037725
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_349
timestamp 1676037725
transform 1 0 33212 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_362
timestamp 1676037725
transform 1 0 34408 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_372
timestamp 1676037725
transform 1 0 35328 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_384
timestamp 1676037725
transform 1 0 36432 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_393
timestamp 1676037725
transform 1 0 37260 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_401
timestamp 1676037725
transform 1 0 37996 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_413
timestamp 1676037725
transform 1 0 39100 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_425
timestamp 1676037725
transform 1 0 40204 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_433
timestamp 1676037725
transform 1 0 40940 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_444
timestamp 1676037725
transform 1 0 41952 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1676037725
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_461
timestamp 1676037725
transform 1 0 43516 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_467
timestamp 1676037725
transform 1 0 44068 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_488
timestamp 1676037725
transform 1 0 46000 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_500
timestamp 1676037725
transform 1 0 47104 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1676037725
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1676037725
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1676037725
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1676037725
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1676037725
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1676037725
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_561
timestamp 1676037725
transform 1 0 52716 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_572
timestamp 1676037725
transform 1 0 53728 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_584
timestamp 1676037725
transform 1 0 54832 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_596
timestamp 1676037725
transform 1 0 55936 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_608
timestamp 1676037725
transform 1 0 57040 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_612
timestamp 1676037725
transform 1 0 57408 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_617
timestamp 1676037725
transform 1 0 57868 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_11
timestamp 1676037725
transform 1 0 2116 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_23
timestamp 1676037725
transform 1 0 3220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_105
timestamp 1676037725
transform 1 0 10764 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_114
timestamp 1676037725
transform 1 0 11592 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_126
timestamp 1676037725
transform 1 0 12696 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_135
timestamp 1676037725
transform 1 0 13524 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1676037725
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_154
timestamp 1676037725
transform 1 0 15272 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_175
timestamp 1676037725
transform 1 0 17204 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_186
timestamp 1676037725
transform 1 0 18216 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1676037725
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_217
timestamp 1676037725
transform 1 0 21068 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_229
timestamp 1676037725
transform 1 0 22172 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_237
timestamp 1676037725
transform 1 0 22908 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_241
timestamp 1676037725
transform 1 0 23276 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1676037725
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_267
timestamp 1676037725
transform 1 0 25668 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_297
timestamp 1676037725
transform 1 0 28428 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_305
timestamp 1676037725
transform 1 0 29164 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_309
timestamp 1676037725
transform 1 0 29532 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_325
timestamp 1676037725
transform 1 0 31004 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_333
timestamp 1676037725
transform 1 0 31740 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_340
timestamp 1676037725
transform 1 0 32384 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_352
timestamp 1676037725
transform 1 0 33488 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_362
timestamp 1676037725
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_365
timestamp 1676037725
transform 1 0 34684 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_371
timestamp 1676037725
transform 1 0 35236 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_381
timestamp 1676037725
transform 1 0 36156 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_393
timestamp 1676037725
transform 1 0 37260 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_401
timestamp 1676037725
transform 1 0 37996 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_411
timestamp 1676037725
transform 1 0 38916 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1676037725
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_421
timestamp 1676037725
transform 1 0 39836 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_445
timestamp 1676037725
transform 1 0 42044 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_457
timestamp 1676037725
transform 1 0 43148 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_465
timestamp 1676037725
transform 1 0 43884 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_474
timestamp 1676037725
transform 1 0 44712 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1676037725
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_498
timestamp 1676037725
transform 1 0 46920 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_510
timestamp 1676037725
transform 1 0 48024 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_522
timestamp 1676037725
transform 1 0 49128 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_530
timestamp 1676037725
transform 1 0 49864 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1676037725
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1676037725
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_557
timestamp 1676037725
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_569
timestamp 1676037725
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1676037725
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1676037725
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_589
timestamp 1676037725
transform 1 0 55292 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_597
timestamp 1676037725
transform 1 0 56028 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_602
timestamp 1676037725
transform 1 0 56488 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_622
timestamp 1676037725
transform 1 0 58328 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_11
timestamp 1676037725
transform 1 0 2116 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_23
timestamp 1676037725
transform 1 0 3220 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_35
timestamp 1676037725
transform 1 0 4324 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_47
timestamp 1676037725
transform 1 0 5428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1676037725
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_101
timestamp 1676037725
transform 1 0 10396 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1676037725
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_122
timestamp 1676037725
transform 1 0 12328 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_130
timestamp 1676037725
transform 1 0 13064 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_136
timestamp 1676037725
transform 1 0 13616 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_147
timestamp 1676037725
transform 1 0 14628 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_158
timestamp 1676037725
transform 1 0 15640 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_165
timestamp 1676037725
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_187
timestamp 1676037725
transform 1 0 18308 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_191
timestamp 1676037725
transform 1 0 18676 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_197
timestamp 1676037725
transform 1 0 19228 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_214
timestamp 1676037725
transform 1 0 20792 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1676037725
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_232
timestamp 1676037725
transform 1 0 22448 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_244
timestamp 1676037725
transform 1 0 23552 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_250
timestamp 1676037725
transform 1 0 24104 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_258
timestamp 1676037725
transform 1 0 24840 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_267
timestamp 1676037725
transform 1 0 25668 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp 1676037725
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_303
timestamp 1676037725
transform 1 0 28980 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_315
timestamp 1676037725
transform 1 0 30084 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_322
timestamp 1676037725
transform 1 0 30728 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1676037725
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1676037725
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_337
timestamp 1676037725
transform 1 0 32108 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_345
timestamp 1676037725
transform 1 0 32844 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_355
timestamp 1676037725
transform 1 0 33764 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_363
timestamp 1676037725
transform 1 0 34500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_381
timestamp 1676037725
transform 1 0 36156 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_389
timestamp 1676037725
transform 1 0 36892 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1676037725
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_405
timestamp 1676037725
transform 1 0 38364 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1676037725
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1676037725
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1676037725
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_449
timestamp 1676037725
transform 1 0 42412 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_465
timestamp 1676037725
transform 1 0 43884 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_477
timestamp 1676037725
transform 1 0 44988 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_481
timestamp 1676037725
transform 1 0 45356 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_499
timestamp 1676037725
transform 1 0 47012 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1676037725
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1676037725
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1676037725
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1676037725
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1676037725
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1676037725
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1676037725
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_561
timestamp 1676037725
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_573
timestamp 1676037725
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_585
timestamp 1676037725
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_597
timestamp 1676037725
transform 1 0 56028 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_605
timestamp 1676037725
transform 1 0 56764 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_614
timestamp 1676037725
transform 1 0 57592 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_617
timestamp 1676037725
transform 1 0 57868 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_9
timestamp 1676037725
transform 1 0 1932 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_17
timestamp 1676037725
transform 1 0 2668 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_25
timestamp 1676037725
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_101
timestamp 1676037725
transform 1 0 10396 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_107
timestamp 1676037725
transform 1 0 10948 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_122
timestamp 1676037725
transform 1 0 12328 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_130
timestamp 1676037725
transform 1 0 13064 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1676037725
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_145
timestamp 1676037725
transform 1 0 14444 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_155
timestamp 1676037725
transform 1 0 15364 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_187
timestamp 1676037725
transform 1 0 18308 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1676037725
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_204
timestamp 1676037725
transform 1 0 19872 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_232
timestamp 1676037725
transform 1 0 22448 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_236
timestamp 1676037725
transform 1 0 22816 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_247
timestamp 1676037725
transform 1 0 23828 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1676037725
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_260
timestamp 1676037725
transform 1 0 25024 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_273
timestamp 1676037725
transform 1 0 26220 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_281
timestamp 1676037725
transform 1 0 26956 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_298
timestamp 1676037725
transform 1 0 28520 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 1676037725
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_309
timestamp 1676037725
transform 1 0 29532 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_319
timestamp 1676037725
transform 1 0 30452 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_329
timestamp 1676037725
transform 1 0 31372 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_336
timestamp 1676037725
transform 1 0 32016 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_346
timestamp 1676037725
transform 1 0 32936 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_358
timestamp 1676037725
transform 1 0 34040 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_18_365
timestamp 1676037725
transform 1 0 34684 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_371
timestamp 1676037725
transform 1 0 35236 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_379
timestamp 1676037725
transform 1 0 35972 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_402
timestamp 1676037725
transform 1 0 38088 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_414
timestamp 1676037725
transform 1 0 39192 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_421
timestamp 1676037725
transform 1 0 39836 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_431
timestamp 1676037725
transform 1 0 40756 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_449
timestamp 1676037725
transform 1 0 42412 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_461
timestamp 1676037725
transform 1 0 43516 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_473
timestamp 1676037725
transform 1 0 44620 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1676037725
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1676037725
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1676037725
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1676037725
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1676037725
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1676037725
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1676037725
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1676037725
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_557
timestamp 1676037725
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_569
timestamp 1676037725
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1676037725
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1676037725
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_589
timestamp 1676037725
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_601
timestamp 1676037725
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_613
timestamp 1676037725
transform 1 0 57500 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_623
timestamp 1676037725
transform 1 0 58420 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1676037725
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_81
timestamp 1676037725
transform 1 0 8556 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_89
timestamp 1676037725
transform 1 0 9292 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_97
timestamp 1676037725
transform 1 0 10028 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_103
timestamp 1676037725
transform 1 0 10580 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1676037725
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_126
timestamp 1676037725
transform 1 0 12696 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_136
timestamp 1676037725
transform 1 0 13616 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1676037725
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_177
timestamp 1676037725
transform 1 0 17388 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_207
timestamp 1676037725
transform 1 0 20148 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_213
timestamp 1676037725
transform 1 0 20700 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_219
timestamp 1676037725
transform 1 0 21252 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1676037725
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_253
timestamp 1676037725
transform 1 0 24380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1676037725
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1676037725
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_291
timestamp 1676037725
transform 1 0 27876 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_295
timestamp 1676037725
transform 1 0 28244 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_319
timestamp 1676037725
transform 1 0 30452 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_323
timestamp 1676037725
transform 1 0 30820 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_328
timestamp 1676037725
transform 1 0 31280 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_337
timestamp 1676037725
transform 1 0 32108 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_352
timestamp 1676037725
transform 1 0 33488 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_372
timestamp 1676037725
transform 1 0 35328 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_376
timestamp 1676037725
transform 1 0 35696 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_384
timestamp 1676037725
transform 1 0 36432 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1676037725
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1676037725
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1676037725
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1676037725
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_441
timestamp 1676037725
transform 1 0 41676 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_446
timestamp 1676037725
transform 1 0 42136 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_449
timestamp 1676037725
transform 1 0 42412 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_458
timestamp 1676037725
transform 1 0 43240 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_470
timestamp 1676037725
transform 1 0 44344 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_482
timestamp 1676037725
transform 1 0 45448 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_494
timestamp 1676037725
transform 1 0 46552 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_502
timestamp 1676037725
transform 1 0 47288 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1676037725
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1676037725
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_529
timestamp 1676037725
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1676037725
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1676037725
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1676037725
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_561
timestamp 1676037725
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_573
timestamp 1676037725
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_585
timestamp 1676037725
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_597
timestamp 1676037725
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1676037725
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1676037725
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_617
timestamp 1676037725
transform 1 0 57868 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_11
timestamp 1676037725
transform 1 0 2116 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_23
timestamp 1676037725
transform 1 0 3220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1676037725
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_108
timestamp 1676037725
transform 1 0 11040 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1676037725
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_162
timestamp 1676037725
transform 1 0 16008 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1676037725
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_208
timestamp 1676037725
transform 1 0 20240 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_242
timestamp 1676037725
transform 1 0 23368 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_246
timestamp 1676037725
transform 1 0 23736 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1676037725
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_262
timestamp 1676037725
transform 1 0 25208 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_270
timestamp 1676037725
transform 1 0 25944 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_291
timestamp 1676037725
transform 1 0 27876 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_298
timestamp 1676037725
transform 1 0 28520 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_306
timestamp 1676037725
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1676037725
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1676037725
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_333
timestamp 1676037725
transform 1 0 31740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_341
timestamp 1676037725
transform 1 0 32476 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_353
timestamp 1676037725
transform 1 0 33580 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_361
timestamp 1676037725
transform 1 0 34316 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1676037725
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_377
timestamp 1676037725
transform 1 0 35788 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_381
timestamp 1676037725
transform 1 0 36156 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_387
timestamp 1676037725
transform 1 0 36708 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_395
timestamp 1676037725
transform 1 0 37444 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_401
timestamp 1676037725
transform 1 0 37996 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_411
timestamp 1676037725
transform 1 0 38916 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1676037725
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1676037725
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1676037725
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_445
timestamp 1676037725
transform 1 0 42044 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_454
timestamp 1676037725
transform 1 0 42872 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_463
timestamp 1676037725
transform 1 0 43700 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1676037725
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1676037725
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1676037725
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1676037725
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1676037725
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1676037725
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1676037725
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_533
timestamp 1676037725
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_545
timestamp 1676037725
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_557
timestamp 1676037725
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_569
timestamp 1676037725
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1676037725
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1676037725
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_589
timestamp 1676037725
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_601
timestamp 1676037725
transform 1 0 56396 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_613
timestamp 1676037725
transform 1 0 57500 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_623
timestamp 1676037725
transform 1 0 58420 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_11
timestamp 1676037725
transform 1 0 2116 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_23
timestamp 1676037725
transform 1 0 3220 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_35
timestamp 1676037725
transform 1 0 4324 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_47
timestamp 1676037725
transform 1 0 5428 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1676037725
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_81
timestamp 1676037725
transform 1 0 8556 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1676037725
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_132
timestamp 1676037725
transform 1 0 13248 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_136
timestamp 1676037725
transform 1 0 13616 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_163
timestamp 1676037725
transform 1 0 16100 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1676037725
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_188
timestamp 1676037725
transform 1 0 18400 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1676037725
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_241
timestamp 1676037725
transform 1 0 23276 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_245
timestamp 1676037725
transform 1 0 23644 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_256
timestamp 1676037725
transform 1 0 24656 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_268
timestamp 1676037725
transform 1 0 25760 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1676037725
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_288
timestamp 1676037725
transform 1 0 27600 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_300
timestamp 1676037725
transform 1 0 28704 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_315
timestamp 1676037725
transform 1 0 30084 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_333
timestamp 1676037725
transform 1 0 31740 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_337
timestamp 1676037725
transform 1 0 32108 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_348
timestamp 1676037725
transform 1 0 33120 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_360
timestamp 1676037725
transform 1 0 34224 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_372
timestamp 1676037725
transform 1 0 35328 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_384
timestamp 1676037725
transform 1 0 36432 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_393
timestamp 1676037725
transform 1 0 37260 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_399
timestamp 1676037725
transform 1 0 37812 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_408
timestamp 1676037725
transform 1 0 38640 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_415
timestamp 1676037725
transform 1 0 39284 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_427
timestamp 1676037725
transform 1 0 40388 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_446
timestamp 1676037725
transform 1 0 42136 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_449
timestamp 1676037725
transform 1 0 42412 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_455
timestamp 1676037725
transform 1 0 42964 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_475
timestamp 1676037725
transform 1 0 44804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_487
timestamp 1676037725
transform 1 0 45908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_499
timestamp 1676037725
transform 1 0 47012 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1676037725
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1676037725
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_517
timestamp 1676037725
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_529
timestamp 1676037725
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_541
timestamp 1676037725
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1676037725
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1676037725
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_561
timestamp 1676037725
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_573
timestamp 1676037725
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_585
timestamp 1676037725
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_597
timestamp 1676037725
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1676037725
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1676037725
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_617
timestamp 1676037725
transform 1 0 57868 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_11
timestamp 1676037725
transform 1 0 2116 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1676037725
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_108
timestamp 1676037725
transform 1 0 11040 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1676037725
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_162
timestamp 1676037725
transform 1 0 16008 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1676037725
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_201
timestamp 1676037725
transform 1 0 19596 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_219
timestamp 1676037725
transform 1 0 21252 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_249
timestamp 1676037725
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_259
timestamp 1676037725
transform 1 0 24932 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_269
timestamp 1676037725
transform 1 0 25852 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_280
timestamp 1676037725
transform 1 0 26864 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1676037725
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_306
timestamp 1676037725
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1676037725
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_328
timestamp 1676037725
transform 1 0 31280 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_332
timestamp 1676037725
transform 1 0 31648 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_336
timestamp 1676037725
transform 1 0 32016 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_362
timestamp 1676037725
transform 1 0 34408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_365
timestamp 1676037725
transform 1 0 34684 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_376
timestamp 1676037725
transform 1 0 35696 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_388
timestamp 1676037725
transform 1 0 36800 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_397
timestamp 1676037725
transform 1 0 37628 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_418
timestamp 1676037725
transform 1 0 39560 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_421
timestamp 1676037725
transform 1 0 39836 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_440
timestamp 1676037725
transform 1 0 41584 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_452
timestamp 1676037725
transform 1 0 42688 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_474
timestamp 1676037725
transform 1 0 44712 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1676037725
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_489
timestamp 1676037725
transform 1 0 46092 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_495
timestamp 1676037725
transform 1 0 46644 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1676037725
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1676037725
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1676037725
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_533
timestamp 1676037725
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_545
timestamp 1676037725
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_557
timestamp 1676037725
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_569
timestamp 1676037725
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1676037725
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1676037725
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_589
timestamp 1676037725
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_601
timestamp 1676037725
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_613
timestamp 1676037725
transform 1 0 57500 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_623
timestamp 1676037725
transform 1 0 58420 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_11
timestamp 1676037725
transform 1 0 2116 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_23
timestamp 1676037725
transform 1 0 3220 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_35
timestamp 1676037725
transform 1 0 4324 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_47
timestamp 1676037725
transform 1 0 5428 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_81
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1676037725
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_147
timestamp 1676037725
transform 1 0 14628 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1676037725
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_187
timestamp 1676037725
transform 1 0 18308 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_193
timestamp 1676037725
transform 1 0 18860 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1676037725
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_253
timestamp 1676037725
transform 1 0 24380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_274
timestamp 1676037725
transform 1 0 26312 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_281
timestamp 1676037725
transform 1 0 26956 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_289
timestamp 1676037725
transform 1 0 27692 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_299
timestamp 1676037725
transform 1 0 28612 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_303
timestamp 1676037725
transform 1 0 28980 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_308
timestamp 1676037725
transform 1 0 29440 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_321
timestamp 1676037725
transform 1 0 30636 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_333
timestamp 1676037725
transform 1 0 31740 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1676037725
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_358
timestamp 1676037725
transform 1 0 34040 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_378
timestamp 1676037725
transform 1 0 35880 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_390
timestamp 1676037725
transform 1 0 36984 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1676037725
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_405
timestamp 1676037725
transform 1 0 38364 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_414
timestamp 1676037725
transform 1 0 39192 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_426
timestamp 1676037725
transform 1 0 40296 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_438
timestamp 1676037725
transform 1 0 41400 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_446
timestamp 1676037725
transform 1 0 42136 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_449
timestamp 1676037725
transform 1 0 42412 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_453
timestamp 1676037725
transform 1 0 42780 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_460
timestamp 1676037725
transform 1 0 43424 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_472
timestamp 1676037725
transform 1 0 44528 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_484
timestamp 1676037725
transform 1 0 45632 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_496
timestamp 1676037725
transform 1 0 46736 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1676037725
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_517
timestamp 1676037725
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_529
timestamp 1676037725
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_541
timestamp 1676037725
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1676037725
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1676037725
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_561
timestamp 1676037725
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_573
timestamp 1676037725
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_585
timestamp 1676037725
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_597
timestamp 1676037725
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1676037725
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1676037725
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_617
timestamp 1676037725
transform 1 0 57868 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_93
timestamp 1676037725
transform 1 0 9660 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_121
timestamp 1676037725
transform 1 0 12236 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_129
timestamp 1676037725
transform 1 0 12972 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1676037725
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_162
timestamp 1676037725
transform 1 0 16008 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1676037725
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_207
timestamp 1676037725
transform 1 0 20148 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_215
timestamp 1676037725
transform 1 0 20884 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_243
timestamp 1676037725
transform 1 0 23460 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1676037725
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_263
timestamp 1676037725
transform 1 0 25300 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_275
timestamp 1676037725
transform 1 0 26404 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_283
timestamp 1676037725
transform 1 0 27140 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1676037725
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1676037725
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1676037725
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_320
timestamp 1676037725
transform 1 0 30544 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_332
timestamp 1676037725
transform 1 0 31648 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_340
timestamp 1676037725
transform 1 0 32384 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_352
timestamp 1676037725
transform 1 0 33488 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1676037725
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_377
timestamp 1676037725
transform 1 0 35788 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_399
timestamp 1676037725
transform 1 0 37812 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_411
timestamp 1676037725
transform 1 0 38916 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1676037725
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1676037725
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_433
timestamp 1676037725
transform 1 0 40940 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_442
timestamp 1676037725
transform 1 0 41768 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_454
timestamp 1676037725
transform 1 0 42872 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_466
timestamp 1676037725
transform 1 0 43976 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_474
timestamp 1676037725
transform 1 0 44712 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1676037725
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_489
timestamp 1676037725
transform 1 0 46092 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_517
timestamp 1676037725
transform 1 0 48668 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_529
timestamp 1676037725
transform 1 0 49772 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_533
timestamp 1676037725
transform 1 0 50140 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_541
timestamp 1676037725
transform 1 0 50876 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_549
timestamp 1676037725
transform 1 0 51612 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_561
timestamp 1676037725
transform 1 0 52716 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_573
timestamp 1676037725
transform 1 0 53820 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_585
timestamp 1676037725
transform 1 0 54924 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_589
timestamp 1676037725
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_601
timestamp 1676037725
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_613
timestamp 1676037725
transform 1 0 57500 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_623
timestamp 1676037725
transform 1 0 58420 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_11
timestamp 1676037725
transform 1 0 2116 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1676037725
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1676037725
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1676037725
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1676037725
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1676037725
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1676037725
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_93
timestamp 1676037725
transform 1 0 9660 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_101
timestamp 1676037725
transform 1 0 10396 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_109
timestamp 1676037725
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_122
timestamp 1676037725
transform 1 0 12328 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_130
timestamp 1676037725
transform 1 0 13064 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_148
timestamp 1676037725
transform 1 0 14720 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_159
timestamp 1676037725
transform 1 0 15732 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1676037725
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_175
timestamp 1676037725
transform 1 0 17204 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_185
timestamp 1676037725
transform 1 0 18124 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_215
timestamp 1676037725
transform 1 0 20884 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1676037725
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_243
timestamp 1676037725
transform 1 0 23460 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1676037725
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1676037725
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_281
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_293
timestamp 1676037725
transform 1 0 28060 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_313
timestamp 1676037725
transform 1 0 29900 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_322
timestamp 1676037725
transform 1 0 30728 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_334
timestamp 1676037725
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1676037725
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_347
timestamp 1676037725
transform 1 0 33028 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_359
timestamp 1676037725
transform 1 0 34132 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_371
timestamp 1676037725
transform 1 0 35236 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_383
timestamp 1676037725
transform 1 0 36340 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1676037725
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_393
timestamp 1676037725
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_402
timestamp 1676037725
transform 1 0 38088 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_413
timestamp 1676037725
transform 1 0 39100 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_428
timestamp 1676037725
transform 1 0 40480 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_446
timestamp 1676037725
transform 1 0 42136 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_449
timestamp 1676037725
transform 1 0 42412 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_458
timestamp 1676037725
transform 1 0 43240 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_466
timestamp 1676037725
transform 1 0 43976 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_488
timestamp 1676037725
transform 1 0 46000 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_501
timestamp 1676037725
transform 1 0 47196 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_505
timestamp 1676037725
transform 1 0 47564 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_516
timestamp 1676037725
transform 1 0 48576 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_528
timestamp 1676037725
transform 1 0 49680 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_540
timestamp 1676037725
transform 1 0 50784 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_558
timestamp 1676037725
transform 1 0 52440 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_561
timestamp 1676037725
transform 1 0 52716 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_569
timestamp 1676037725
transform 1 0 53452 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_577
timestamp 1676037725
transform 1 0 54188 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_585
timestamp 1676037725
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_597
timestamp 1676037725
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1676037725
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1676037725
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_617
timestamp 1676037725
transform 1 0 57868 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_11
timestamp 1676037725
transform 1 0 2116 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_23
timestamp 1676037725
transform 1 0 3220 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1676037725
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1676037725
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1676037725
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1676037725
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_90
timestamp 1676037725
transform 1 0 9384 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_102
timestamp 1676037725
transform 1 0 10488 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_125
timestamp 1676037725
transform 1 0 12604 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1676037725
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_147
timestamp 1676037725
transform 1 0 14628 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_164
timestamp 1676037725
transform 1 0 16192 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1676037725
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_231
timestamp 1676037725
transform 1 0 22356 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_243
timestamp 1676037725
transform 1 0 23460 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1676037725
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_262
timestamp 1676037725
transform 1 0 25208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_266
timestamp 1676037725
transform 1 0 25576 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_283
timestamp 1676037725
transform 1 0 27140 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_296
timestamp 1676037725
transform 1 0 28336 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_305
timestamp 1676037725
transform 1 0 29164 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1676037725
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1676037725
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_333
timestamp 1676037725
transform 1 0 31740 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_342
timestamp 1676037725
transform 1 0 32568 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_362
timestamp 1676037725
transform 1 0 34408 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1676037725
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_377
timestamp 1676037725
transform 1 0 35788 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_390
timestamp 1676037725
transform 1 0 36984 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_410
timestamp 1676037725
transform 1 0 38824 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_418
timestamp 1676037725
transform 1 0 39560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_421
timestamp 1676037725
transform 1 0 39836 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_427
timestamp 1676037725
transform 1 0 40388 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_435
timestamp 1676037725
transform 1 0 41124 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_446
timestamp 1676037725
transform 1 0 42136 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_458
timestamp 1676037725
transform 1 0 43240 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_470
timestamp 1676037725
transform 1 0 44344 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_477
timestamp 1676037725
transform 1 0 44988 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_496
timestamp 1676037725
transform 1 0 46736 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_508
timestamp 1676037725
transform 1 0 47840 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_520
timestamp 1676037725
transform 1 0 48944 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_533
timestamp 1676037725
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_545
timestamp 1676037725
transform 1 0 51244 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_551
timestamp 1676037725
transform 1 0 51796 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_559
timestamp 1676037725
transform 1 0 52532 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_566
timestamp 1676037725
transform 1 0 53176 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_586
timestamp 1676037725
transform 1 0 55016 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_589
timestamp 1676037725
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_601
timestamp 1676037725
transform 1 0 56396 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_613
timestamp 1676037725
transform 1 0 57500 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_623
timestamp 1676037725
transform 1 0 58420 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_11
timestamp 1676037725
transform 1 0 2116 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1676037725
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1676037725
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1676037725
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1676037725
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_66
timestamp 1676037725
transform 1 0 7176 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_74
timestamp 1676037725
transform 1 0 7912 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_96
timestamp 1676037725
transform 1 0 9936 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_108
timestamp 1676037725
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_121
timestamp 1676037725
transform 1 0 12236 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_150
timestamp 1676037725
transform 1 0 14904 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_158
timestamp 1676037725
transform 1 0 15640 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1676037725
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_176
timestamp 1676037725
transform 1 0 17296 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_206
timestamp 1676037725
transform 1 0 20056 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_211
timestamp 1676037725
transform 1 0 20516 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1676037725
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_253
timestamp 1676037725
transform 1 0 24380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_266
timestamp 1676037725
transform 1 0 25576 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_277
timestamp 1676037725
transform 1 0 26588 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_285
timestamp 1676037725
transform 1 0 27324 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_294
timestamp 1676037725
transform 1 0 28152 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_306
timestamp 1676037725
transform 1 0 29256 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_310
timestamp 1676037725
transform 1 0 29624 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_320
timestamp 1676037725
transform 1 0 30544 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_332
timestamp 1676037725
transform 1 0 31648 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1676037725
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_346
timestamp 1676037725
transform 1 0 32936 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_371
timestamp 1676037725
transform 1 0 35236 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_383
timestamp 1676037725
transform 1 0 36340 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1676037725
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_393
timestamp 1676037725
transform 1 0 37260 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_401
timestamp 1676037725
transform 1 0 37996 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_412
timestamp 1676037725
transform 1 0 39008 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_424
timestamp 1676037725
transform 1 0 40112 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_428
timestamp 1676037725
transform 1 0 40480 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_438
timestamp 1676037725
transform 1 0 41400 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_446
timestamp 1676037725
transform 1 0 42136 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1676037725
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1676037725
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1676037725
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1676037725
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1676037725
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1676037725
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1676037725
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_517
timestamp 1676037725
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_529
timestamp 1676037725
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_541
timestamp 1676037725
transform 1 0 50876 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_545
timestamp 1676037725
transform 1 0 51244 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_551
timestamp 1676037725
transform 1 0 51796 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1676037725
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_561
timestamp 1676037725
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_573
timestamp 1676037725
transform 1 0 53820 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_579
timestamp 1676037725
transform 1 0 54372 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_590
timestamp 1676037725
transform 1 0 55384 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_599
timestamp 1676037725
transform 1 0 56212 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_607
timestamp 1676037725
transform 1 0 56948 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_614
timestamp 1676037725
transform 1 0 57592 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_617
timestamp 1676037725
transform 1 0 57868 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_11
timestamp 1676037725
transform 1 0 2116 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_23
timestamp 1676037725
transform 1 0 3220 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_53
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_61
timestamp 1676037725
transform 1 0 6716 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_71
timestamp 1676037725
transform 1 0 7636 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1676037725
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_94
timestamp 1676037725
transform 1 0 9752 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_124
timestamp 1676037725
transform 1 0 12512 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_134
timestamp 1676037725
transform 1 0 13432 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_150
timestamp 1676037725
transform 1 0 14904 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_159
timestamp 1676037725
transform 1 0 15732 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1676037725
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1676037725
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_202
timestamp 1676037725
transform 1 0 19688 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_232
timestamp 1676037725
transform 1 0 22448 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1676037725
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1676037725
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_264
timestamp 1676037725
transform 1 0 25392 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_288
timestamp 1676037725
transform 1 0 27600 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_292
timestamp 1676037725
transform 1 0 27968 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1676037725
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1676037725
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_309
timestamp 1676037725
transform 1 0 29532 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_315
timestamp 1676037725
transform 1 0 30084 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_325
timestamp 1676037725
transform 1 0 31004 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_335
timestamp 1676037725
transform 1 0 31924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_344
timestamp 1676037725
transform 1 0 32752 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_348
timestamp 1676037725
transform 1 0 33120 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_359
timestamp 1676037725
transform 1 0 34132 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1676037725
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_365
timestamp 1676037725
transform 1 0 34684 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_372
timestamp 1676037725
transform 1 0 35328 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_384
timestamp 1676037725
transform 1 0 36432 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_396
timestamp 1676037725
transform 1 0 37536 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_408
timestamp 1676037725
transform 1 0 38640 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_418
timestamp 1676037725
transform 1 0 39560 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_421
timestamp 1676037725
transform 1 0 39836 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_425
timestamp 1676037725
transform 1 0 40204 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_442
timestamp 1676037725
transform 1 0 41768 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_454
timestamp 1676037725
transform 1 0 42872 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_466
timestamp 1676037725
transform 1 0 43976 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_474
timestamp 1676037725
transform 1 0 44712 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1676037725
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1676037725
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_501
timestamp 1676037725
transform 1 0 47196 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_507
timestamp 1676037725
transform 1 0 47748 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_515
timestamp 1676037725
transform 1 0 48484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_527
timestamp 1676037725
transform 1 0 49588 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1676037725
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_533
timestamp 1676037725
transform 1 0 50140 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_543
timestamp 1676037725
transform 1 0 51060 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_563
timestamp 1676037725
transform 1 0 52900 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_575
timestamp 1676037725
transform 1 0 54004 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1676037725
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_589
timestamp 1676037725
transform 1 0 55292 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_597
timestamp 1676037725
transform 1 0 56028 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_605
timestamp 1676037725
transform 1 0 56764 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_622
timestamp 1676037725
transform 1 0 58328 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1676037725
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1676037725
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1676037725
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1676037725
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1676037725
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_76
timestamp 1676037725
transform 1 0 8096 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_80
timestamp 1676037725
transform 1 0 8464 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_107
timestamp 1676037725
transform 1 0 10948 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1676037725
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_123
timestamp 1676037725
transform 1 0 12420 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_153
timestamp 1676037725
transform 1 0 15180 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1676037725
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_173
timestamp 1676037725
transform 1 0 17020 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_191
timestamp 1676037725
transform 1 0 18676 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_195
timestamp 1676037725
transform 1 0 19044 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1676037725
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_236
timestamp 1676037725
transform 1 0 22816 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_242
timestamp 1676037725
transform 1 0 23368 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_248
timestamp 1676037725
transform 1 0 23920 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1676037725
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_281
timestamp 1676037725
transform 1 0 26956 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_304
timestamp 1676037725
transform 1 0 29072 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_316
timestamp 1676037725
transform 1 0 30176 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_322
timestamp 1676037725
transform 1 0 30728 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_332
timestamp 1676037725
transform 1 0 31648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_363
timestamp 1676037725
transform 1 0 34500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_367
timestamp 1676037725
transform 1 0 34868 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_378
timestamp 1676037725
transform 1 0 35880 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_390
timestamp 1676037725
transform 1 0 36984 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1676037725
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_405
timestamp 1676037725
transform 1 0 38364 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_428
timestamp 1676037725
transform 1 0 40480 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_436
timestamp 1676037725
transform 1 0 41216 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_446
timestamp 1676037725
transform 1 0 42136 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_449
timestamp 1676037725
transform 1 0 42412 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_459
timestamp 1676037725
transform 1 0 43332 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_471
timestamp 1676037725
transform 1 0 44436 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_483
timestamp 1676037725
transform 1 0 45540 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_493
timestamp 1676037725
transform 1 0 46460 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_501
timestamp 1676037725
transform 1 0 47196 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_505
timestamp 1676037725
transform 1 0 47564 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_513
timestamp 1676037725
transform 1 0 48300 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_532
timestamp 1676037725
transform 1 0 50048 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_544
timestamp 1676037725
transform 1 0 51152 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_556
timestamp 1676037725
transform 1 0 52256 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_561
timestamp 1676037725
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_573
timestamp 1676037725
transform 1 0 53820 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_577
timestamp 1676037725
transform 1 0 54188 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_586
timestamp 1676037725
transform 1 0 55016 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_29_610
timestamp 1676037725
transform 1 0 57224 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_617
timestamp 1676037725
transform 1 0 57868 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_11
timestamp 1676037725
transform 1 0 2116 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1676037725
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1676037725
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_53
timestamp 1676037725
transform 1 0 5980 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1676037725
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_104
timestamp 1676037725
transform 1 0 10672 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1676037725
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_162
timestamp 1676037725
transform 1 0 16008 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1676037725
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1676037725
transform 1 0 20884 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1676037725
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1676037725
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_258
timestamp 1676037725
transform 1 0 24840 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_262
timestamp 1676037725
transform 1 0 25208 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_272
timestamp 1676037725
transform 1 0 26128 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_302
timestamp 1676037725
transform 1 0 28888 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_309
timestamp 1676037725
transform 1 0 29532 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_334
timestamp 1676037725
transform 1 0 31832 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_343
timestamp 1676037725
transform 1 0 32660 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_361
timestamp 1676037725
transform 1 0 34316 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_365
timestamp 1676037725
transform 1 0 34684 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_373
timestamp 1676037725
transform 1 0 35420 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_377
timestamp 1676037725
transform 1 0 35788 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_381
timestamp 1676037725
transform 1 0 36156 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_385
timestamp 1676037725
transform 1 0 36524 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_397
timestamp 1676037725
transform 1 0 37628 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_405
timestamp 1676037725
transform 1 0 38364 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1676037725
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1676037725
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_421
timestamp 1676037725
transform 1 0 39836 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_438
timestamp 1676037725
transform 1 0 41400 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_450
timestamp 1676037725
transform 1 0 42504 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_460
timestamp 1676037725
transform 1 0 43424 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_472
timestamp 1676037725
transform 1 0 44528 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_477
timestamp 1676037725
transform 1 0 44988 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_484
timestamp 1676037725
transform 1 0 45632 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_495
timestamp 1676037725
transform 1 0 46644 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_505
timestamp 1676037725
transform 1 0 47564 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_518
timestamp 1676037725
transform 1 0 48760 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_530
timestamp 1676037725
transform 1 0 49864 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_533
timestamp 1676037725
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_545
timestamp 1676037725
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_557
timestamp 1676037725
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_569
timestamp 1676037725
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1676037725
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1676037725
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_589
timestamp 1676037725
transform 1 0 55292 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_596
timestamp 1676037725
transform 1 0 55936 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_604
timestamp 1676037725
transform 1 0 56672 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_613
timestamp 1676037725
transform 1 0 57500 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_623
timestamp 1676037725
transform 1 0 58420 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_11
timestamp 1676037725
transform 1 0 2116 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1676037725
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1676037725
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1676037725
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1676037725
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1676037725
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_61
timestamp 1676037725
transform 1 0 6716 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_79
timestamp 1676037725
transform 1 0 8372 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_83
timestamp 1676037725
transform 1 0 8740 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1676037725
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_136
timestamp 1676037725
transform 1 0 13616 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1676037725
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_190
timestamp 1676037725
transform 1 0 18584 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1676037725
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_248
timestamp 1676037725
transform 1 0 23920 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1676037725
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1676037725
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_309
timestamp 1676037725
transform 1 0 29532 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_334
timestamp 1676037725
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_337
timestamp 1676037725
transform 1 0 32108 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_358
timestamp 1676037725
transform 1 0 34040 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_362
timestamp 1676037725
transform 1 0 34408 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_373
timestamp 1676037725
transform 1 0 35420 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_377
timestamp 1676037725
transform 1 0 35788 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_388
timestamp 1676037725
transform 1 0 36800 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1676037725
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1676037725
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_417
timestamp 1676037725
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1676037725
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_446
timestamp 1676037725
transform 1 0 42136 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_449
timestamp 1676037725
transform 1 0 42412 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_459
timestamp 1676037725
transform 1 0 43332 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_469
timestamp 1676037725
transform 1 0 44252 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_498
timestamp 1676037725
transform 1 0 46920 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_505
timestamp 1676037725
transform 1 0 47564 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_513
timestamp 1676037725
transform 1 0 48300 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_525
timestamp 1676037725
transform 1 0 49404 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_531
timestamp 1676037725
transform 1 0 49956 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_537
timestamp 1676037725
transform 1 0 50508 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_548
timestamp 1676037725
transform 1 0 51520 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_557
timestamp 1676037725
transform 1 0 52348 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_561
timestamp 1676037725
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_573
timestamp 1676037725
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_585
timestamp 1676037725
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_597
timestamp 1676037725
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1676037725
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1676037725
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_617
timestamp 1676037725
transform 1 0 57868 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_11
timestamp 1676037725
transform 1 0 2116 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_23
timestamp 1676037725
transform 1 0 3220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1676037725
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_53
timestamp 1676037725
transform 1 0 5980 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1676037725
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_93
timestamp 1676037725
transform 1 0 9660 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_97
timestamp 1676037725
transform 1 0 10028 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_105
timestamp 1676037725
transform 1 0 10764 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_111
timestamp 1676037725
transform 1 0 11316 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1676037725
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_164
timestamp 1676037725
transform 1 0 16192 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1676037725
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_216
timestamp 1676037725
transform 1 0 20976 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_248
timestamp 1676037725
transform 1 0 23920 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_267
timestamp 1676037725
transform 1 0 25668 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_273
timestamp 1676037725
transform 1 0 26220 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_300
timestamp 1676037725
transform 1 0 28704 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1676037725
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_316
timestamp 1676037725
transform 1 0 30176 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_320
timestamp 1676037725
transform 1 0 30544 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_347
timestamp 1676037725
transform 1 0 33028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_359
timestamp 1676037725
transform 1 0 34132 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1676037725
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_365
timestamp 1676037725
transform 1 0 34684 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_373
timestamp 1676037725
transform 1 0 35420 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_394
timestamp 1676037725
transform 1 0 37352 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_407
timestamp 1676037725
transform 1 0 38548 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1676037725
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_421
timestamp 1676037725
transform 1 0 39836 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_425
timestamp 1676037725
transform 1 0 40204 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_431
timestamp 1676037725
transform 1 0 40756 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_452
timestamp 1676037725
transform 1 0 42688 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_472
timestamp 1676037725
transform 1 0 44528 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_477
timestamp 1676037725
transform 1 0 44988 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_485
timestamp 1676037725
transform 1 0 45724 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_506
timestamp 1676037725
transform 1 0 47656 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_515
timestamp 1676037725
transform 1 0 48484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_527
timestamp 1676037725
transform 1 0 49588 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1676037725
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_533
timestamp 1676037725
transform 1 0 50140 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_542
timestamp 1676037725
transform 1 0 50968 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_546
timestamp 1676037725
transform 1 0 51336 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_564
timestamp 1676037725
transform 1 0 52992 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_572
timestamp 1676037725
transform 1 0 53728 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_580
timestamp 1676037725
transform 1 0 54464 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_589
timestamp 1676037725
transform 1 0 55292 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_598
timestamp 1676037725
transform 1 0 56120 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_602
timestamp 1676037725
transform 1 0 56488 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_619
timestamp 1676037725
transform 1 0 58052 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_11
timestamp 1676037725
transform 1 0 2116 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_23
timestamp 1676037725
transform 1 0 3220 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_35
timestamp 1676037725
transform 1 0 4324 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_47
timestamp 1676037725
transform 1 0 5428 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1676037725
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_69
timestamp 1676037725
transform 1 0 7452 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_33_101
timestamp 1676037725
transform 1 0 10396 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1676037725
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_119
timestamp 1676037725
transform 1 0 12052 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_136
timestamp 1676037725
transform 1 0 13616 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1676037725
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_185
timestamp 1676037725
transform 1 0 18124 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_215
timestamp 1676037725
transform 1 0 20884 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1676037725
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_243
timestamp 1676037725
transform 1 0 23460 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_251
timestamp 1676037725
transform 1 0 24196 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1676037725
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1676037725
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_300
timestamp 1676037725
transform 1 0 28704 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_334
timestamp 1676037725
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1676037725
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_349
timestamp 1676037725
transform 1 0 33212 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_355
timestamp 1676037725
transform 1 0 33764 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_367
timestamp 1676037725
transform 1 0 34868 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_389
timestamp 1676037725
transform 1 0 36892 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_393
timestamp 1676037725
transform 1 0 37260 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_400
timestamp 1676037725
transform 1 0 37904 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_404
timestamp 1676037725
transform 1 0 38272 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_424
timestamp 1676037725
transform 1 0 40112 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1676037725
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1676037725
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_449
timestamp 1676037725
transform 1 0 42412 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_468
timestamp 1676037725
transform 1 0 44160 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_480
timestamp 1676037725
transform 1 0 45264 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_486
timestamp 1676037725
transform 1 0 45816 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_493
timestamp 1676037725
transform 1 0 46460 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_502
timestamp 1676037725
transform 1 0 47288 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_505
timestamp 1676037725
transform 1 0 47564 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_33_528
timestamp 1676037725
transform 1 0 49680 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_551
timestamp 1676037725
transform 1 0 51796 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1676037725
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_561
timestamp 1676037725
transform 1 0 52716 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_581
timestamp 1676037725
transform 1 0 54556 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_601
timestamp 1676037725
transform 1 0 56396 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_613
timestamp 1676037725
transform 1 0 57500 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_617
timestamp 1676037725
transform 1 0 57868 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1676037725
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1676037725
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1676037725
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1676037725
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1676037725
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1676037725
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1676037725
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1676037725
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_109
timestamp 1676037725
transform 1 0 11132 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_113
timestamp 1676037725
transform 1 0 11500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_121
timestamp 1676037725
transform 1 0 12236 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1676037725
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1676037725
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_153
timestamp 1676037725
transform 1 0 15180 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_157
timestamp 1676037725
transform 1 0 15548 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_164
timestamp 1676037725
transform 1 0 16192 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1676037725
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_207
timestamp 1676037725
transform 1 0 20148 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_241
timestamp 1676037725
transform 1 0 23276 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1676037725
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_271
timestamp 1676037725
transform 1 0 26036 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_279
timestamp 1676037725
transform 1 0 26772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_283
timestamp 1676037725
transform 1 0 27140 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_294
timestamp 1676037725
transform 1 0 28152 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_303
timestamp 1676037725
transform 1 0 28980 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1676037725
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_309
timestamp 1676037725
transform 1 0 29532 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_317
timestamp 1676037725
transform 1 0 30268 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_330
timestamp 1676037725
transform 1 0 31464 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_342
timestamp 1676037725
transform 1 0 32568 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_354
timestamp 1676037725
transform 1 0 33672 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 1676037725
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_365
timestamp 1676037725
transform 1 0 34684 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_393
timestamp 1676037725
transform 1 0 37260 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_401
timestamp 1676037725
transform 1 0 37996 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_409
timestamp 1676037725
transform 1 0 38732 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_417
timestamp 1676037725
transform 1 0 39468 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1676037725
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_433
timestamp 1676037725
transform 1 0 40940 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_448
timestamp 1676037725
transform 1 0 42320 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_457
timestamp 1676037725
transform 1 0 43148 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_466
timestamp 1676037725
transform 1 0 43976 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_474
timestamp 1676037725
transform 1 0 44712 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1676037725
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1676037725
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_501
timestamp 1676037725
transform 1 0 47196 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_511
timestamp 1676037725
transform 1 0 48116 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_523
timestamp 1676037725
transform 1 0 49220 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1676037725
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_533
timestamp 1676037725
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_545
timestamp 1676037725
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_557
timestamp 1676037725
transform 1 0 52348 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_568
timestamp 1676037725
transform 1 0 53360 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_577
timestamp 1676037725
transform 1 0 54188 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_586
timestamp 1676037725
transform 1 0 55016 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_589
timestamp 1676037725
transform 1 0 55292 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_597
timestamp 1676037725
transform 1 0 56028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_609
timestamp 1676037725
transform 1 0 57132 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_623
timestamp 1676037725
transform 1 0 58420 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_9
timestamp 1676037725
transform 1 0 1932 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_21
timestamp 1676037725
transform 1 0 3036 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_33
timestamp 1676037725
transform 1 0 4140 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_45
timestamp 1676037725
transform 1 0 5244 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1676037725
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1676037725
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1676037725
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1676037725
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1676037725
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1676037725
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_120
timestamp 1676037725
transform 1 0 12144 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_126
timestamp 1676037725
transform 1 0 12696 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_134
timestamp 1676037725
transform 1 0 13432 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_146
timestamp 1676037725
transform 1 0 14536 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_152
timestamp 1676037725
transform 1 0 15088 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_156
timestamp 1676037725
transform 1 0 15456 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_162
timestamp 1676037725
transform 1 0 16008 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1676037725
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_188
timestamp 1676037725
transform 1 0 18400 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_218
timestamp 1676037725
transform 1 0 21160 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_236
timestamp 1676037725
transform 1 0 22816 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_270
timestamp 1676037725
transform 1 0 25944 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1676037725
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_281
timestamp 1676037725
transform 1 0 26956 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_285
timestamp 1676037725
transform 1 0 27324 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_295
timestamp 1676037725
transform 1 0 28244 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_325
timestamp 1676037725
transform 1 0 31004 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_333
timestamp 1676037725
transform 1 0 31740 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1676037725
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1676037725
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_361
timestamp 1676037725
transform 1 0 34316 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_369
timestamp 1676037725
transform 1 0 35052 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_373
timestamp 1676037725
transform 1 0 35420 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_384
timestamp 1676037725
transform 1 0 36432 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_35_393
timestamp 1676037725
transform 1 0 37260 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_399
timestamp 1676037725
transform 1 0 37812 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_402
timestamp 1676037725
transform 1 0 38088 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_413
timestamp 1676037725
transform 1 0 39100 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_425
timestamp 1676037725
transform 1 0 40204 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_437
timestamp 1676037725
transform 1 0 41308 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_445
timestamp 1676037725
transform 1 0 42044 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1676037725
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1676037725
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1676037725
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1676037725
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1676037725
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1676037725
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_505
timestamp 1676037725
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_517
timestamp 1676037725
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_529
timestamp 1676037725
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_541
timestamp 1676037725
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1676037725
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1676037725
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_561
timestamp 1676037725
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_573
timestamp 1676037725
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_585
timestamp 1676037725
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_597
timestamp 1676037725
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1676037725
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1676037725
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_617
timestamp 1676037725
transform 1 0 57868 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_623
timestamp 1676037725
transform 1 0 58420 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_11
timestamp 1676037725
transform 1 0 2116 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_23
timestamp 1676037725
transform 1 0 3220 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1676037725
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1676037725
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1676037725
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1676037725
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1676037725
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1676037725
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_96
timestamp 1676037725
transform 1 0 9936 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_108
timestamp 1676037725
transform 1 0 11040 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_120
timestamp 1676037725
transform 1 0 12144 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_132
timestamp 1676037725
transform 1 0 13248 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1676037725
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_165
timestamp 1676037725
transform 1 0 16284 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1676037725
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_208
timestamp 1676037725
transform 1 0 20240 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1676037725
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1676037725
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1676037725
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1676037725
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_265
timestamp 1676037725
transform 1 0 25484 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_275
timestamp 1676037725
transform 1 0 26404 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_287
timestamp 1676037725
transform 1 0 27508 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_299
timestamp 1676037725
transform 1 0 28612 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1676037725
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1676037725
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1676037725
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1676037725
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1676037725
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1676037725
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1676037725
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1676037725
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1676037725
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1676037725
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_401
timestamp 1676037725
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1676037725
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1676037725
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1676037725
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1676037725
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1676037725
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1676037725
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1676037725
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1676037725
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1676037725
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1676037725
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1676037725
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_513
timestamp 1676037725
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1676037725
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1676037725
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_533
timestamp 1676037725
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_545
timestamp 1676037725
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_557
timestamp 1676037725
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_569
timestamp 1676037725
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1676037725
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1676037725
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_589
timestamp 1676037725
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_601
timestamp 1676037725
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_613
timestamp 1676037725
transform 1 0 57500 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_623
timestamp 1676037725
transform 1 0 58420 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_11
timestamp 1676037725
transform 1 0 2116 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_23
timestamp 1676037725
transform 1 0 3220 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_35
timestamp 1676037725
transform 1 0 4324 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_47
timestamp 1676037725
transform 1 0 5428 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1676037725
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1676037725
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1676037725
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1676037725
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1676037725
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1676037725
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1676037725
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1676037725
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1676037725
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1676037725
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1676037725
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_178
timestamp 1676037725
transform 1 0 17480 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_190
timestamp 1676037725
transform 1 0 18584 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_198
timestamp 1676037725
transform 1 0 19320 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_204
timestamp 1676037725
transform 1 0 19872 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_216
timestamp 1676037725
transform 1 0 20976 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1676037725
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1676037725
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_261
timestamp 1676037725
transform 1 0 25116 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_267
timestamp 1676037725
transform 1 0 25668 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1676037725
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1676037725
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1676037725
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1676037725
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1676037725
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1676037725
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1676037725
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1676037725
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1676037725
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1676037725
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1676037725
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1676037725
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1676037725
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1676037725
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1676037725
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_405
timestamp 1676037725
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_417
timestamp 1676037725
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_429
timestamp 1676037725
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1676037725
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1676037725
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1676037725
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1676037725
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1676037725
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1676037725
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1676037725
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1676037725
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1676037725
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_517
timestamp 1676037725
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_529
timestamp 1676037725
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_541
timestamp 1676037725
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1676037725
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1676037725
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_561
timestamp 1676037725
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_573
timestamp 1676037725
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_585
timestamp 1676037725
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_597
timestamp 1676037725
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1676037725
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1676037725
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_617
timestamp 1676037725
transform 1 0 57868 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_623
timestamp 1676037725
transform 1 0 58420 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_11
timestamp 1676037725
transform 1 0 2116 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_23
timestamp 1676037725
transform 1 0 3220 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1676037725
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1676037725
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1676037725
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1676037725
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1676037725
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1676037725
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_97
timestamp 1676037725
transform 1 0 10028 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_105
timestamp 1676037725
transform 1 0 10764 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_111
timestamp 1676037725
transform 1 0 11316 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_117
timestamp 1676037725
transform 1 0 11868 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_123
timestamp 1676037725
transform 1 0 12420 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_135
timestamp 1676037725
transform 1 0 13524 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1676037725
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1676037725
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1676037725
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_177
timestamp 1676037725
transform 1 0 17388 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_185
timestamp 1676037725
transform 1 0 18124 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_190
timestamp 1676037725
transform 1 0 18584 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1676037725
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1676037725
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1676037725
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1676037725
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1676037725
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1676037725
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1676037725
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1676037725
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1676037725
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1676037725
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1676037725
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1676037725
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1676037725
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1676037725
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1676037725
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1676037725
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1676037725
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1676037725
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1676037725
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_401
timestamp 1676037725
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1676037725
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1676037725
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1676037725
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1676037725
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_445
timestamp 1676037725
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_457
timestamp 1676037725
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1676037725
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1676037725
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1676037725
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1676037725
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1676037725
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_513
timestamp 1676037725
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1676037725
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1676037725
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_533
timestamp 1676037725
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_545
timestamp 1676037725
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_557
timestamp 1676037725
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_569
timestamp 1676037725
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1676037725
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1676037725
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_589
timestamp 1676037725
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_601
timestamp 1676037725
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_613
timestamp 1676037725
transform 1 0 57500 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_623
timestamp 1676037725
transform 1 0 58420 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1676037725
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1676037725
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1676037725
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1676037725
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1676037725
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1676037725
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1676037725
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1676037725
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1676037725
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1676037725
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_119
timestamp 1676037725
transform 1 0 12052 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_129
timestamp 1676037725
transform 1 0 12972 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_141
timestamp 1676037725
transform 1 0 14076 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_153
timestamp 1676037725
transform 1 0 15180 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_165
timestamp 1676037725
transform 1 0 16284 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1676037725
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1676037725
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1676037725
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1676037725
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1676037725
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1676037725
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1676037725
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1676037725
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1676037725
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1676037725
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1676037725
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1676037725
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1676037725
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1676037725
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1676037725
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1676037725
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1676037725
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1676037725
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1676037725
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1676037725
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1676037725
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1676037725
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1676037725
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_405
timestamp 1676037725
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_417
timestamp 1676037725
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_429
timestamp 1676037725
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1676037725
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1676037725
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1676037725
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1676037725
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1676037725
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1676037725
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1676037725
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1676037725
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_505
timestamp 1676037725
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_517
timestamp 1676037725
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_529
timestamp 1676037725
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_541
timestamp 1676037725
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1676037725
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1676037725
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_561
timestamp 1676037725
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_573
timestamp 1676037725
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_585
timestamp 1676037725
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_597
timestamp 1676037725
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1676037725
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1676037725
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_617
timestamp 1676037725
transform 1 0 57868 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_11
timestamp 1676037725
transform 1 0 2116 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_24
timestamp 1676037725
transform 1 0 3312 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1676037725
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1676037725
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1676037725
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1676037725
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1676037725
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1676037725
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1676037725
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1676037725
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1676037725
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1676037725
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1676037725
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1676037725
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1676037725
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1676037725
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1676037725
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1676037725
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1676037725
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1676037725
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1676037725
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1676037725
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1676037725
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1676037725
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1676037725
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1676037725
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1676037725
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1676037725
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1676037725
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1676037725
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1676037725
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1676037725
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1676037725
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1676037725
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1676037725
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1676037725
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1676037725
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1676037725
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1676037725
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1676037725
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_433
timestamp 1676037725
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_445
timestamp 1676037725
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_457
timestamp 1676037725
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1676037725
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1676037725
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1676037725
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1676037725
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1676037725
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_513
timestamp 1676037725
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1676037725
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1676037725
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_533
timestamp 1676037725
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_545
timestamp 1676037725
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_557
timestamp 1676037725
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_569
timestamp 1676037725
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1676037725
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1676037725
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_589
timestamp 1676037725
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_601
timestamp 1676037725
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_613
timestamp 1676037725
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1676037725
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_11
timestamp 1676037725
transform 1 0 2116 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_23
timestamp 1676037725
transform 1 0 3220 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_35
timestamp 1676037725
transform 1 0 4324 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_47
timestamp 1676037725
transform 1 0 5428 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1676037725
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1676037725
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1676037725
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1676037725
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1676037725
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1676037725
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1676037725
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1676037725
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1676037725
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1676037725
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1676037725
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1676037725
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1676037725
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1676037725
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1676037725
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1676037725
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1676037725
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1676037725
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1676037725
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1676037725
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1676037725
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1676037725
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1676037725
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1676037725
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1676037725
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1676037725
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1676037725
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1676037725
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1676037725
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1676037725
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1676037725
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1676037725
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1676037725
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1676037725
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1676037725
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1676037725
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1676037725
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1676037725
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_405
timestamp 1676037725
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_417
timestamp 1676037725
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_429
timestamp 1676037725
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1676037725
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1676037725
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1676037725
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1676037725
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1676037725
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1676037725
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1676037725
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1676037725
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_505
timestamp 1676037725
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_517
timestamp 1676037725
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_529
timestamp 1676037725
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1676037725
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1676037725
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1676037725
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_561
timestamp 1676037725
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_573
timestamp 1676037725
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_585
timestamp 1676037725
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_597
timestamp 1676037725
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1676037725
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1676037725
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_617
timestamp 1676037725
transform 1 0 57868 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_623
timestamp 1676037725
transform 1 0 58420 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1676037725
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_11
timestamp 1676037725
transform 1 0 2116 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_20
timestamp 1676037725
transform 1 0 2944 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1676037725
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1676037725
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1676037725
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1676037725
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1676037725
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1676037725
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1676037725
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1676037725
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1676037725
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1676037725
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1676037725
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1676037725
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1676037725
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1676037725
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1676037725
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1676037725
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1676037725
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1676037725
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1676037725
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1676037725
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1676037725
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1676037725
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1676037725
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1676037725
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1676037725
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1676037725
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1676037725
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1676037725
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1676037725
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1676037725
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1676037725
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1676037725
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1676037725
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1676037725
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1676037725
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1676037725
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1676037725
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1676037725
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1676037725
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_401
timestamp 1676037725
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1676037725
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1676037725
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1676037725
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1676037725
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1676037725
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1676037725
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1676037725
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1676037725
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1676037725
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1676037725
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1676037725
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_513
timestamp 1676037725
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1676037725
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1676037725
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_533
timestamp 1676037725
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_545
timestamp 1676037725
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_557
timestamp 1676037725
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_569
timestamp 1676037725
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1676037725
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1676037725
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_589
timestamp 1676037725
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_601
timestamp 1676037725
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_613
timestamp 1676037725
transform 1 0 57500 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_623
timestamp 1676037725
transform 1 0 58420 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_3
timestamp 1676037725
transform 1 0 1380 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_11
timestamp 1676037725
transform 1 0 2116 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_23
timestamp 1676037725
transform 1 0 3220 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_35
timestamp 1676037725
transform 1 0 4324 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_47
timestamp 1676037725
transform 1 0 5428 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1676037725
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1676037725
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1676037725
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1676037725
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_93
timestamp 1676037725
transform 1 0 9660 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_101
timestamp 1676037725
transform 1 0 10396 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_109
timestamp 1676037725
transform 1 0 11132 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1676037725
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1676037725
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1676037725
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1676037725
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1676037725
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1676037725
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1676037725
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1676037725
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1676037725
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1676037725
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1676037725
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1676037725
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1676037725
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1676037725
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1676037725
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1676037725
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1676037725
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1676037725
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1676037725
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1676037725
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1676037725
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1676037725
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1676037725
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1676037725
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1676037725
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1676037725
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1676037725
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1676037725
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1676037725
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1676037725
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1676037725
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 1676037725
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_417
timestamp 1676037725
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1676037725
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1676037725
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1676037725
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1676037725
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1676037725
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1676037725
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1676037725
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1676037725
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1676037725
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1676037725
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1676037725
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1676037725
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1676037725
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1676037725
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1676037725
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_561
timestamp 1676037725
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_573
timestamp 1676037725
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_585
timestamp 1676037725
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_597
timestamp 1676037725
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1676037725
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1676037725
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_617
timestamp 1676037725
transform 1 0 57868 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_623
timestamp 1676037725
transform 1 0 58420 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1676037725
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1676037725
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1676037725
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1676037725
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1676037725
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1676037725
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1676037725
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1676037725
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1676037725
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1676037725
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1676037725
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1676037725
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1676037725
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1676037725
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1676037725
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1676037725
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1676037725
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1676037725
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1676037725
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1676037725
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1676037725
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1676037725
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1676037725
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1676037725
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1676037725
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1676037725
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1676037725
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1676037725
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1676037725
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1676037725
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1676037725
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1676037725
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1676037725
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1676037725
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1676037725
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1676037725
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1676037725
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1676037725
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1676037725
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1676037725
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1676037725
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1676037725
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_401
timestamp 1676037725
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1676037725
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1676037725
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1676037725
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1676037725
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1676037725
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1676037725
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1676037725
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1676037725
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1676037725
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1676037725
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1676037725
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_513
timestamp 1676037725
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1676037725
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1676037725
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_533
timestamp 1676037725
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_545
timestamp 1676037725
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_557
timestamp 1676037725
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_569
timestamp 1676037725
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1676037725
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1676037725
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_589
timestamp 1676037725
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_601
timestamp 1676037725
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_613
timestamp 1676037725
transform 1 0 57500 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_623
timestamp 1676037725
transform 1 0 58420 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1676037725
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_11
timestamp 1676037725
transform 1 0 2116 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_20
timestamp 1676037725
transform 1 0 2944 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_32
timestamp 1676037725
transform 1 0 4048 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_44
timestamp 1676037725
transform 1 0 5152 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1676037725
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1676037725
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1676037725
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1676037725
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1676037725
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1676037725
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1676037725
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1676037725
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1676037725
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1676037725
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1676037725
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1676037725
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1676037725
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1676037725
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1676037725
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1676037725
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1676037725
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1676037725
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_225
timestamp 1676037725
transform 1 0 21804 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_233
timestamp 1676037725
transform 1 0 22540 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_244
timestamp 1676037725
transform 1 0 23552 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_256
timestamp 1676037725
transform 1 0 24656 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_268
timestamp 1676037725
transform 1 0 25760 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1676037725
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1676037725
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1676037725
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1676037725
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1676037725
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1676037725
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1676037725
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1676037725
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1676037725
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1676037725
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1676037725
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1676037725
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1676037725
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1676037725
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1676037725
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1676037725
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1676037725
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1676037725
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1676037725
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1676037725
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1676037725
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1676037725
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1676037725
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1676037725
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1676037725
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_517
timestamp 1676037725
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_529
timestamp 1676037725
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_541
timestamp 1676037725
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1676037725
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1676037725
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_561
timestamp 1676037725
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_573
timestamp 1676037725
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_585
timestamp 1676037725
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_597
timestamp 1676037725
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1676037725
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1676037725
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_617
timestamp 1676037725
transform 1 0 57868 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1676037725
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_11
timestamp 1676037725
transform 1 0 2116 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_23
timestamp 1676037725
transform 1 0 3220 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1676037725
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1676037725
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1676037725
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1676037725
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1676037725
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1676037725
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1676037725
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1676037725
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1676037725
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1676037725
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1676037725
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1676037725
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1676037725
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1676037725
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1676037725
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1676037725
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1676037725
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1676037725
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1676037725
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1676037725
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1676037725
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1676037725
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_233
timestamp 1676037725
transform 1 0 22540 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_247
timestamp 1676037725
transform 1 0 23828 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1676037725
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1676037725
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1676037725
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1676037725
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1676037725
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1676037725
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1676037725
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1676037725
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1676037725
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1676037725
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1676037725
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1676037725
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1676037725
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1676037725
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1676037725
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1676037725
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_401
timestamp 1676037725
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1676037725
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1676037725
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1676037725
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1676037725
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1676037725
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1676037725
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1676037725
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1676037725
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1676037725
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1676037725
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1676037725
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_513
timestamp 1676037725
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1676037725
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1676037725
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_533
timestamp 1676037725
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_545
timestamp 1676037725
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_557
timestamp 1676037725
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_569
timestamp 1676037725
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1676037725
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1676037725
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_589
timestamp 1676037725
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_601
timestamp 1676037725
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_613
timestamp 1676037725
transform 1 0 57500 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_623
timestamp 1676037725
transform 1 0 58420 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1676037725
transform 1 0 1380 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_11
timestamp 1676037725
transform 1 0 2116 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_23
timestamp 1676037725
transform 1 0 3220 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_35
timestamp 1676037725
transform 1 0 4324 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_47
timestamp 1676037725
transform 1 0 5428 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1676037725
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1676037725
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1676037725
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1676037725
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1676037725
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1676037725
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1676037725
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1676037725
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1676037725
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1676037725
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1676037725
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1676037725
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1676037725
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1676037725
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1676037725
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1676037725
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1676037725
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1676037725
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1676037725
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1676037725
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_237
timestamp 1676037725
transform 1 0 22908 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_246
timestamp 1676037725
transform 1 0 23736 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_258
timestamp 1676037725
transform 1 0 24840 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_270
timestamp 1676037725
transform 1 0 25944 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_278
timestamp 1676037725
transform 1 0 26680 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1676037725
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1676037725
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1676037725
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1676037725
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1676037725
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1676037725
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1676037725
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1676037725
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1676037725
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1676037725
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1676037725
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1676037725
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1676037725
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1676037725
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1676037725
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1676037725
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1676037725
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1676037725
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1676037725
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1676037725
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1676037725
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1676037725
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1676037725
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1676037725
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1676037725
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_517
timestamp 1676037725
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_529
timestamp 1676037725
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_541
timestamp 1676037725
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1676037725
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1676037725
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_561
timestamp 1676037725
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_573
timestamp 1676037725
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_585
timestamp 1676037725
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_597
timestamp 1676037725
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 1676037725
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1676037725
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_617
timestamp 1676037725
transform 1 0 57868 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_3
timestamp 1676037725
transform 1 0 1380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_11
timestamp 1676037725
transform 1 0 2116 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_20
timestamp 1676037725
transform 1 0 2944 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1676037725
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1676037725
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1676037725
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1676037725
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1676037725
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1676037725
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1676037725
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1676037725
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1676037725
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1676037725
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1676037725
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1676037725
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1676037725
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1676037725
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1676037725
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1676037725
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1676037725
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1676037725
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1676037725
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1676037725
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1676037725
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1676037725
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1676037725
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1676037725
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1676037725
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1676037725
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1676037725
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1676037725
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1676037725
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1676037725
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1676037725
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1676037725
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1676037725
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1676037725
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1676037725
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1676037725
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1676037725
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1676037725
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1676037725
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_401
timestamp 1676037725
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1676037725
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1676037725
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1676037725
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1676037725
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1676037725
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1676037725
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1676037725
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1676037725
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1676037725
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1676037725
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1676037725
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_513
timestamp 1676037725
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1676037725
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1676037725
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_533
timestamp 1676037725
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_545
timestamp 1676037725
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_557
timestamp 1676037725
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_569
timestamp 1676037725
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1676037725
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1676037725
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_589
timestamp 1676037725
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_601
timestamp 1676037725
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_613
timestamp 1676037725
transform 1 0 57500 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_623
timestamp 1676037725
transform 1 0 58420 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1676037725
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1676037725
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1676037725
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1676037725
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1676037725
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1676037725
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1676037725
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1676037725
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_81
timestamp 1676037725
transform 1 0 8556 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_94
timestamp 1676037725
transform 1 0 9752 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_106
timestamp 1676037725
transform 1 0 10856 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1676037725
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1676037725
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1676037725
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1676037725
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1676037725
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1676037725
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1676037725
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1676037725
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1676037725
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1676037725
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1676037725
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1676037725
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1676037725
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1676037725
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1676037725
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1676037725
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1676037725
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1676037725
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1676037725
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1676037725
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1676037725
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1676037725
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1676037725
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1676037725
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1676037725
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1676037725
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1676037725
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1676037725
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1676037725
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1676037725
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1676037725
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1676037725
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1676037725
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1676037725
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1676037725
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1676037725
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1676037725
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1676037725
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1676037725
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1676037725
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1676037725
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1676037725
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1676037725
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_517
timestamp 1676037725
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_529
timestamp 1676037725
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_541
timestamp 1676037725
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1676037725
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1676037725
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_561
timestamp 1676037725
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_573
timestamp 1676037725
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_585
timestamp 1676037725
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_597
timestamp 1676037725
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 1676037725
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1676037725
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_617
timestamp 1676037725
transform 1 0 57868 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1676037725
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_11
timestamp 1676037725
transform 1 0 2116 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_23
timestamp 1676037725
transform 1 0 3220 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1676037725
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1676037725
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1676037725
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1676037725
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1676037725
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1676037725
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1676037725
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1676037725
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1676037725
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1676037725
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1676037725
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1676037725
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1676037725
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1676037725
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1676037725
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1676037725
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1676037725
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1676037725
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1676037725
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1676037725
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1676037725
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_221
timestamp 1676037725
transform 1 0 21436 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_229
timestamp 1676037725
transform 1 0 22172 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_240
timestamp 1676037725
transform 1 0 23184 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1676037725
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1676037725
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1676037725
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1676037725
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1676037725
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1676037725
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1676037725
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1676037725
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1676037725
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1676037725
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1676037725
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1676037725
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1676037725
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1676037725
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1676037725
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1676037725
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1676037725
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1676037725
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1676037725
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1676037725
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1676037725
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1676037725
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1676037725
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1676037725
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1676037725
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1676037725
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1676037725
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_513
timestamp 1676037725
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1676037725
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1676037725
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_533
timestamp 1676037725
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_545
timestamp 1676037725
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_557
timestamp 1676037725
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_569
timestamp 1676037725
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1676037725
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1676037725
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_589
timestamp 1676037725
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_601
timestamp 1676037725
transform 1 0 56396 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_613
timestamp 1676037725
transform 1 0 57500 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_623
timestamp 1676037725
transform 1 0 58420 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_3
timestamp 1676037725
transform 1 0 1380 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_11
timestamp 1676037725
transform 1 0 2116 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_23
timestamp 1676037725
transform 1 0 3220 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_35
timestamp 1676037725
transform 1 0 4324 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_47
timestamp 1676037725
transform 1 0 5428 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1676037725
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1676037725
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1676037725
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1676037725
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1676037725
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1676037725
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1676037725
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1676037725
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1676037725
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1676037725
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1676037725
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1676037725
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1676037725
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1676037725
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_181
timestamp 1676037725
transform 1 0 17756 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_189
timestamp 1676037725
transform 1 0 18492 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_199
timestamp 1676037725
transform 1 0 19412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_211
timestamp 1676037725
transform 1 0 20516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1676037725
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_225
timestamp 1676037725
transform 1 0 21804 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_229
timestamp 1676037725
transform 1 0 22172 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_239
timestamp 1676037725
transform 1 0 23092 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_251
timestamp 1676037725
transform 1 0 24196 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_263
timestamp 1676037725
transform 1 0 25300 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_275
timestamp 1676037725
transform 1 0 26404 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1676037725
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1676037725
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1676037725
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1676037725
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1676037725
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1676037725
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1676037725
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1676037725
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1676037725
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1676037725
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1676037725
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1676037725
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1676037725
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1676037725
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1676037725
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_417
timestamp 1676037725
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_429
timestamp 1676037725
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1676037725
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1676037725
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1676037725
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1676037725
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1676037725
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1676037725
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1676037725
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1676037725
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1676037725
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_517
timestamp 1676037725
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_529
timestamp 1676037725
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_541
timestamp 1676037725
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1676037725
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1676037725
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_561
timestamp 1676037725
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_573
timestamp 1676037725
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_585
timestamp 1676037725
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_597
timestamp 1676037725
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1676037725
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1676037725
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_617
timestamp 1676037725
transform 1 0 57868 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1676037725
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_9
timestamp 1676037725
transform 1 0 1932 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_21
timestamp 1676037725
transform 1 0 3036 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1676037725
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1676037725
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1676037725
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1676037725
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1676037725
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1676037725
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1676037725
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1676037725
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1676037725
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1676037725
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1676037725
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1676037725
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1676037725
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1676037725
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1676037725
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1676037725
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1676037725
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1676037725
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1676037725
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_197
timestamp 1676037725
transform 1 0 19228 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_208
timestamp 1676037725
transform 1 0 20240 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_220
timestamp 1676037725
transform 1 0 21344 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_234
timestamp 1676037725
transform 1 0 22632 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1676037725
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1676037725
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1676037725
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1676037725
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1676037725
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1676037725
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1676037725
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1676037725
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1676037725
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1676037725
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1676037725
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1676037725
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1676037725
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1676037725
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1676037725
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1676037725
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1676037725
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_401
timestamp 1676037725
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1676037725
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1676037725
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1676037725
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1676037725
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1676037725
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1676037725
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1676037725
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1676037725
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1676037725
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1676037725
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1676037725
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_513
timestamp 1676037725
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1676037725
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1676037725
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_533
timestamp 1676037725
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_545
timestamp 1676037725
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_557
timestamp 1676037725
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_569
timestamp 1676037725
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1676037725
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1676037725
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_589
timestamp 1676037725
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_601
timestamp 1676037725
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_613
timestamp 1676037725
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1676037725
transform 1 0 1380 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_9
timestamp 1676037725
transform 1 0 1932 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_21
timestamp 1676037725
transform 1 0 3036 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_33
timestamp 1676037725
transform 1 0 4140 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_45
timestamp 1676037725
transform 1 0 5244 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_53
timestamp 1676037725
transform 1 0 5980 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1676037725
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1676037725
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1676037725
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1676037725
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1676037725
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1676037725
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1676037725
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1676037725
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1676037725
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1676037725
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1676037725
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1676037725
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1676037725
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1676037725
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1676037725
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1676037725
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1676037725
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1676037725
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1676037725
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1676037725
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_249
timestamp 1676037725
transform 1 0 24012 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_258
timestamp 1676037725
transform 1 0 24840 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_270
timestamp 1676037725
transform 1 0 25944 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_278
timestamp 1676037725
transform 1 0 26680 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1676037725
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1676037725
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1676037725
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1676037725
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1676037725
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1676037725
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1676037725
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1676037725
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1676037725
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1676037725
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1676037725
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1676037725
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1676037725
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1676037725
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1676037725
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1676037725
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1676037725
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1676037725
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1676037725
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1676037725
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1676037725
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1676037725
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1676037725
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1676037725
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1676037725
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_517
timestamp 1676037725
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_529
timestamp 1676037725
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_541
timestamp 1676037725
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1676037725
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1676037725
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_561
timestamp 1676037725
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_573
timestamp 1676037725
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_585
timestamp 1676037725
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_597
timestamp 1676037725
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1676037725
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1676037725
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_617
timestamp 1676037725
transform 1 0 57868 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_623
timestamp 1676037725
transform 1 0 58420 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1676037725
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1676037725
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1676037725
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1676037725
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1676037725
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1676037725
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1676037725
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1676037725
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1676037725
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1676037725
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1676037725
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1676037725
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1676037725
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1676037725
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1676037725
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1676037725
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1676037725
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1676037725
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1676037725
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1676037725
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1676037725
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1676037725
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1676037725
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_221
timestamp 1676037725
transform 1 0 21436 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_229
timestamp 1676037725
transform 1 0 22172 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_233
timestamp 1676037725
transform 1 0 22540 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_242
timestamp 1676037725
transform 1 0 23368 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_250
timestamp 1676037725
transform 1 0 24104 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1676037725
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1676037725
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1676037725
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1676037725
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1676037725
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1676037725
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1676037725
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1676037725
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1676037725
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1676037725
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1676037725
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1676037725
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1676037725
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1676037725
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1676037725
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_401
timestamp 1676037725
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1676037725
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1676037725
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1676037725
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1676037725
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1676037725
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1676037725
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1676037725
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1676037725
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1676037725
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1676037725
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1676037725
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_513
timestamp 1676037725
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1676037725
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1676037725
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_533
timestamp 1676037725
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_545
timestamp 1676037725
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_557
timestamp 1676037725
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_569
timestamp 1676037725
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1676037725
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1676037725
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_589
timestamp 1676037725
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_601
timestamp 1676037725
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_613
timestamp 1676037725
transform 1 0 57500 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_623
timestamp 1676037725
transform 1 0 58420 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1676037725
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_9
timestamp 1676037725
transform 1 0 1932 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_21
timestamp 1676037725
transform 1 0 3036 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_33
timestamp 1676037725
transform 1 0 4140 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_45
timestamp 1676037725
transform 1 0 5244 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_53
timestamp 1676037725
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1676037725
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1676037725
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1676037725
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1676037725
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1676037725
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1676037725
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1676037725
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1676037725
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1676037725
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1676037725
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1676037725
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1676037725
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1676037725
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1676037725
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1676037725
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1676037725
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1676037725
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1676037725
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1676037725
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1676037725
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1676037725
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1676037725
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1676037725
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1676037725
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1676037725
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1676037725
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1676037725
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1676037725
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1676037725
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1676037725
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1676037725
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1676037725
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1676037725
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1676037725
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1676037725
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1676037725
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1676037725
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1676037725
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_417
timestamp 1676037725
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1676037725
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1676037725
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1676037725
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1676037725
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1676037725
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1676037725
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1676037725
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1676037725
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1676037725
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1676037725
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_517
timestamp 1676037725
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_529
timestamp 1676037725
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1676037725
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1676037725
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1676037725
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_561
timestamp 1676037725
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_573
timestamp 1676037725
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_585
timestamp 1676037725
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_597
timestamp 1676037725
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1676037725
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1676037725
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_617
timestamp 1676037725
transform 1 0 57868 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1676037725
transform 1 0 1380 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_9
timestamp 1676037725
transform 1 0 1932 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_21
timestamp 1676037725
transform 1 0 3036 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1676037725
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1676037725
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1676037725
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1676037725
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1676037725
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1676037725
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1676037725
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1676037725
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1676037725
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1676037725
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1676037725
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1676037725
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1676037725
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1676037725
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1676037725
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1676037725
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1676037725
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1676037725
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1676037725
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1676037725
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1676037725
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_221
timestamp 1676037725
transform 1 0 21436 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_234
timestamp 1676037725
transform 1 0 22632 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_246
timestamp 1676037725
transform 1 0 23736 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_253
timestamp 1676037725
transform 1 0 24380 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_266
timestamp 1676037725
transform 1 0 25576 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_278
timestamp 1676037725
transform 1 0 26680 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_290
timestamp 1676037725
transform 1 0 27784 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_302
timestamp 1676037725
transform 1 0 28888 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1676037725
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1676037725
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1676037725
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1676037725
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1676037725
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1676037725
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1676037725
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1676037725
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1676037725
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1676037725
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1676037725
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1676037725
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1676037725
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1676037725
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1676037725
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1676037725
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1676037725
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1676037725
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1676037725
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1676037725
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1676037725
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_513
timestamp 1676037725
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1676037725
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1676037725
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_533
timestamp 1676037725
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_545
timestamp 1676037725
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_557
timestamp 1676037725
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_569
timestamp 1676037725
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1676037725
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1676037725
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_589
timestamp 1676037725
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_601
timestamp 1676037725
transform 1 0 56396 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_613
timestamp 1676037725
transform 1 0 57500 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_623
timestamp 1676037725
transform 1 0 58420 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_3
timestamp 1676037725
transform 1 0 1380 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_9
timestamp 1676037725
transform 1 0 1932 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_21
timestamp 1676037725
transform 1 0 3036 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_33
timestamp 1676037725
transform 1 0 4140 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_45
timestamp 1676037725
transform 1 0 5244 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_53
timestamp 1676037725
transform 1 0 5980 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1676037725
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1676037725
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1676037725
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1676037725
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1676037725
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1676037725
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1676037725
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1676037725
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1676037725
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1676037725
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1676037725
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1676037725
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1676037725
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1676037725
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1676037725
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_205
timestamp 1676037725
transform 1 0 19964 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_57_213
timestamp 1676037725
transform 1 0 20700 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_222
timestamp 1676037725
transform 1 0 21528 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_225
timestamp 1676037725
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_235
timestamp 1676037725
transform 1 0 22724 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_247
timestamp 1676037725
transform 1 0 23828 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_259
timestamp 1676037725
transform 1 0 24932 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_271
timestamp 1676037725
transform 1 0 26036 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1676037725
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1676037725
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1676037725
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1676037725
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1676037725
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1676037725
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1676037725
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1676037725
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1676037725
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1676037725
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_373
timestamp 1676037725
transform 1 0 35420 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1676037725
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1676037725
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1676037725
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1676037725
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1676037725
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1676037725
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1676037725
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1676037725
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1676037725
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1676037725
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1676037725
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1676037725
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1676037725
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1676037725
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1676037725
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_517
timestamp 1676037725
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_529
timestamp 1676037725
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_541
timestamp 1676037725
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1676037725
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1676037725
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_561
timestamp 1676037725
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_573
timestamp 1676037725
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_585
timestamp 1676037725
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_597
timestamp 1676037725
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1676037725
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1676037725
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_617
timestamp 1676037725
transform 1 0 57868 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_3
timestamp 1676037725
transform 1 0 1380 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_9
timestamp 1676037725
transform 1 0 1932 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_21
timestamp 1676037725
transform 1 0 3036 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1676037725
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1676037725
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1676037725
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1676037725
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1676037725
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1676037725
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1676037725
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1676037725
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1676037725
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1676037725
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1676037725
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1676037725
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1676037725
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1676037725
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1676037725
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1676037725
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1676037725
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1676037725
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1676037725
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1676037725
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_209
timestamp 1676037725
transform 1 0 20332 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_217
timestamp 1676037725
transform 1 0 21068 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_229
timestamp 1676037725
transform 1 0 22172 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_242
timestamp 1676037725
transform 1 0 23368 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_250
timestamp 1676037725
transform 1 0 24104 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1676037725
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_263
timestamp 1676037725
transform 1 0 25300 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_275
timestamp 1676037725
transform 1 0 26404 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_287
timestamp 1676037725
transform 1 0 27508 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_299
timestamp 1676037725
transform 1 0 28612 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1676037725
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1676037725
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1676037725
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1676037725
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1676037725
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1676037725
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1676037725
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1676037725
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1676037725
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1676037725
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_401
timestamp 1676037725
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1676037725
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1676037725
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1676037725
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1676037725
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1676037725
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1676037725
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1676037725
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1676037725
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1676037725
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1676037725
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1676037725
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_513
timestamp 1676037725
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1676037725
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1676037725
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_533
timestamp 1676037725
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_545
timestamp 1676037725
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_557
timestamp 1676037725
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_569
timestamp 1676037725
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1676037725
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1676037725
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_589
timestamp 1676037725
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_601
timestamp 1676037725
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_613
timestamp 1676037725
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1676037725
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1676037725
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1676037725
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1676037725
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1676037725
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1676037725
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1676037725
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1676037725
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1676037725
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1676037725
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1676037725
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1676037725
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1676037725
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1676037725
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1676037725
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1676037725
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1676037725
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1676037725
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1676037725
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1676037725
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1676037725
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1676037725
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1676037725
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1676037725
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1676037725
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1676037725
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1676037725
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1676037725
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1676037725
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1676037725
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1676037725
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1676037725
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1676037725
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1676037725
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1676037725
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1676037725
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1676037725
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1676037725
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1676037725
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1676037725
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1676037725
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1676037725
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1676037725
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1676037725
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1676037725
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1676037725
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1676037725
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1676037725
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1676037725
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1676037725
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1676037725
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1676037725
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1676037725
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1676037725
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1676037725
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_517
timestamp 1676037725
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_529
timestamp 1676037725
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_541
timestamp 1676037725
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1676037725
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1676037725
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_561
timestamp 1676037725
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_573
timestamp 1676037725
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_585
timestamp 1676037725
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_597
timestamp 1676037725
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1676037725
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1676037725
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_617
timestamp 1676037725
transform 1 0 57868 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_623
timestamp 1676037725
transform 1 0 58420 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_3
timestamp 1676037725
transform 1 0 1380 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_9
timestamp 1676037725
transform 1 0 1932 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_21
timestamp 1676037725
transform 1 0 3036 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1676037725
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1676037725
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1676037725
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1676037725
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1676037725
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1676037725
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1676037725
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1676037725
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1676037725
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1676037725
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1676037725
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1676037725
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1676037725
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1676037725
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1676037725
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1676037725
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1676037725
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1676037725
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1676037725
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1676037725
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1676037725
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1676037725
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_240
timestamp 1676037725
transform 1 0 23184 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1676037725
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1676037725
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1676037725
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1676037725
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1676037725
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1676037725
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1676037725
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1676037725
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1676037725
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1676037725
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1676037725
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1676037725
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1676037725
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1676037725
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1676037725
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_401
timestamp 1676037725
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1676037725
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1676037725
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_421
timestamp 1676037725
transform 1 0 39836 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_430
timestamp 1676037725
transform 1 0 40664 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_442
timestamp 1676037725
transform 1 0 41768 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_454
timestamp 1676037725
transform 1 0 42872 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_466
timestamp 1676037725
transform 1 0 43976 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_474
timestamp 1676037725
transform 1 0 44712 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1676037725
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1676037725
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1676037725
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_513
timestamp 1676037725
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1676037725
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1676037725
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_533
timestamp 1676037725
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_545
timestamp 1676037725
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_557
timestamp 1676037725
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_569
timestamp 1676037725
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1676037725
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1676037725
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_589
timestamp 1676037725
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_601
timestamp 1676037725
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_613
timestamp 1676037725
transform 1 0 57500 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_623
timestamp 1676037725
transform 1 0 58420 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_3
timestamp 1676037725
transform 1 0 1380 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_9
timestamp 1676037725
transform 1 0 1932 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_21
timestamp 1676037725
transform 1 0 3036 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_33
timestamp 1676037725
transform 1 0 4140 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_45
timestamp 1676037725
transform 1 0 5244 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_53
timestamp 1676037725
transform 1 0 5980 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1676037725
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1676037725
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1676037725
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1676037725
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1676037725
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1676037725
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1676037725
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1676037725
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1676037725
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1676037725
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1676037725
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1676037725
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1676037725
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1676037725
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_193
timestamp 1676037725
transform 1 0 18860 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_202
timestamp 1676037725
transform 1 0 19688 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_211
timestamp 1676037725
transform 1 0 20516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1676037725
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_225
timestamp 1676037725
transform 1 0 21804 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_233
timestamp 1676037725
transform 1 0 22540 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_246
timestamp 1676037725
transform 1 0 23736 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_258
timestamp 1676037725
transform 1 0 24840 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_270
timestamp 1676037725
transform 1 0 25944 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_278
timestamp 1676037725
transform 1 0 26680 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1676037725
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1676037725
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1676037725
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1676037725
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1676037725
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1676037725
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1676037725
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1676037725
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1676037725
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1676037725
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1676037725
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1676037725
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1676037725
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1676037725
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_417
timestamp 1676037725
transform 1 0 39468 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_61_432
timestamp 1676037725
transform 1 0 40848 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_444
timestamp 1676037725
transform 1 0 41952 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1676037725
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1676037725
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1676037725
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1676037725
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1676037725
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1676037725
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1676037725
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_517
timestamp 1676037725
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_529
timestamp 1676037725
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_541
timestamp 1676037725
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1676037725
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1676037725
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_561
timestamp 1676037725
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_573
timestamp 1676037725
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_585
timestamp 1676037725
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_597
timestamp 1676037725
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1676037725
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1676037725
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_617
timestamp 1676037725
transform 1 0 57868 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1676037725
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_9
timestamp 1676037725
transform 1 0 1932 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_23
timestamp 1676037725
transform 1 0 3220 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1676037725
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1676037725
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1676037725
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1676037725
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1676037725
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1676037725
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1676037725
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1676037725
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1676037725
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1676037725
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1676037725
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1676037725
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1676037725
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1676037725
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1676037725
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1676037725
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1676037725
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1676037725
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1676037725
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_197
timestamp 1676037725
transform 1 0 19228 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_205
timestamp 1676037725
transform 1 0 19964 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_216
timestamp 1676037725
transform 1 0 20976 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_228
timestamp 1676037725
transform 1 0 22080 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_236
timestamp 1676037725
transform 1 0 22816 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_240
timestamp 1676037725
transform 1 0 23184 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_248
timestamp 1676037725
transform 1 0 23920 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_253
timestamp 1676037725
transform 1 0 24380 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_262
timestamp 1676037725
transform 1 0 25208 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_274
timestamp 1676037725
transform 1 0 26312 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_286
timestamp 1676037725
transform 1 0 27416 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_298
timestamp 1676037725
transform 1 0 28520 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_306
timestamp 1676037725
transform 1 0 29256 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1676037725
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1676037725
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1676037725
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1676037725
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1676037725
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1676037725
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1676037725
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1676037725
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1676037725
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_401
timestamp 1676037725
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1676037725
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1676037725
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1676037725
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1676037725
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1676037725
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1676037725
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1676037725
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1676037725
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1676037725
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1676037725
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1676037725
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_513
timestamp 1676037725
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1676037725
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1676037725
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_533
timestamp 1676037725
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_545
timestamp 1676037725
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_557
timestamp 1676037725
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_569
timestamp 1676037725
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1676037725
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1676037725
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_589
timestamp 1676037725
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_601
timestamp 1676037725
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_613
timestamp 1676037725
transform 1 0 57500 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_623
timestamp 1676037725
transform 1 0 58420 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1676037725
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_9
timestamp 1676037725
transform 1 0 1932 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_21
timestamp 1676037725
transform 1 0 3036 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_33
timestamp 1676037725
transform 1 0 4140 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_45
timestamp 1676037725
transform 1 0 5244 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_53
timestamp 1676037725
transform 1 0 5980 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1676037725
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1676037725
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1676037725
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1676037725
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1676037725
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1676037725
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1676037725
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1676037725
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1676037725
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1676037725
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1676037725
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1676037725
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1676037725
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_181
timestamp 1676037725
transform 1 0 17756 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_187
timestamp 1676037725
transform 1 0 18308 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_195
timestamp 1676037725
transform 1 0 19044 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_219
timestamp 1676037725
transform 1 0 21252 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1676037725
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1676037725
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_237
timestamp 1676037725
transform 1 0 22908 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_241
timestamp 1676037725
transform 1 0 23276 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_244
timestamp 1676037725
transform 1 0 23552 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_252
timestamp 1676037725
transform 1 0 24288 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_264
timestamp 1676037725
transform 1 0 25392 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_276
timestamp 1676037725
transform 1 0 26496 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1676037725
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1676037725
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1676037725
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1676037725
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1676037725
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1676037725
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1676037725
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1676037725
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1676037725
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1676037725
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1676037725
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1676037725
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1676037725
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1676037725
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1676037725
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1676037725
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1676037725
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1676037725
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1676037725
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1676037725
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1676037725
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1676037725
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1676037725
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1676037725
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1676037725
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_517
timestamp 1676037725
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_529
timestamp 1676037725
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_541
timestamp 1676037725
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1676037725
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1676037725
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_561
timestamp 1676037725
transform 1 0 52716 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_569
timestamp 1676037725
transform 1 0 53452 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_579
timestamp 1676037725
transform 1 0 54372 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_591
timestamp 1676037725
transform 1 0 55476 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_603
timestamp 1676037725
transform 1 0 56580 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1676037725
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_617
timestamp 1676037725
transform 1 0 57868 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1676037725
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_9
timestamp 1676037725
transform 1 0 1932 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_21
timestamp 1676037725
transform 1 0 3036 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1676037725
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1676037725
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_41
timestamp 1676037725
transform 1 0 4876 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_64
timestamp 1676037725
transform 1 0 6992 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_76
timestamp 1676037725
transform 1 0 8096 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1676037725
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1676037725
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1676037725
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1676037725
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1676037725
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1676037725
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1676037725
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1676037725
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1676037725
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1676037725
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1676037725
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1676037725
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_197
timestamp 1676037725
transform 1 0 19228 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_209
timestamp 1676037725
transform 1 0 20332 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_225
timestamp 1676037725
transform 1 0 21804 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_237
timestamp 1676037725
transform 1 0 22908 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_249
timestamp 1676037725
transform 1 0 24012 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1676037725
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1676037725
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_277
timestamp 1676037725
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_289
timestamp 1676037725
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1676037725
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1676037725
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1676037725
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1676037725
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_333
timestamp 1676037725
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_345
timestamp 1676037725
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1676037725
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1676037725
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1676037725
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1676037725
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_389
timestamp 1676037725
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_401
timestamp 1676037725
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1676037725
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1676037725
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1676037725
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1676037725
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1676037725
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1676037725
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1676037725
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1676037725
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1676037725
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1676037725
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1676037725
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_513
timestamp 1676037725
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1676037725
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1676037725
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_533
timestamp 1676037725
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_545
timestamp 1676037725
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_557
timestamp 1676037725
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_569
timestamp 1676037725
transform 1 0 53452 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_581
timestamp 1676037725
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 1676037725
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_589
timestamp 1676037725
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_601
timestamp 1676037725
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_613
timestamp 1676037725
transform 1 0 57500 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_623
timestamp 1676037725
transform 1 0 58420 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_65_3
timestamp 1676037725
transform 1 0 1380 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_9
timestamp 1676037725
transform 1 0 1932 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_17
timestamp 1676037725
transform 1 0 2668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_29
timestamp 1676037725
transform 1 0 3772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_41
timestamp 1676037725
transform 1 0 4876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_53
timestamp 1676037725
transform 1 0 5980 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1676037725
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1676037725
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1676037725
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1676037725
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1676037725
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1676037725
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1676037725
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1676037725
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1676037725
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1676037725
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1676037725
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1676037725
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1676037725
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1676037725
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_193
timestamp 1676037725
transform 1 0 18860 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_197
timestamp 1676037725
transform 1 0 19228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_206
timestamp 1676037725
transform 1 0 20056 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_210
timestamp 1676037725
transform 1 0 20424 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_65_218
timestamp 1676037725
transform 1 0 21160 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_65_225
timestamp 1676037725
transform 1 0 21804 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_65_233
timestamp 1676037725
transform 1 0 22540 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_242
timestamp 1676037725
transform 1 0 23368 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_255
timestamp 1676037725
transform 1 0 24564 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_266
timestamp 1676037725
transform 1 0 25576 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_278
timestamp 1676037725
transform 1 0 26680 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1676037725
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_293
timestamp 1676037725
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_305
timestamp 1676037725
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_317
timestamp 1676037725
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1676037725
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1676037725
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_337
timestamp 1676037725
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_349
timestamp 1676037725
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_361
timestamp 1676037725
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_373
timestamp 1676037725
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1676037725
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1676037725
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1676037725
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1676037725
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1676037725
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1676037725
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1676037725
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1676037725
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1676037725
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1676037725
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1676037725
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1676037725
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1676037725
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1676037725
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_505
timestamp 1676037725
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_517
timestamp 1676037725
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_529
timestamp 1676037725
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_541
timestamp 1676037725
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 1676037725
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1676037725
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_561
timestamp 1676037725
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_573
timestamp 1676037725
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_585
timestamp 1676037725
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_597
timestamp 1676037725
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_609
timestamp 1676037725
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1676037725
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_617
timestamp 1676037725
transform 1 0 57868 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_623
timestamp 1676037725
transform 1 0 58420 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_3
timestamp 1676037725
transform 1 0 1380 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_66_9
timestamp 1676037725
transform 1 0 1932 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_15
timestamp 1676037725
transform 1 0 2484 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_21
timestamp 1676037725
transform 1 0 3036 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1676037725
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1676037725
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1676037725
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1676037725
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1676037725
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1676037725
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1676037725
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1676037725
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1676037725
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1676037725
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1676037725
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1676037725
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1676037725
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1676037725
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1676037725
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1676037725
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1676037725
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1676037725
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1676037725
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_197
timestamp 1676037725
transform 1 0 19228 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_205
timestamp 1676037725
transform 1 0 19964 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_213
timestamp 1676037725
transform 1 0 20700 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_219
timestamp 1676037725
transform 1 0 21252 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_230
timestamp 1676037725
transform 1 0 22264 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_247
timestamp 1676037725
transform 1 0 23828 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1676037725
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1676037725
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_265
timestamp 1676037725
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_277
timestamp 1676037725
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_289
timestamp 1676037725
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1676037725
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1676037725
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_309
timestamp 1676037725
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_321
timestamp 1676037725
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_333
timestamp 1676037725
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_345
timestamp 1676037725
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1676037725
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1676037725
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1676037725
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1676037725
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_389
timestamp 1676037725
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_401
timestamp 1676037725
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1676037725
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1676037725
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1676037725
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1676037725
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1676037725
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1676037725
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1676037725
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1676037725
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1676037725
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1676037725
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1676037725
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_513
timestamp 1676037725
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 1676037725
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1676037725
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_533
timestamp 1676037725
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_545
timestamp 1676037725
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_557
timestamp 1676037725
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_569
timestamp 1676037725
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_581
timestamp 1676037725
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 1676037725
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_589
timestamp 1676037725
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_601
timestamp 1676037725
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_613
timestamp 1676037725
transform 1 0 57500 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_623
timestamp 1676037725
transform 1 0 58420 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_3
timestamp 1676037725
transform 1 0 1380 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_9
timestamp 1676037725
transform 1 0 1932 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_21
timestamp 1676037725
transform 1 0 3036 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_33
timestamp 1676037725
transform 1 0 4140 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_45
timestamp 1676037725
transform 1 0 5244 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_53
timestamp 1676037725
transform 1 0 5980 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1676037725
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1676037725
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1676037725
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1676037725
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1676037725
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1676037725
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1676037725
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1676037725
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1676037725
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1676037725
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1676037725
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1676037725
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1676037725
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1676037725
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1676037725
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1676037725
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1676037725
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1676037725
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1676037725
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_245
timestamp 1676037725
transform 1 0 23644 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_257
timestamp 1676037725
transform 1 0 24748 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_269
timestamp 1676037725
transform 1 0 25852 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_277
timestamp 1676037725
transform 1 0 26588 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1676037725
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_293
timestamp 1676037725
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_305
timestamp 1676037725
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_317
timestamp 1676037725
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1676037725
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1676037725
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_337
timestamp 1676037725
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_349
timestamp 1676037725
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_361
timestamp 1676037725
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_373
timestamp 1676037725
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1676037725
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1676037725
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1676037725
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1676037725
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1676037725
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1676037725
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1676037725
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1676037725
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1676037725
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1676037725
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1676037725
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1676037725
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1676037725
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1676037725
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_505
timestamp 1676037725
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_517
timestamp 1676037725
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_529
timestamp 1676037725
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_541
timestamp 1676037725
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1676037725
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1676037725
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_561
timestamp 1676037725
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_573
timestamp 1676037725
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_585
timestamp 1676037725
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_597
timestamp 1676037725
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_609
timestamp 1676037725
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 1676037725
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_617
timestamp 1676037725
transform 1 0 57868 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_3
timestamp 1676037725
transform 1 0 1380 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_9
timestamp 1676037725
transform 1 0 1932 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_21
timestamp 1676037725
transform 1 0 3036 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1676037725
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1676037725
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1676037725
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1676037725
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1676037725
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1676037725
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1676037725
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1676037725
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1676037725
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1676037725
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1676037725
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1676037725
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1676037725
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1676037725
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1676037725
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1676037725
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1676037725
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1676037725
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1676037725
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1676037725
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1676037725
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1676037725
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_233
timestamp 1676037725
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1676037725
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1676037725
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1676037725
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1676037725
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_277
timestamp 1676037725
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_289
timestamp 1676037725
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1676037725
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1676037725
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 1676037725
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_321
timestamp 1676037725
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_333
timestamp 1676037725
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_345
timestamp 1676037725
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1676037725
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1676037725
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1676037725
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1676037725
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1676037725
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_401
timestamp 1676037725
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1676037725
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1676037725
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1676037725
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1676037725
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1676037725
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1676037725
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1676037725
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1676037725
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1676037725
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1676037725
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1676037725
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_513
timestamp 1676037725
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_525
timestamp 1676037725
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_531
timestamp 1676037725
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_533
timestamp 1676037725
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_545
timestamp 1676037725
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_557
timestamp 1676037725
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_569
timestamp 1676037725
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_581
timestamp 1676037725
transform 1 0 54556 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_587
timestamp 1676037725
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_589
timestamp 1676037725
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_601
timestamp 1676037725
transform 1 0 56396 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_613
timestamp 1676037725
transform 1 0 57500 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_623
timestamp 1676037725
transform 1 0 58420 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1676037725
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1676037725
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1676037725
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1676037725
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1676037725
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1676037725
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1676037725
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1676037725
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1676037725
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1676037725
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1676037725
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1676037725
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1676037725
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1676037725
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1676037725
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1676037725
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1676037725
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1676037725
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1676037725
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1676037725
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1676037725
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_205
timestamp 1676037725
transform 1 0 19964 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_213
timestamp 1676037725
transform 1 0 20700 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_222
timestamp 1676037725
transform 1 0 21528 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1676037725
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1676037725
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1676037725
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_261
timestamp 1676037725
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1676037725
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1676037725
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_281
timestamp 1676037725
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_293
timestamp 1676037725
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_305
timestamp 1676037725
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_317
timestamp 1676037725
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1676037725
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1676037725
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1676037725
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1676037725
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1676037725
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1676037725
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1676037725
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1676037725
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1676037725
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1676037725
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1676037725
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1676037725
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1676037725
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1676037725
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1676037725
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1676037725
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1676037725
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1676037725
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1676037725
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1676037725
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_505
timestamp 1676037725
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_517
timestamp 1676037725
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_529
timestamp 1676037725
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_541
timestamp 1676037725
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_553
timestamp 1676037725
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 1676037725
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_561
timestamp 1676037725
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_573
timestamp 1676037725
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_585
timestamp 1676037725
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_597
timestamp 1676037725
transform 1 0 56028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_609
timestamp 1676037725
transform 1 0 57132 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_615
timestamp 1676037725
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_617
timestamp 1676037725
transform 1 0 57868 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_3
timestamp 1676037725
transform 1 0 1380 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_9
timestamp 1676037725
transform 1 0 1932 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_21
timestamp 1676037725
transform 1 0 3036 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1676037725
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1676037725
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1676037725
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1676037725
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1676037725
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1676037725
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1676037725
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1676037725
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1676037725
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1676037725
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1676037725
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1676037725
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1676037725
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1676037725
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1676037725
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1676037725
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1676037725
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1676037725
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1676037725
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1676037725
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1676037725
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1676037725
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1676037725
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1676037725
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1676037725
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1676037725
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_265
timestamp 1676037725
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_277
timestamp 1676037725
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_289
timestamp 1676037725
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1676037725
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1676037725
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_309
timestamp 1676037725
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_321
timestamp 1676037725
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_333
timestamp 1676037725
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_345
timestamp 1676037725
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1676037725
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1676037725
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1676037725
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1676037725
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_389
timestamp 1676037725
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_401
timestamp 1676037725
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1676037725
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1676037725
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1676037725
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1676037725
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1676037725
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1676037725
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1676037725
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1676037725
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1676037725
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1676037725
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1676037725
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_513
timestamp 1676037725
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_525
timestamp 1676037725
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_531
timestamp 1676037725
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_533
timestamp 1676037725
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_545
timestamp 1676037725
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_557
timestamp 1676037725
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_569
timestamp 1676037725
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_581
timestamp 1676037725
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_587
timestamp 1676037725
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_589
timestamp 1676037725
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_601
timestamp 1676037725
transform 1 0 56396 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_70_613
timestamp 1676037725
transform 1 0 57500 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_623
timestamp 1676037725
transform 1 0 58420 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_3
timestamp 1676037725
transform 1 0 1380 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_9
timestamp 1676037725
transform 1 0 1932 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_21
timestamp 1676037725
transform 1 0 3036 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_33
timestamp 1676037725
transform 1 0 4140 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_45
timestamp 1676037725
transform 1 0 5244 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_53
timestamp 1676037725
transform 1 0 5980 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1676037725
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1676037725
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1676037725
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1676037725
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1676037725
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1676037725
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1676037725
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1676037725
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1676037725
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1676037725
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1676037725
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1676037725
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1676037725
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1676037725
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1676037725
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1676037725
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1676037725
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1676037725
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1676037725
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1676037725
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_249
timestamp 1676037725
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_261
timestamp 1676037725
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1676037725
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1676037725
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_281
timestamp 1676037725
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_293
timestamp 1676037725
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_305
timestamp 1676037725
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_317
timestamp 1676037725
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1676037725
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1676037725
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1676037725
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_349
timestamp 1676037725
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1676037725
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1676037725
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1676037725
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1676037725
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1676037725
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1676037725
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1676037725
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1676037725
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1676037725
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1676037725
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1676037725
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1676037725
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1676037725
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1676037725
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1676037725
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1676037725
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_505
timestamp 1676037725
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_517
timestamp 1676037725
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_529
timestamp 1676037725
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_541
timestamp 1676037725
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_553
timestamp 1676037725
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_559
timestamp 1676037725
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_561
timestamp 1676037725
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_573
timestamp 1676037725
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_585
timestamp 1676037725
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_597
timestamp 1676037725
transform 1 0 56028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_609
timestamp 1676037725
transform 1 0 57132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_615
timestamp 1676037725
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_617
timestamp 1676037725
transform 1 0 57868 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_3
timestamp 1676037725
transform 1 0 1380 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_11
timestamp 1676037725
transform 1 0 2116 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_23
timestamp 1676037725
transform 1 0 3220 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1676037725
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1676037725
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1676037725
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1676037725
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1676037725
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1676037725
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1676037725
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1676037725
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1676037725
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1676037725
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1676037725
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1676037725
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1676037725
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1676037725
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1676037725
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1676037725
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1676037725
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1676037725
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1676037725
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1676037725
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1676037725
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1676037725
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1676037725
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1676037725
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1676037725
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1676037725
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_265
timestamp 1676037725
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_277
timestamp 1676037725
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_289
timestamp 1676037725
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1676037725
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1676037725
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1676037725
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_321
timestamp 1676037725
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_333
timestamp 1676037725
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_345
timestamp 1676037725
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1676037725
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1676037725
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_365
timestamp 1676037725
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_377
timestamp 1676037725
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_389
timestamp 1676037725
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_401
timestamp 1676037725
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1676037725
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1676037725
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1676037725
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1676037725
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1676037725
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1676037725
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1676037725
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1676037725
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1676037725
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1676037725
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1676037725
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_513
timestamp 1676037725
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_525
timestamp 1676037725
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_531
timestamp 1676037725
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_533
timestamp 1676037725
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_545
timestamp 1676037725
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_557
timestamp 1676037725
transform 1 0 52348 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_569
timestamp 1676037725
transform 1 0 53452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_581
timestamp 1676037725
transform 1 0 54556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_587
timestamp 1676037725
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_589
timestamp 1676037725
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_601
timestamp 1676037725
transform 1 0 56396 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_613
timestamp 1676037725
transform 1 0 57500 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_623
timestamp 1676037725
transform 1 0 58420 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_3
timestamp 1676037725
transform 1 0 1380 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_9
timestamp 1676037725
transform 1 0 1932 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_21
timestamp 1676037725
transform 1 0 3036 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_33
timestamp 1676037725
transform 1 0 4140 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_45
timestamp 1676037725
transform 1 0 5244 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_53
timestamp 1676037725
transform 1 0 5980 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1676037725
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1676037725
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1676037725
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1676037725
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1676037725
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1676037725
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1676037725
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1676037725
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1676037725
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1676037725
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1676037725
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1676037725
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1676037725
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1676037725
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1676037725
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1676037725
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1676037725
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1676037725
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1676037725
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1676037725
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1676037725
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_261
timestamp 1676037725
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1676037725
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1676037725
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_281
timestamp 1676037725
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_293
timestamp 1676037725
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_305
timestamp 1676037725
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_317
timestamp 1676037725
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1676037725
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1676037725
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1676037725
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_349
timestamp 1676037725
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_361
timestamp 1676037725
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_373
timestamp 1676037725
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1676037725
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1676037725
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1676037725
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1676037725
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1676037725
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1676037725
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1676037725
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1676037725
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1676037725
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1676037725
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1676037725
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1676037725
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1676037725
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1676037725
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_505
timestamp 1676037725
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_517
timestamp 1676037725
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_529
timestamp 1676037725
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_541
timestamp 1676037725
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_553
timestamp 1676037725
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_559
timestamp 1676037725
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_561
timestamp 1676037725
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_573
timestamp 1676037725
transform 1 0 53820 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_585
timestamp 1676037725
transform 1 0 54924 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_597
timestamp 1676037725
transform 1 0 56028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_609
timestamp 1676037725
transform 1 0 57132 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_615
timestamp 1676037725
transform 1 0 57684 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_617
timestamp 1676037725
transform 1 0 57868 0 -1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1676037725
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1676037725
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1676037725
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1676037725
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1676037725
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1676037725
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1676037725
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1676037725
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1676037725
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1676037725
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1676037725
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1676037725
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1676037725
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1676037725
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1676037725
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1676037725
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1676037725
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1676037725
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1676037725
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1676037725
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1676037725
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1676037725
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1676037725
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1676037725
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1676037725
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1676037725
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1676037725
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1676037725
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_265
timestamp 1676037725
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_277
timestamp 1676037725
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_289
timestamp 1676037725
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1676037725
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1676037725
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1676037725
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1676037725
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_333
timestamp 1676037725
transform 1 0 31740 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_341
timestamp 1676037725
transform 1 0 32476 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_359
timestamp 1676037725
transform 1 0 34132 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1676037725
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_365
timestamp 1676037725
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_377
timestamp 1676037725
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_389
timestamp 1676037725
transform 1 0 36892 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_400
timestamp 1676037725
transform 1 0 37904 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_412
timestamp 1676037725
transform 1 0 39008 0 1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1676037725
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1676037725
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1676037725
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1676037725
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1676037725
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1676037725
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1676037725
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1676037725
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1676037725
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_513
timestamp 1676037725
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_525
timestamp 1676037725
transform 1 0 49404 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_531
timestamp 1676037725
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_533
timestamp 1676037725
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_545
timestamp 1676037725
transform 1 0 51244 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_557
timestamp 1676037725
transform 1 0 52348 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_569
timestamp 1676037725
transform 1 0 53452 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_581
timestamp 1676037725
transform 1 0 54556 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_587
timestamp 1676037725
transform 1 0 55108 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_589
timestamp 1676037725
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_601
timestamp 1676037725
transform 1 0 56396 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_613
timestamp 1676037725
transform 1 0 57500 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_623
timestamp 1676037725
transform 1 0 58420 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_3
timestamp 1676037725
transform 1 0 1380 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_9
timestamp 1676037725
transform 1 0 1932 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_21
timestamp 1676037725
transform 1 0 3036 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_33
timestamp 1676037725
transform 1 0 4140 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_45
timestamp 1676037725
transform 1 0 5244 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_53
timestamp 1676037725
transform 1 0 5980 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1676037725
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1676037725
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1676037725
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1676037725
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1676037725
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1676037725
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1676037725
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1676037725
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1676037725
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1676037725
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1676037725
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1676037725
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1676037725
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1676037725
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1676037725
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1676037725
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1676037725
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1676037725
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1676037725
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1676037725
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1676037725
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_261
timestamp 1676037725
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1676037725
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1676037725
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1676037725
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_293
timestamp 1676037725
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_305
timestamp 1676037725
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_317
timestamp 1676037725
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1676037725
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1676037725
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_337
timestamp 1676037725
transform 1 0 32108 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_347
timestamp 1676037725
transform 1 0 33028 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_359
timestamp 1676037725
transform 1 0 34132 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_371
timestamp 1676037725
transform 1 0 35236 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_383
timestamp 1676037725
transform 1 0 36340 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1676037725
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1676037725
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1676037725
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1676037725
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1676037725
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1676037725
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1676037725
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1676037725
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1676037725
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1676037725
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1676037725
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1676037725
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1676037725
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_505
timestamp 1676037725
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_517
timestamp 1676037725
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_529
timestamp 1676037725
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_541
timestamp 1676037725
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_553
timestamp 1676037725
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_559
timestamp 1676037725
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_561
timestamp 1676037725
transform 1 0 52716 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_573
timestamp 1676037725
transform 1 0 53820 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_585
timestamp 1676037725
transform 1 0 54924 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_597
timestamp 1676037725
transform 1 0 56028 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_609
timestamp 1676037725
transform 1 0 57132 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_615
timestamp 1676037725
transform 1 0 57684 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_617
timestamp 1676037725
transform 1 0 57868 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_3
timestamp 1676037725
transform 1 0 1380 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_9
timestamp 1676037725
transform 1 0 1932 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_21
timestamp 1676037725
transform 1 0 3036 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1676037725
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1676037725
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1676037725
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1676037725
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1676037725
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1676037725
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1676037725
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1676037725
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1676037725
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1676037725
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1676037725
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1676037725
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1676037725
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1676037725
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1676037725
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1676037725
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1676037725
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1676037725
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1676037725
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1676037725
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1676037725
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_221
timestamp 1676037725
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1676037725
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1676037725
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1676037725
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1676037725
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_265
timestamp 1676037725
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_277
timestamp 1676037725
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_289
timestamp 1676037725
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1676037725
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1676037725
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_309
timestamp 1676037725
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_321
timestamp 1676037725
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_333
timestamp 1676037725
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_345
timestamp 1676037725
transform 1 0 32844 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_353
timestamp 1676037725
transform 1 0 33580 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_362
timestamp 1676037725
transform 1 0 34408 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1676037725
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_377
timestamp 1676037725
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_389
timestamp 1676037725
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_401
timestamp 1676037725
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1676037725
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1676037725
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1676037725
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1676037725
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1676037725
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1676037725
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1676037725
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1676037725
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1676037725
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1676037725
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1676037725
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_513
timestamp 1676037725
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_525
timestamp 1676037725
transform 1 0 49404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_531
timestamp 1676037725
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_533
timestamp 1676037725
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_545
timestamp 1676037725
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_557
timestamp 1676037725
transform 1 0 52348 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_569
timestamp 1676037725
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_581
timestamp 1676037725
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_587
timestamp 1676037725
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_589
timestamp 1676037725
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_601
timestamp 1676037725
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_613
timestamp 1676037725
transform 1 0 57500 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_623
timestamp 1676037725
transform 1 0 58420 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_3
timestamp 1676037725
transform 1 0 1380 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_9
timestamp 1676037725
transform 1 0 1932 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_21
timestamp 1676037725
transform 1 0 3036 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_33
timestamp 1676037725
transform 1 0 4140 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_45
timestamp 1676037725
transform 1 0 5244 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_53
timestamp 1676037725
transform 1 0 5980 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1676037725
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1676037725
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1676037725
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1676037725
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1676037725
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1676037725
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1676037725
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1676037725
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1676037725
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1676037725
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1676037725
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1676037725
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1676037725
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1676037725
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1676037725
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1676037725
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1676037725
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1676037725
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1676037725
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1676037725
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_249
timestamp 1676037725
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_261
timestamp 1676037725
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1676037725
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1676037725
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1676037725
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1676037725
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1676037725
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1676037725
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1676037725
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1676037725
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1676037725
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_349
timestamp 1676037725
transform 1 0 33212 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_357
timestamp 1676037725
transform 1 0 33948 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_366
timestamp 1676037725
transform 1 0 34776 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_378
timestamp 1676037725
transform 1 0 35880 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_390
timestamp 1676037725
transform 1 0 36984 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1676037725
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_405
timestamp 1676037725
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_417
timestamp 1676037725
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_429
timestamp 1676037725
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1676037725
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1676037725
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1676037725
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1676037725
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1676037725
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1676037725
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1676037725
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1676037725
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_505
timestamp 1676037725
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_517
timestamp 1676037725
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_529
timestamp 1676037725
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_541
timestamp 1676037725
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_553
timestamp 1676037725
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_559
timestamp 1676037725
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_561
timestamp 1676037725
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_573
timestamp 1676037725
transform 1 0 53820 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_585
timestamp 1676037725
transform 1 0 54924 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_597
timestamp 1676037725
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_609
timestamp 1676037725
transform 1 0 57132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_615
timestamp 1676037725
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_617
timestamp 1676037725
transform 1 0 57868 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_3
timestamp 1676037725
transform 1 0 1380 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_11
timestamp 1676037725
transform 1 0 2116 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_23
timestamp 1676037725
transform 1 0 3220 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1676037725
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1676037725
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1676037725
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1676037725
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1676037725
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1676037725
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1676037725
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1676037725
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1676037725
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1676037725
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1676037725
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1676037725
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1676037725
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1676037725
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1676037725
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1676037725
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1676037725
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1676037725
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1676037725
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1676037725
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1676037725
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1676037725
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1676037725
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1676037725
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1676037725
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1676037725
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1676037725
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_277
timestamp 1676037725
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_289
timestamp 1676037725
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1676037725
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1676037725
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1676037725
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1676037725
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1676037725
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1676037725
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1676037725
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1676037725
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_365
timestamp 1676037725
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_377
timestamp 1676037725
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_389
timestamp 1676037725
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_401
timestamp 1676037725
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1676037725
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1676037725
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1676037725
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1676037725
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1676037725
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1676037725
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1676037725
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1676037725
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1676037725
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1676037725
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1676037725
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_513
timestamp 1676037725
transform 1 0 48300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_525
timestamp 1676037725
transform 1 0 49404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_531
timestamp 1676037725
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_533
timestamp 1676037725
transform 1 0 50140 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_545
timestamp 1676037725
transform 1 0 51244 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_557
timestamp 1676037725
transform 1 0 52348 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_569
timestamp 1676037725
transform 1 0 53452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_581
timestamp 1676037725
transform 1 0 54556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_587
timestamp 1676037725
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_589
timestamp 1676037725
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_601
timestamp 1676037725
transform 1 0 56396 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_78_613
timestamp 1676037725
transform 1 0 57500 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_623
timestamp 1676037725
transform 1 0 58420 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1676037725
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1676037725
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1676037725
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1676037725
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1676037725
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1676037725
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1676037725
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1676037725
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1676037725
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1676037725
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1676037725
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1676037725
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1676037725
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1676037725
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1676037725
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1676037725
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1676037725
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1676037725
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_169
timestamp 1676037725
transform 1 0 16652 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_182
timestamp 1676037725
transform 1 0 17848 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_194
timestamp 1676037725
transform 1 0 18952 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_206
timestamp 1676037725
transform 1 0 20056 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_218
timestamp 1676037725
transform 1 0 21160 0 -1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1676037725
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1676037725
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1676037725
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_261
timestamp 1676037725
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1676037725
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1676037725
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1676037725
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1676037725
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_305
timestamp 1676037725
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_317
timestamp 1676037725
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1676037725
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1676037725
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_337
timestamp 1676037725
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_349
timestamp 1676037725
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1676037725
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_373
timestamp 1676037725
transform 1 0 35420 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_381
timestamp 1676037725
transform 1 0 36156 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_390
timestamp 1676037725
transform 1 0 36984 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_393
timestamp 1676037725
transform 1 0 37260 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_399
timestamp 1676037725
transform 1 0 37812 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_409
timestamp 1676037725
transform 1 0 38732 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_421
timestamp 1676037725
transform 1 0 39836 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_433
timestamp 1676037725
transform 1 0 40940 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_445
timestamp 1676037725
transform 1 0 42044 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1676037725
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1676037725
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1676037725
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1676037725
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1676037725
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1676037725
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_505
timestamp 1676037725
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_517
timestamp 1676037725
transform 1 0 48668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_529
timestamp 1676037725
transform 1 0 49772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_541
timestamp 1676037725
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_553
timestamp 1676037725
transform 1 0 51980 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_559
timestamp 1676037725
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_561
timestamp 1676037725
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_573
timestamp 1676037725
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_585
timestamp 1676037725
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_597
timestamp 1676037725
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_609
timestamp 1676037725
transform 1 0 57132 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_615
timestamp 1676037725
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_617
timestamp 1676037725
transform 1 0 57868 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_623
timestamp 1676037725
transform 1 0 58420 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_3
timestamp 1676037725
transform 1 0 1380 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_9
timestamp 1676037725
transform 1 0 1932 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_21
timestamp 1676037725
transform 1 0 3036 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1676037725
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1676037725
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1676037725
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1676037725
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1676037725
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1676037725
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1676037725
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1676037725
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1676037725
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1676037725
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1676037725
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1676037725
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1676037725
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1676037725
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1676037725
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1676037725
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_177
timestamp 1676037725
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1676037725
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1676037725
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1676037725
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1676037725
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1676037725
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_233
timestamp 1676037725
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1676037725
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1676037725
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_253
timestamp 1676037725
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_265
timestamp 1676037725
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_277
timestamp 1676037725
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_289
timestamp 1676037725
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1676037725
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1676037725
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_309
timestamp 1676037725
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_321
timestamp 1676037725
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_333
timestamp 1676037725
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_345
timestamp 1676037725
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1676037725
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1676037725
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_365
timestamp 1676037725
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_377
timestamp 1676037725
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_389
timestamp 1676037725
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_401
timestamp 1676037725
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_413
timestamp 1676037725
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1676037725
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1676037725
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1676037725
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1676037725
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1676037725
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1676037725
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1676037725
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1676037725
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1676037725
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_501
timestamp 1676037725
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_513
timestamp 1676037725
transform 1 0 48300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_525
timestamp 1676037725
transform 1 0 49404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_531
timestamp 1676037725
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_533
timestamp 1676037725
transform 1 0 50140 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_545
timestamp 1676037725
transform 1 0 51244 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_557
timestamp 1676037725
transform 1 0 52348 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_569
timestamp 1676037725
transform 1 0 53452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_581
timestamp 1676037725
transform 1 0 54556 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_587
timestamp 1676037725
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_589
timestamp 1676037725
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_601
timestamp 1676037725
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_613
timestamp 1676037725
transform 1 0 57500 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_623
timestamp 1676037725
transform 1 0 58420 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_3
timestamp 1676037725
transform 1 0 1380 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_9
timestamp 1676037725
transform 1 0 1932 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_21
timestamp 1676037725
transform 1 0 3036 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_33
timestamp 1676037725
transform 1 0 4140 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_45
timestamp 1676037725
transform 1 0 5244 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_53
timestamp 1676037725
transform 1 0 5980 0 -1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1676037725
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1676037725
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1676037725
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1676037725
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1676037725
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1676037725
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1676037725
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1676037725
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1676037725
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1676037725
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1676037725
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1676037725
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1676037725
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1676037725
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1676037725
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1676037725
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1676037725
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1676037725
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1676037725
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1676037725
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1676037725
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_261
timestamp 1676037725
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1676037725
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1676037725
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1676037725
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_293
timestamp 1676037725
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_305
timestamp 1676037725
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_317
timestamp 1676037725
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1676037725
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1676037725
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_337
timestamp 1676037725
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_349
timestamp 1676037725
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_361
timestamp 1676037725
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_373
timestamp 1676037725
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1676037725
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1676037725
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1676037725
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1676037725
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1676037725
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1676037725
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1676037725
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1676037725
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1676037725
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1676037725
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1676037725
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 1676037725
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1676037725
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1676037725
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_505
timestamp 1676037725
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_517
timestamp 1676037725
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_529
timestamp 1676037725
transform 1 0 49772 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_541
timestamp 1676037725
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_553
timestamp 1676037725
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_559
timestamp 1676037725
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_561
timestamp 1676037725
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_573
timestamp 1676037725
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_585
timestamp 1676037725
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_597
timestamp 1676037725
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_609
timestamp 1676037725
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_615
timestamp 1676037725
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_617
timestamp 1676037725
transform 1 0 57868 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_3
timestamp 1676037725
transform 1 0 1380 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_9
timestamp 1676037725
transform 1 0 1932 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_21
timestamp 1676037725
transform 1 0 3036 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1676037725
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1676037725
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1676037725
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1676037725
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1676037725
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1676037725
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1676037725
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1676037725
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1676037725
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_109
timestamp 1676037725
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_121
timestamp 1676037725
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1676037725
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1676037725
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1676037725
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1676037725
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1676037725
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1676037725
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1676037725
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1676037725
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1676037725
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1676037725
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1676037725
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1676037725
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1676037725
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1676037725
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_253
timestamp 1676037725
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_265
timestamp 1676037725
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_277
timestamp 1676037725
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_289
timestamp 1676037725
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1676037725
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1676037725
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_309
timestamp 1676037725
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_321
timestamp 1676037725
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_333
timestamp 1676037725
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_345
timestamp 1676037725
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1676037725
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1676037725
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1676037725
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_377
timestamp 1676037725
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_389
timestamp 1676037725
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_401
timestamp 1676037725
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1676037725
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1676037725
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1676037725
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1676037725
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_445
timestamp 1676037725
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_457
timestamp 1676037725
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1676037725
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1676037725
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 1676037725
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_489
timestamp 1676037725
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_501
timestamp 1676037725
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_513
timestamp 1676037725
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_525
timestamp 1676037725
transform 1 0 49404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_531
timestamp 1676037725
transform 1 0 49956 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_533
timestamp 1676037725
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_545
timestamp 1676037725
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_557
timestamp 1676037725
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_569
timestamp 1676037725
transform 1 0 53452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_581
timestamp 1676037725
transform 1 0 54556 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_587
timestamp 1676037725
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_589
timestamp 1676037725
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_601
timestamp 1676037725
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_613
timestamp 1676037725
transform 1 0 57500 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_83_3
timestamp 1676037725
transform 1 0 1380 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_9
timestamp 1676037725
transform 1 0 1932 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_21
timestamp 1676037725
transform 1 0 3036 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_33
timestamp 1676037725
transform 1 0 4140 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_45
timestamp 1676037725
transform 1 0 5244 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_53
timestamp 1676037725
transform 1 0 5980 0 -1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1676037725
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1676037725
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1676037725
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_93
timestamp 1676037725
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1676037725
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1676037725
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1676037725
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1676037725
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1676037725
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1676037725
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1676037725
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1676037725
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1676037725
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1676037725
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1676037725
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1676037725
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1676037725
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1676037725
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1676037725
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1676037725
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_249
timestamp 1676037725
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_261
timestamp 1676037725
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_273
timestamp 1676037725
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 1676037725
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_281
timestamp 1676037725
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_293
timestamp 1676037725
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_305
timestamp 1676037725
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_317
timestamp 1676037725
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1676037725
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1676037725
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_337
timestamp 1676037725
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_349
timestamp 1676037725
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_361
timestamp 1676037725
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_373
timestamp 1676037725
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_385
timestamp 1676037725
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1676037725
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_393
timestamp 1676037725
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_405
timestamp 1676037725
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_417
timestamp 1676037725
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_429
timestamp 1676037725
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_441
timestamp 1676037725
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1676037725
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_449
timestamp 1676037725
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_461
timestamp 1676037725
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_473
timestamp 1676037725
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_485
timestamp 1676037725
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_497
timestamp 1676037725
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1676037725
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_505
timestamp 1676037725
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_517
timestamp 1676037725
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_529
timestamp 1676037725
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_541
timestamp 1676037725
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_553
timestamp 1676037725
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_559
timestamp 1676037725
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_561
timestamp 1676037725
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_573
timestamp 1676037725
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_585
timestamp 1676037725
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_597
timestamp 1676037725
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_609
timestamp 1676037725
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_615
timestamp 1676037725
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_617
timestamp 1676037725
transform 1 0 57868 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_623
timestamp 1676037725
transform 1 0 58420 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_84_3
timestamp 1676037725
transform 1 0 1380 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_9
timestamp 1676037725
transform 1 0 1932 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_18
timestamp 1676037725
transform 1 0 2760 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_26
timestamp 1676037725
transform 1 0 3496 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1676037725
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1676037725
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1676037725
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1676037725
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1676037725
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1676037725
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1676037725
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1676037725
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1676037725
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1676037725
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1676037725
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1676037725
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1676037725
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1676037725
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1676037725
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1676037725
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1676037725
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1676037725
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1676037725
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1676037725
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1676037725
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1676037725
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1676037725
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1676037725
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_253
timestamp 1676037725
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_265
timestamp 1676037725
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_277
timestamp 1676037725
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_289
timestamp 1676037725
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 1676037725
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1676037725
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_309
timestamp 1676037725
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_321
timestamp 1676037725
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_333
timestamp 1676037725
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_345
timestamp 1676037725
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_357
timestamp 1676037725
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1676037725
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_365
timestamp 1676037725
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_377
timestamp 1676037725
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_389
timestamp 1676037725
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_401
timestamp 1676037725
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_413
timestamp 1676037725
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1676037725
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_421
timestamp 1676037725
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_433
timestamp 1676037725
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_445
timestamp 1676037725
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_457
timestamp 1676037725
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1676037725
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1676037725
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_477
timestamp 1676037725
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_489
timestamp 1676037725
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_501
timestamp 1676037725
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_513
timestamp 1676037725
transform 1 0 48300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_525
timestamp 1676037725
transform 1 0 49404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_531
timestamp 1676037725
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_533
timestamp 1676037725
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_545
timestamp 1676037725
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_557
timestamp 1676037725
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_569
timestamp 1676037725
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_581
timestamp 1676037725
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_587
timestamp 1676037725
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_589
timestamp 1676037725
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_601
timestamp 1676037725
transform 1 0 56396 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_613
timestamp 1676037725
transform 1 0 57500 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_84_623
timestamp 1676037725
transform 1 0 58420 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_3
timestamp 1676037725
transform 1 0 1380 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_9
timestamp 1676037725
transform 1 0 1932 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_21
timestamp 1676037725
transform 1 0 3036 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_33
timestamp 1676037725
transform 1 0 4140 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_45
timestamp 1676037725
transform 1 0 5244 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_85_53
timestamp 1676037725
transform 1 0 5980 0 -1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1676037725
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1676037725
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1676037725
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1676037725
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1676037725
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1676037725
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1676037725
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1676037725
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1676037725
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1676037725
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1676037725
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1676037725
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1676037725
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1676037725
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1676037725
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1676037725
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1676037725
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1676037725
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1676037725
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1676037725
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1676037725
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_261
timestamp 1676037725
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 1676037725
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1676037725
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_281
timestamp 1676037725
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_293
timestamp 1676037725
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_305
timestamp 1676037725
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_317
timestamp 1676037725
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_329
timestamp 1676037725
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1676037725
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_337
timestamp 1676037725
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_349
timestamp 1676037725
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_361
timestamp 1676037725
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_373
timestamp 1676037725
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 1676037725
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1676037725
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_393
timestamp 1676037725
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_405
timestamp 1676037725
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_417
timestamp 1676037725
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_429
timestamp 1676037725
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 1676037725
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1676037725
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_449
timestamp 1676037725
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_461
timestamp 1676037725
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_473
timestamp 1676037725
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_485
timestamp 1676037725
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 1676037725
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1676037725
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_505
timestamp 1676037725
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_517
timestamp 1676037725
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_529
timestamp 1676037725
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_541
timestamp 1676037725
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_553
timestamp 1676037725
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_559
timestamp 1676037725
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_561
timestamp 1676037725
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_573
timestamp 1676037725
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_585
timestamp 1676037725
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_597
timestamp 1676037725
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_609
timestamp 1676037725
transform 1 0 57132 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_615
timestamp 1676037725
transform 1 0 57684 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_617
timestamp 1676037725
transform 1 0 57868 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_3
timestamp 1676037725
transform 1 0 1380 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_9
timestamp 1676037725
transform 1 0 1932 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_21
timestamp 1676037725
transform 1 0 3036 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1676037725
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1676037725
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1676037725
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1676037725
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1676037725
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1676037725
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1676037725
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1676037725
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1676037725
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1676037725
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1676037725
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1676037725
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1676037725
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1676037725
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1676037725
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1676037725
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1676037725
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1676037725
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1676037725
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1676037725
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1676037725
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1676037725
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1676037725
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1676037725
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1676037725
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_253
timestamp 1676037725
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_265
timestamp 1676037725
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_277
timestamp 1676037725
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_289
timestamp 1676037725
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 1676037725
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1676037725
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_309
timestamp 1676037725
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_321
timestamp 1676037725
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_333
timestamp 1676037725
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_345
timestamp 1676037725
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_357
timestamp 1676037725
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1676037725
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_365
timestamp 1676037725
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_377
timestamp 1676037725
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_389
timestamp 1676037725
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_401
timestamp 1676037725
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_413
timestamp 1676037725
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1676037725
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1676037725
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1676037725
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_445
timestamp 1676037725
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_457
timestamp 1676037725
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1676037725
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1676037725
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_477
timestamp 1676037725
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_489
timestamp 1676037725
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_501
timestamp 1676037725
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_513
timestamp 1676037725
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_525
timestamp 1676037725
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_531
timestamp 1676037725
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_533
timestamp 1676037725
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_545
timestamp 1676037725
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_557
timestamp 1676037725
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_569
timestamp 1676037725
transform 1 0 53452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_581
timestamp 1676037725
transform 1 0 54556 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_587
timestamp 1676037725
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_589
timestamp 1676037725
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_601
timestamp 1676037725
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_613
timestamp 1676037725
transform 1 0 57500 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_623
timestamp 1676037725
transform 1 0 58420 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_3
timestamp 1676037725
transform 1 0 1380 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_9
timestamp 1676037725
transform 1 0 1932 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_21
timestamp 1676037725
transform 1 0 3036 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_33
timestamp 1676037725
transform 1 0 4140 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_45
timestamp 1676037725
transform 1 0 5244 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_87_53
timestamp 1676037725
transform 1 0 5980 0 -1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1676037725
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1676037725
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1676037725
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1676037725
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1676037725
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1676037725
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1676037725
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1676037725
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1676037725
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1676037725
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1676037725
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1676037725
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1676037725
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1676037725
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1676037725
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1676037725
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1676037725
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1676037725
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1676037725
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1676037725
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_249
timestamp 1676037725
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_261
timestamp 1676037725
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_273
timestamp 1676037725
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1676037725
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_281
timestamp 1676037725
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_293
timestamp 1676037725
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_305
timestamp 1676037725
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_317
timestamp 1676037725
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 1676037725
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1676037725
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_337
timestamp 1676037725
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_349
timestamp 1676037725
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_361
timestamp 1676037725
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_373
timestamp 1676037725
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 1676037725
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1676037725
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_393
timestamp 1676037725
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_405
timestamp 1676037725
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_417
timestamp 1676037725
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_429
timestamp 1676037725
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1676037725
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1676037725
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_449
timestamp 1676037725
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_461
timestamp 1676037725
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_473
timestamp 1676037725
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_485
timestamp 1676037725
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1676037725
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1676037725
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_505
timestamp 1676037725
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_517
timestamp 1676037725
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_529
timestamp 1676037725
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_541
timestamp 1676037725
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_553
timestamp 1676037725
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_559
timestamp 1676037725
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_561
timestamp 1676037725
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_573
timestamp 1676037725
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_585
timestamp 1676037725
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_597
timestamp 1676037725
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_609
timestamp 1676037725
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_615
timestamp 1676037725
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_617
timestamp 1676037725
transform 1 0 57868 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_3
timestamp 1676037725
transform 1 0 1380 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_9
timestamp 1676037725
transform 1 0 1932 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_21
timestamp 1676037725
transform 1 0 3036 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1676037725
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1676037725
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1676037725
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1676037725
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1676037725
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1676037725
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1676037725
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1676037725
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1676037725
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1676037725
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1676037725
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1676037725
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1676037725
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1676037725
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1676037725
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1676037725
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1676037725
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1676037725
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1676037725
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1676037725
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1676037725
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1676037725
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1676037725
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1676037725
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1676037725
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_253
timestamp 1676037725
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_265
timestamp 1676037725
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_277
timestamp 1676037725
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_289
timestamp 1676037725
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_301
timestamp 1676037725
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1676037725
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_309
timestamp 1676037725
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_321
timestamp 1676037725
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_333
timestamp 1676037725
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_345
timestamp 1676037725
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 1676037725
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1676037725
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_365
timestamp 1676037725
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_377
timestamp 1676037725
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_389
timestamp 1676037725
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_401
timestamp 1676037725
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1676037725
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1676037725
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1676037725
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1676037725
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_445
timestamp 1676037725
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_457
timestamp 1676037725
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1676037725
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1676037725
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_477
timestamp 1676037725
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_489
timestamp 1676037725
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_501
timestamp 1676037725
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_513
timestamp 1676037725
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_525
timestamp 1676037725
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_531
timestamp 1676037725
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_533
timestamp 1676037725
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_545
timestamp 1676037725
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_557
timestamp 1676037725
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_569
timestamp 1676037725
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_581
timestamp 1676037725
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_587
timestamp 1676037725
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_589
timestamp 1676037725
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_601
timestamp 1676037725
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_613
timestamp 1676037725
transform 1 0 57500 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_88_623
timestamp 1676037725
transform 1 0 58420 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1676037725
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1676037725
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_89_27
timestamp 1676037725
transform 1 0 3588 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_36
timestamp 1676037725
transform 1 0 4416 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_48
timestamp 1676037725
transform 1 0 5520 0 -1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1676037725
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1676037725
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1676037725
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1676037725
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1676037725
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1676037725
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1676037725
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1676037725
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1676037725
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1676037725
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1676037725
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1676037725
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1676037725
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1676037725
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1676037725
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1676037725
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1676037725
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1676037725
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1676037725
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1676037725
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_249
timestamp 1676037725
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_261
timestamp 1676037725
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_273
timestamp 1676037725
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1676037725
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_281
timestamp 1676037725
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_293
timestamp 1676037725
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_305
timestamp 1676037725
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_317
timestamp 1676037725
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1676037725
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1676037725
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_337
timestamp 1676037725
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_349
timestamp 1676037725
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_361
timestamp 1676037725
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_373
timestamp 1676037725
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1676037725
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1676037725
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_393
timestamp 1676037725
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_405
timestamp 1676037725
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_417
timestamp 1676037725
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_429
timestamp 1676037725
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1676037725
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1676037725
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_449
timestamp 1676037725
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_461
timestamp 1676037725
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_473
timestamp 1676037725
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_485
timestamp 1676037725
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1676037725
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1676037725
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_505
timestamp 1676037725
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_517
timestamp 1676037725
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_529
timestamp 1676037725
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_541
timestamp 1676037725
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_553
timestamp 1676037725
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_559
timestamp 1676037725
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_561
timestamp 1676037725
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_573
timestamp 1676037725
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_585
timestamp 1676037725
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_597
timestamp 1676037725
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_609
timestamp 1676037725
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_615
timestamp 1676037725
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_617
timestamp 1676037725
transform 1 0 57868 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_90_3
timestamp 1676037725
transform 1 0 1380 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_9
timestamp 1676037725
transform 1 0 1932 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_21
timestamp 1676037725
transform 1 0 3036 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1676037725
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1676037725
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1676037725
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1676037725
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1676037725
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1676037725
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1676037725
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1676037725
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1676037725
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1676037725
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1676037725
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1676037725
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1676037725
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1676037725
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1676037725
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1676037725
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1676037725
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1676037725
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1676037725
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1676037725
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_90_209
timestamp 1676037725
transform 1 0 20332 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_220
timestamp 1676037725
transform 1 0 21344 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_232
timestamp 1676037725
transform 1 0 22448 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_244
timestamp 1676037725
transform 1 0 23552 0 1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_90_253
timestamp 1676037725
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_265
timestamp 1676037725
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_277
timestamp 1676037725
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_289
timestamp 1676037725
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_301
timestamp 1676037725
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1676037725
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_309
timestamp 1676037725
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_321
timestamp 1676037725
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_333
timestamp 1676037725
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_345
timestamp 1676037725
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 1676037725
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1676037725
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_365
timestamp 1676037725
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_377
timestamp 1676037725
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_389
timestamp 1676037725
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_401
timestamp 1676037725
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1676037725
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1676037725
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1676037725
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_433
timestamp 1676037725
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_445
timestamp 1676037725
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_457
timestamp 1676037725
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1676037725
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1676037725
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_477
timestamp 1676037725
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_489
timestamp 1676037725
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_501
timestamp 1676037725
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_513
timestamp 1676037725
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_525
timestamp 1676037725
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_531
timestamp 1676037725
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_533
timestamp 1676037725
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_545
timestamp 1676037725
transform 1 0 51244 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_557
timestamp 1676037725
transform 1 0 52348 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_569
timestamp 1676037725
transform 1 0 53452 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_581
timestamp 1676037725
transform 1 0 54556 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_587
timestamp 1676037725
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_589
timestamp 1676037725
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_601
timestamp 1676037725
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_613
timestamp 1676037725
transform 1 0 57500 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_619
timestamp 1676037725
transform 1 0 58052 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_623
timestamp 1676037725
transform 1 0 58420 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_3
timestamp 1676037725
transform 1 0 1380 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_9
timestamp 1676037725
transform 1 0 1932 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_21
timestamp 1676037725
transform 1 0 3036 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_33
timestamp 1676037725
transform 1 0 4140 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_45
timestamp 1676037725
transform 1 0 5244 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_91_53
timestamp 1676037725
transform 1 0 5980 0 -1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1676037725
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_91_69
timestamp 1676037725
transform 1 0 7452 0 -1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_91_79
timestamp 1676037725
transform 1 0 8372 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_91
timestamp 1676037725
transform 1 0 9476 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_103
timestamp 1676037725
transform 1 0 10580 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1676037725
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1676037725
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1676037725
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1676037725
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1676037725
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1676037725
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1676037725
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1676037725
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1676037725
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1676037725
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1676037725
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1676037725
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1676037725
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1676037725
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1676037725
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1676037725
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_261
timestamp 1676037725
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 1676037725
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1676037725
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_281
timestamp 1676037725
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_293
timestamp 1676037725
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_305
timestamp 1676037725
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_317
timestamp 1676037725
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 1676037725
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1676037725
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_337
timestamp 1676037725
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_349
timestamp 1676037725
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_361
timestamp 1676037725
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_373
timestamp 1676037725
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1676037725
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1676037725
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_393
timestamp 1676037725
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_405
timestamp 1676037725
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_417
timestamp 1676037725
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_429
timestamp 1676037725
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1676037725
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1676037725
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_449
timestamp 1676037725
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_461
timestamp 1676037725
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_473
timestamp 1676037725
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_485
timestamp 1676037725
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1676037725
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1676037725
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_505
timestamp 1676037725
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_517
timestamp 1676037725
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_529
timestamp 1676037725
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_541
timestamp 1676037725
transform 1 0 50876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_553
timestamp 1676037725
transform 1 0 51980 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_559
timestamp 1676037725
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_561
timestamp 1676037725
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_573
timestamp 1676037725
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_585
timestamp 1676037725
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_597
timestamp 1676037725
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_609
timestamp 1676037725
transform 1 0 57132 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_615
timestamp 1676037725
transform 1 0 57684 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_617
timestamp 1676037725
transform 1 0 57868 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_92_3
timestamp 1676037725
transform 1 0 1380 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_11
timestamp 1676037725
transform 1 0 2116 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_23
timestamp 1676037725
transform 1 0 3220 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1676037725
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1676037725
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1676037725
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1676037725
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_65
timestamp 1676037725
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1676037725
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1676037725
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1676037725
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1676037725
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1676037725
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1676037725
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1676037725
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1676037725
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1676037725
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1676037725
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1676037725
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1676037725
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1676037725
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1676037725
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1676037725
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1676037725
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1676037725
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1676037725
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1676037725
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1676037725
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_253
timestamp 1676037725
transform 1 0 24380 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_261
timestamp 1676037725
transform 1 0 25116 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_273
timestamp 1676037725
transform 1 0 26220 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_285
timestamp 1676037725
transform 1 0 27324 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_297
timestamp 1676037725
transform 1 0 28428 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_92_305
timestamp 1676037725
transform 1 0 29164 0 1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_92_309
timestamp 1676037725
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_321
timestamp 1676037725
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_333
timestamp 1676037725
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_345
timestamp 1676037725
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1676037725
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1676037725
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_365
timestamp 1676037725
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_377
timestamp 1676037725
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_389
timestamp 1676037725
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_401
timestamp 1676037725
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1676037725
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1676037725
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1676037725
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_433
timestamp 1676037725
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_445
timestamp 1676037725
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_457
timestamp 1676037725
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_469
timestamp 1676037725
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1676037725
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_477
timestamp 1676037725
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_489
timestamp 1676037725
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_501
timestamp 1676037725
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_513
timestamp 1676037725
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_525
timestamp 1676037725
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_531
timestamp 1676037725
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_533
timestamp 1676037725
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_545
timestamp 1676037725
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_557
timestamp 1676037725
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_569
timestamp 1676037725
transform 1 0 53452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_581
timestamp 1676037725
transform 1 0 54556 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_587
timestamp 1676037725
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_589
timestamp 1676037725
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_601
timestamp 1676037725
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_613
timestamp 1676037725
transform 1 0 57500 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_3
timestamp 1676037725
transform 1 0 1380 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_9
timestamp 1676037725
transform 1 0 1932 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_21
timestamp 1676037725
transform 1 0 3036 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_33
timestamp 1676037725
transform 1 0 4140 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_45
timestamp 1676037725
transform 1 0 5244 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_93_53
timestamp 1676037725
transform 1 0 5980 0 -1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1676037725
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_69
timestamp 1676037725
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_81
timestamp 1676037725
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_93
timestamp 1676037725
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1676037725
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1676037725
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1676037725
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1676037725
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1676037725
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1676037725
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1676037725
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1676037725
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1676037725
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1676037725
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1676037725
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1676037725
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1676037725
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1676037725
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1676037725
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_237
timestamp 1676037725
transform 1 0 22908 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_243
timestamp 1676037725
transform 1 0 23460 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_251
timestamp 1676037725
transform 1 0 24196 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_93_261
timestamp 1676037725
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_273
timestamp 1676037725
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_279
timestamp 1676037725
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_281
timestamp 1676037725
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_293
timestamp 1676037725
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_305
timestamp 1676037725
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_317
timestamp 1676037725
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_329
timestamp 1676037725
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 1676037725
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_337
timestamp 1676037725
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_349
timestamp 1676037725
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_361
timestamp 1676037725
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_373
timestamp 1676037725
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1676037725
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1676037725
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_393
timestamp 1676037725
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_405
timestamp 1676037725
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_417
timestamp 1676037725
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_429
timestamp 1676037725
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_441
timestamp 1676037725
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1676037725
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_449
timestamp 1676037725
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_461
timestamp 1676037725
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_473
timestamp 1676037725
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_485
timestamp 1676037725
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_497
timestamp 1676037725
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1676037725
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_505
timestamp 1676037725
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_517
timestamp 1676037725
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_529
timestamp 1676037725
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_541
timestamp 1676037725
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_553
timestamp 1676037725
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_559
timestamp 1676037725
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_561
timestamp 1676037725
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_573
timestamp 1676037725
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_585
timestamp 1676037725
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_597
timestamp 1676037725
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_609
timestamp 1676037725
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_615
timestamp 1676037725
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_93_617
timestamp 1676037725
transform 1 0 57868 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_93_623
timestamp 1676037725
transform 1 0 58420 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_3
timestamp 1676037725
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_15
timestamp 1676037725
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1676037725
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1676037725
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1676037725
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1676037725
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_65
timestamp 1676037725
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1676037725
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1676037725
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1676037725
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_97
timestamp 1676037725
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_109
timestamp 1676037725
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1676037725
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1676037725
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1676037725
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1676037725
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1676037725
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1676037725
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1676037725
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1676037725
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1676037725
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1676037725
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1676037725
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_221
timestamp 1676037725
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_233
timestamp 1676037725
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_245
timestamp 1676037725
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 1676037725
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_253
timestamp 1676037725
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_265
timestamp 1676037725
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_277
timestamp 1676037725
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_289
timestamp 1676037725
transform 1 0 27692 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_301
timestamp 1676037725
transform 1 0 28796 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_307
timestamp 1676037725
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_309
timestamp 1676037725
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_321
timestamp 1676037725
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_333
timestamp 1676037725
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_345
timestamp 1676037725
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_357
timestamp 1676037725
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_363
timestamp 1676037725
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_365
timestamp 1676037725
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_377
timestamp 1676037725
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_389
timestamp 1676037725
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_401
timestamp 1676037725
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_413
timestamp 1676037725
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_419
timestamp 1676037725
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_421
timestamp 1676037725
transform 1 0 39836 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_425
timestamp 1676037725
transform 1 0 40204 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_434
timestamp 1676037725
transform 1 0 41032 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_438
timestamp 1676037725
transform 1 0 41400 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_450
timestamp 1676037725
transform 1 0 42504 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_462
timestamp 1676037725
transform 1 0 43608 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_94_474
timestamp 1676037725
transform 1 0 44712 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_477
timestamp 1676037725
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_489
timestamp 1676037725
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_501
timestamp 1676037725
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_513
timestamp 1676037725
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_525
timestamp 1676037725
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_531
timestamp 1676037725
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_533
timestamp 1676037725
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_545
timestamp 1676037725
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_557
timestamp 1676037725
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_569
timestamp 1676037725
transform 1 0 53452 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_581
timestamp 1676037725
transform 1 0 54556 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_587
timestamp 1676037725
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_589
timestamp 1676037725
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_601
timestamp 1676037725
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_613
timestamp 1676037725
transform 1 0 57500 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_3
timestamp 1676037725
transform 1 0 1380 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_95_9
timestamp 1676037725
transform 1 0 1932 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_21
timestamp 1676037725
transform 1 0 3036 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_33
timestamp 1676037725
transform 1 0 4140 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_45
timestamp 1676037725
transform 1 0 5244 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_95_53
timestamp 1676037725
transform 1 0 5980 0 -1 54400
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_95_57
timestamp 1676037725
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_69
timestamp 1676037725
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_81
timestamp 1676037725
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_93
timestamp 1676037725
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_105
timestamp 1676037725
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 1676037725
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_113
timestamp 1676037725
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_125
timestamp 1676037725
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_137
timestamp 1676037725
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_149
timestamp 1676037725
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_161
timestamp 1676037725
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 1676037725
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_169
timestamp 1676037725
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_181
timestamp 1676037725
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_193
timestamp 1676037725
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_205
timestamp 1676037725
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_217
timestamp 1676037725
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1676037725
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_225
timestamp 1676037725
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_237
timestamp 1676037725
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_249
timestamp 1676037725
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_261
timestamp 1676037725
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_273
timestamp 1676037725
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_279
timestamp 1676037725
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_281
timestamp 1676037725
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_293
timestamp 1676037725
transform 1 0 28060 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_305
timestamp 1676037725
transform 1 0 29164 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_317
timestamp 1676037725
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_329
timestamp 1676037725
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_335
timestamp 1676037725
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_337
timestamp 1676037725
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_349
timestamp 1676037725
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_361
timestamp 1676037725
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_373
timestamp 1676037725
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_385
timestamp 1676037725
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_391
timestamp 1676037725
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_393
timestamp 1676037725
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_405
timestamp 1676037725
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_417
timestamp 1676037725
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_429
timestamp 1676037725
transform 1 0 40572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_441
timestamp 1676037725
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_447
timestamp 1676037725
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_449
timestamp 1676037725
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_461
timestamp 1676037725
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_473
timestamp 1676037725
transform 1 0 44620 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_485
timestamp 1676037725
transform 1 0 45724 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_497
timestamp 1676037725
transform 1 0 46828 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_503
timestamp 1676037725
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_505
timestamp 1676037725
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_517
timestamp 1676037725
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_529
timestamp 1676037725
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_541
timestamp 1676037725
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_553
timestamp 1676037725
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_559
timestamp 1676037725
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_561
timestamp 1676037725
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_573
timestamp 1676037725
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_585
timestamp 1676037725
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_597
timestamp 1676037725
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_609
timestamp 1676037725
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_615
timestamp 1676037725
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_95_617
timestamp 1676037725
transform 1 0 57868 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_96_3
timestamp 1676037725
transform 1 0 1380 0 1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_96_9
timestamp 1676037725
transform 1 0 1932 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_21
timestamp 1676037725
transform 1 0 3036 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1676037725
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1676037725
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_41
timestamp 1676037725
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_53
timestamp 1676037725
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_65
timestamp 1676037725
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1676037725
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1676037725
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_85
timestamp 1676037725
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_97
timestamp 1676037725
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_109
timestamp 1676037725
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_121
timestamp 1676037725
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_133
timestamp 1676037725
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1676037725
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_141
timestamp 1676037725
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_153
timestamp 1676037725
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_165
timestamp 1676037725
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_177
timestamp 1676037725
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_189
timestamp 1676037725
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_195
timestamp 1676037725
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_197
timestamp 1676037725
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_209
timestamp 1676037725
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_221
timestamp 1676037725
transform 1 0 21436 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_96_233
timestamp 1676037725
transform 1 0 22540 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_96_250
timestamp 1676037725
transform 1 0 24104 0 1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_96_253
timestamp 1676037725
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_265
timestamp 1676037725
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_277
timestamp 1676037725
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_289
timestamp 1676037725
transform 1 0 27692 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_301
timestamp 1676037725
transform 1 0 28796 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_307
timestamp 1676037725
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_309
timestamp 1676037725
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_321
timestamp 1676037725
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_333
timestamp 1676037725
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_345
timestamp 1676037725
transform 1 0 32844 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_357
timestamp 1676037725
transform 1 0 33948 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_363
timestamp 1676037725
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_365
timestamp 1676037725
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_377
timestamp 1676037725
transform 1 0 35788 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_389
timestamp 1676037725
transform 1 0 36892 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_401
timestamp 1676037725
transform 1 0 37996 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_413
timestamp 1676037725
transform 1 0 39100 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_419
timestamp 1676037725
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_421
timestamp 1676037725
transform 1 0 39836 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_433
timestamp 1676037725
transform 1 0 40940 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_445
timestamp 1676037725
transform 1 0 42044 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_457
timestamp 1676037725
transform 1 0 43148 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_469
timestamp 1676037725
transform 1 0 44252 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_475
timestamp 1676037725
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_477
timestamp 1676037725
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_489
timestamp 1676037725
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_501
timestamp 1676037725
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_513
timestamp 1676037725
transform 1 0 48300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_525
timestamp 1676037725
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_531
timestamp 1676037725
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_533
timestamp 1676037725
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_545
timestamp 1676037725
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_557
timestamp 1676037725
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_569
timestamp 1676037725
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_581
timestamp 1676037725
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_587
timestamp 1676037725
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_589
timestamp 1676037725
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_601
timestamp 1676037725
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_613
timestamp 1676037725
transform 1 0 57500 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_619
timestamp 1676037725
transform 1 0 58052 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_96_623
timestamp 1676037725
transform 1 0 58420 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_3
timestamp 1676037725
transform 1 0 1380 0 -1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_97_9
timestamp 1676037725
transform 1 0 1932 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_21
timestamp 1676037725
transform 1 0 3036 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_33
timestamp 1676037725
transform 1 0 4140 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_45
timestamp 1676037725
transform 1 0 5244 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_97_53
timestamp 1676037725
transform 1 0 5980 0 -1 55488
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_97_57
timestamp 1676037725
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_69
timestamp 1676037725
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_81
timestamp 1676037725
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_93
timestamp 1676037725
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_105
timestamp 1676037725
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_111
timestamp 1676037725
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_113
timestamp 1676037725
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_125
timestamp 1676037725
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_137
timestamp 1676037725
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_149
timestamp 1676037725
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_161
timestamp 1676037725
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_167
timestamp 1676037725
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_169
timestamp 1676037725
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_181
timestamp 1676037725
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_193
timestamp 1676037725
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_205
timestamp 1676037725
transform 1 0 19964 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_217
timestamp 1676037725
transform 1 0 21068 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_223
timestamp 1676037725
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_225
timestamp 1676037725
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_237
timestamp 1676037725
transform 1 0 22908 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_249
timestamp 1676037725
transform 1 0 24012 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_261
timestamp 1676037725
transform 1 0 25116 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_273
timestamp 1676037725
transform 1 0 26220 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_279
timestamp 1676037725
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_281
timestamp 1676037725
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_293
timestamp 1676037725
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_305
timestamp 1676037725
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_317
timestamp 1676037725
transform 1 0 30268 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_329
timestamp 1676037725
transform 1 0 31372 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_335
timestamp 1676037725
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_337
timestamp 1676037725
transform 1 0 32108 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_349
timestamp 1676037725
transform 1 0 33212 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_361
timestamp 1676037725
transform 1 0 34316 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_373
timestamp 1676037725
transform 1 0 35420 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_385
timestamp 1676037725
transform 1 0 36524 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_391
timestamp 1676037725
transform 1 0 37076 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_393
timestamp 1676037725
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_405
timestamp 1676037725
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_417
timestamp 1676037725
transform 1 0 39468 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_97_429
timestamp 1676037725
transform 1 0 40572 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_97_440
timestamp 1676037725
transform 1 0 41584 0 -1 55488
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_97_449
timestamp 1676037725
transform 1 0 42412 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_461
timestamp 1676037725
transform 1 0 43516 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_473
timestamp 1676037725
transform 1 0 44620 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_485
timestamp 1676037725
transform 1 0 45724 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_497
timestamp 1676037725
transform 1 0 46828 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_503
timestamp 1676037725
transform 1 0 47380 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_505
timestamp 1676037725
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_517
timestamp 1676037725
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_529
timestamp 1676037725
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_541
timestamp 1676037725
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_553
timestamp 1676037725
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_559
timestamp 1676037725
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_561
timestamp 1676037725
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_573
timestamp 1676037725
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_585
timestamp 1676037725
transform 1 0 54924 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_597
timestamp 1676037725
transform 1 0 56028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_609
timestamp 1676037725
transform 1 0 57132 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_615
timestamp 1676037725
transform 1 0 57684 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_97_617
timestamp 1676037725
transform 1 0 57868 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_98_3
timestamp 1676037725
transform 1 0 1380 0 1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_98_9
timestamp 1676037725
transform 1 0 1932 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_21
timestamp 1676037725
transform 1 0 3036 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1676037725
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1676037725
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_41
timestamp 1676037725
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_53
timestamp 1676037725
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_65
timestamp 1676037725
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1676037725
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1676037725
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_85
timestamp 1676037725
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_97
timestamp 1676037725
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_109
timestamp 1676037725
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_121
timestamp 1676037725
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_133
timestamp 1676037725
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_139
timestamp 1676037725
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_141
timestamp 1676037725
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_153
timestamp 1676037725
transform 1 0 15180 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_165
timestamp 1676037725
transform 1 0 16284 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_177
timestamp 1676037725
transform 1 0 17388 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_189
timestamp 1676037725
transform 1 0 18492 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_195
timestamp 1676037725
transform 1 0 19044 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_197
timestamp 1676037725
transform 1 0 19228 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_209
timestamp 1676037725
transform 1 0 20332 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_221
timestamp 1676037725
transform 1 0 21436 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_233
timestamp 1676037725
transform 1 0 22540 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_245
timestamp 1676037725
transform 1 0 23644 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_251
timestamp 1676037725
transform 1 0 24196 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_98_253
timestamp 1676037725
transform 1 0 24380 0 1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_98_269
timestamp 1676037725
transform 1 0 25852 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_281
timestamp 1676037725
transform 1 0 26956 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_293
timestamp 1676037725
transform 1 0 28060 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_98_305
timestamp 1676037725
transform 1 0 29164 0 1 55488
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_98_309
timestamp 1676037725
transform 1 0 29532 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_321
timestamp 1676037725
transform 1 0 30636 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_333
timestamp 1676037725
transform 1 0 31740 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_345
timestamp 1676037725
transform 1 0 32844 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_357
timestamp 1676037725
transform 1 0 33948 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_363
timestamp 1676037725
transform 1 0 34500 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_365
timestamp 1676037725
transform 1 0 34684 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_377
timestamp 1676037725
transform 1 0 35788 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_389
timestamp 1676037725
transform 1 0 36892 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_401
timestamp 1676037725
transform 1 0 37996 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_413
timestamp 1676037725
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_419
timestamp 1676037725
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_421
timestamp 1676037725
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_433
timestamp 1676037725
transform 1 0 40940 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_445
timestamp 1676037725
transform 1 0 42044 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_457
timestamp 1676037725
transform 1 0 43148 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_469
timestamp 1676037725
transform 1 0 44252 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_475
timestamp 1676037725
transform 1 0 44804 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_477
timestamp 1676037725
transform 1 0 44988 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_489
timestamp 1676037725
transform 1 0 46092 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_501
timestamp 1676037725
transform 1 0 47196 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_513
timestamp 1676037725
transform 1 0 48300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_525
timestamp 1676037725
transform 1 0 49404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_531
timestamp 1676037725
transform 1 0 49956 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_533
timestamp 1676037725
transform 1 0 50140 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_545
timestamp 1676037725
transform 1 0 51244 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_557
timestamp 1676037725
transform 1 0 52348 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_569
timestamp 1676037725
transform 1 0 53452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_581
timestamp 1676037725
transform 1 0 54556 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_587
timestamp 1676037725
transform 1 0 55108 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_589
timestamp 1676037725
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_601
timestamp 1676037725
transform 1 0 56396 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_613
timestamp 1676037725
transform 1 0 57500 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_619
timestamp 1676037725
transform 1 0 58052 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_98_623
timestamp 1676037725
transform 1 0 58420 0 1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_99_3
timestamp 1676037725
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_15
timestamp 1676037725
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_27
timestamp 1676037725
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_39
timestamp 1676037725
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_51
timestamp 1676037725
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1676037725
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_57
timestamp 1676037725
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_69
timestamp 1676037725
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_81
timestamp 1676037725
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_93
timestamp 1676037725
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_105
timestamp 1676037725
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 1676037725
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_113
timestamp 1676037725
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_125
timestamp 1676037725
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_137
timestamp 1676037725
transform 1 0 13708 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_149
timestamp 1676037725
transform 1 0 14812 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_161
timestamp 1676037725
transform 1 0 15916 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_167
timestamp 1676037725
transform 1 0 16468 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_169
timestamp 1676037725
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_181
timestamp 1676037725
transform 1 0 17756 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_193
timestamp 1676037725
transform 1 0 18860 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_205
timestamp 1676037725
transform 1 0 19964 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_217
timestamp 1676037725
transform 1 0 21068 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_223
timestamp 1676037725
transform 1 0 21620 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_225
timestamp 1676037725
transform 1 0 21804 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_237
timestamp 1676037725
transform 1 0 22908 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_99_245
timestamp 1676037725
transform 1 0 23644 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_260
timestamp 1676037725
transform 1 0 25024 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_272
timestamp 1676037725
transform 1 0 26128 0 -1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_99_281
timestamp 1676037725
transform 1 0 26956 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_293
timestamp 1676037725
transform 1 0 28060 0 -1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_99_315
timestamp 1676037725
transform 1 0 30084 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_327
timestamp 1676037725
transform 1 0 31188 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_99_335
timestamp 1676037725
transform 1 0 31924 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_337
timestamp 1676037725
transform 1 0 32108 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_349
timestamp 1676037725
transform 1 0 33212 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_361
timestamp 1676037725
transform 1 0 34316 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_373
timestamp 1676037725
transform 1 0 35420 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_385
timestamp 1676037725
transform 1 0 36524 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_391
timestamp 1676037725
transform 1 0 37076 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_393
timestamp 1676037725
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_405
timestamp 1676037725
transform 1 0 38364 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_417
timestamp 1676037725
transform 1 0 39468 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_99_429
timestamp 1676037725
transform 1 0 40572 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_99_446
timestamp 1676037725
transform 1 0 42136 0 -1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_99_449
timestamp 1676037725
transform 1 0 42412 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_461
timestamp 1676037725
transform 1 0 43516 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_473
timestamp 1676037725
transform 1 0 44620 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_485
timestamp 1676037725
transform 1 0 45724 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_497
timestamp 1676037725
transform 1 0 46828 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_503
timestamp 1676037725
transform 1 0 47380 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_505
timestamp 1676037725
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_517
timestamp 1676037725
transform 1 0 48668 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_529
timestamp 1676037725
transform 1 0 49772 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_541
timestamp 1676037725
transform 1 0 50876 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_553
timestamp 1676037725
transform 1 0 51980 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_559
timestamp 1676037725
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_561
timestamp 1676037725
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_573
timestamp 1676037725
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_585
timestamp 1676037725
transform 1 0 54924 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_597
timestamp 1676037725
transform 1 0 56028 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_609
timestamp 1676037725
transform 1 0 57132 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_615
timestamp 1676037725
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_99_617
timestamp 1676037725
transform 1 0 57868 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_623
timestamp 1676037725
transform 1 0 58420 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_100_3
timestamp 1676037725
transform 1 0 1380 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_11
timestamp 1676037725
transform 1 0 2116 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_23
timestamp 1676037725
transform 1 0 3220 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1676037725
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_29
timestamp 1676037725
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_41
timestamp 1676037725
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_53
timestamp 1676037725
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_65
timestamp 1676037725
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_77
timestamp 1676037725
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1676037725
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_85
timestamp 1676037725
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_97
timestamp 1676037725
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_109
timestamp 1676037725
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_121
timestamp 1676037725
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_133
timestamp 1676037725
transform 1 0 13340 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_139
timestamp 1676037725
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_141
timestamp 1676037725
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_153
timestamp 1676037725
transform 1 0 15180 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_165
timestamp 1676037725
transform 1 0 16284 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_177
timestamp 1676037725
transform 1 0 17388 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_189
timestamp 1676037725
transform 1 0 18492 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_195
timestamp 1676037725
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_197
timestamp 1676037725
transform 1 0 19228 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_209
timestamp 1676037725
transform 1 0 20332 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_221
timestamp 1676037725
transform 1 0 21436 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_233
timestamp 1676037725
transform 1 0 22540 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_245
timestamp 1676037725
transform 1 0 23644 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_251
timestamp 1676037725
transform 1 0 24196 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_253
timestamp 1676037725
transform 1 0 24380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_265
timestamp 1676037725
transform 1 0 25484 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_277
timestamp 1676037725
transform 1 0 26588 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_289
timestamp 1676037725
transform 1 0 27692 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_301
timestamp 1676037725
transform 1 0 28796 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_307
timestamp 1676037725
transform 1 0 29348 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_309
timestamp 1676037725
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_321
timestamp 1676037725
transform 1 0 30636 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_333
timestamp 1676037725
transform 1 0 31740 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_339
timestamp 1676037725
transform 1 0 32292 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_100_354
timestamp 1676037725
transform 1 0 33672 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_362
timestamp 1676037725
transform 1 0 34408 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_365
timestamp 1676037725
transform 1 0 34684 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_377
timestamp 1676037725
transform 1 0 35788 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_389
timestamp 1676037725
transform 1 0 36892 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_401
timestamp 1676037725
transform 1 0 37996 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_413
timestamp 1676037725
transform 1 0 39100 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_419
timestamp 1676037725
transform 1 0 39652 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_421
timestamp 1676037725
transform 1 0 39836 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_433
timestamp 1676037725
transform 1 0 40940 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_445
timestamp 1676037725
transform 1 0 42044 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_457
timestamp 1676037725
transform 1 0 43148 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_469
timestamp 1676037725
transform 1 0 44252 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_475
timestamp 1676037725
transform 1 0 44804 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_477
timestamp 1676037725
transform 1 0 44988 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_489
timestamp 1676037725
transform 1 0 46092 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_501
timestamp 1676037725
transform 1 0 47196 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_513
timestamp 1676037725
transform 1 0 48300 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_525
timestamp 1676037725
transform 1 0 49404 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_531
timestamp 1676037725
transform 1 0 49956 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_533
timestamp 1676037725
transform 1 0 50140 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_545
timestamp 1676037725
transform 1 0 51244 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_557
timestamp 1676037725
transform 1 0 52348 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_569
timestamp 1676037725
transform 1 0 53452 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_581
timestamp 1676037725
transform 1 0 54556 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_587
timestamp 1676037725
transform 1 0 55108 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_589
timestamp 1676037725
transform 1 0 55292 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_601
timestamp 1676037725
transform 1 0 56396 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_613
timestamp 1676037725
transform 1 0 57500 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_623
timestamp 1676037725
transform 1 0 58420 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_3
timestamp 1676037725
transform 1 0 1380 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_9
timestamp 1676037725
transform 1 0 1932 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_21
timestamp 1676037725
transform 1 0 3036 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_33
timestamp 1676037725
transform 1 0 4140 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_45
timestamp 1676037725
transform 1 0 5244 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_53
timestamp 1676037725
transform 1 0 5980 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_57
timestamp 1676037725
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_69
timestamp 1676037725
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_81
timestamp 1676037725
transform 1 0 8556 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_93
timestamp 1676037725
transform 1 0 9660 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_105
timestamp 1676037725
transform 1 0 10764 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_111
timestamp 1676037725
transform 1 0 11316 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_113
timestamp 1676037725
transform 1 0 11500 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_125
timestamp 1676037725
transform 1 0 12604 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_137
timestamp 1676037725
transform 1 0 13708 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_149
timestamp 1676037725
transform 1 0 14812 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_161
timestamp 1676037725
transform 1 0 15916 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_167
timestamp 1676037725
transform 1 0 16468 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_169
timestamp 1676037725
transform 1 0 16652 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_181
timestamp 1676037725
transform 1 0 17756 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_193
timestamp 1676037725
transform 1 0 18860 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_205
timestamp 1676037725
transform 1 0 19964 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_217
timestamp 1676037725
transform 1 0 21068 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_223
timestamp 1676037725
transform 1 0 21620 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_225
timestamp 1676037725
transform 1 0 21804 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_237
timestamp 1676037725
transform 1 0 22908 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_249
timestamp 1676037725
transform 1 0 24012 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_261
timestamp 1676037725
transform 1 0 25116 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_273
timestamp 1676037725
transform 1 0 26220 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_279
timestamp 1676037725
transform 1 0 26772 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_281
timestamp 1676037725
transform 1 0 26956 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_293
timestamp 1676037725
transform 1 0 28060 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_305
timestamp 1676037725
transform 1 0 29164 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_317
timestamp 1676037725
transform 1 0 30268 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_329
timestamp 1676037725
transform 1 0 31372 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_335
timestamp 1676037725
transform 1 0 31924 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_337
timestamp 1676037725
transform 1 0 32108 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_349
timestamp 1676037725
transform 1 0 33212 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_361
timestamp 1676037725
transform 1 0 34316 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_373
timestamp 1676037725
transform 1 0 35420 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_384
timestamp 1676037725
transform 1 0 36432 0 -1 57664
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_101_393
timestamp 1676037725
transform 1 0 37260 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_405
timestamp 1676037725
transform 1 0 38364 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_417
timestamp 1676037725
transform 1 0 39468 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_429
timestamp 1676037725
transform 1 0 40572 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_441
timestamp 1676037725
transform 1 0 41676 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_447
timestamp 1676037725
transform 1 0 42228 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_449
timestamp 1676037725
transform 1 0 42412 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_461
timestamp 1676037725
transform 1 0 43516 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_473
timestamp 1676037725
transform 1 0 44620 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_485
timestamp 1676037725
transform 1 0 45724 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_497
timestamp 1676037725
transform 1 0 46828 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_503
timestamp 1676037725
transform 1 0 47380 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_505
timestamp 1676037725
transform 1 0 47564 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_517
timestamp 1676037725
transform 1 0 48668 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_529
timestamp 1676037725
transform 1 0 49772 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_541
timestamp 1676037725
transform 1 0 50876 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_553
timestamp 1676037725
transform 1 0 51980 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_559
timestamp 1676037725
transform 1 0 52532 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_561
timestamp 1676037725
transform 1 0 52716 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_573
timestamp 1676037725
transform 1 0 53820 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_585
timestamp 1676037725
transform 1 0 54924 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_597
timestamp 1676037725
transform 1 0 56028 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_609
timestamp 1676037725
transform 1 0 57132 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_615
timestamp 1676037725
transform 1 0 57684 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_617
timestamp 1676037725
transform 1 0 57868 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_102_3
timestamp 1676037725
transform 1 0 1380 0 1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_102_11
timestamp 1676037725
transform 1 0 2116 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_102_23
timestamp 1676037725
transform 1 0 3220 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_102_27
timestamp 1676037725
transform 1 0 3588 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_29
timestamp 1676037725
transform 1 0 3772 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_41
timestamp 1676037725
transform 1 0 4876 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_53
timestamp 1676037725
transform 1 0 5980 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_65
timestamp 1676037725
transform 1 0 7084 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_77
timestamp 1676037725
transform 1 0 8188 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_83
timestamp 1676037725
transform 1 0 8740 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_85
timestamp 1676037725
transform 1 0 8924 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_97
timestamp 1676037725
transform 1 0 10028 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_109
timestamp 1676037725
transform 1 0 11132 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_121
timestamp 1676037725
transform 1 0 12236 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_133
timestamp 1676037725
transform 1 0 13340 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_139
timestamp 1676037725
transform 1 0 13892 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_141
timestamp 1676037725
transform 1 0 14076 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_153
timestamp 1676037725
transform 1 0 15180 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_165
timestamp 1676037725
transform 1 0 16284 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_177
timestamp 1676037725
transform 1 0 17388 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_189
timestamp 1676037725
transform 1 0 18492 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_195
timestamp 1676037725
transform 1 0 19044 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_197
timestamp 1676037725
transform 1 0 19228 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_209
timestamp 1676037725
transform 1 0 20332 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_221
timestamp 1676037725
transform 1 0 21436 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_233
timestamp 1676037725
transform 1 0 22540 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_245
timestamp 1676037725
transform 1 0 23644 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_251
timestamp 1676037725
transform 1 0 24196 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_253
timestamp 1676037725
transform 1 0 24380 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_265
timestamp 1676037725
transform 1 0 25484 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_277
timestamp 1676037725
transform 1 0 26588 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_289
timestamp 1676037725
transform 1 0 27692 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_301
timestamp 1676037725
transform 1 0 28796 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_307
timestamp 1676037725
transform 1 0 29348 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_309
timestamp 1676037725
transform 1 0 29532 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_321
timestamp 1676037725
transform 1 0 30636 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_333
timestamp 1676037725
transform 1 0 31740 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_345
timestamp 1676037725
transform 1 0 32844 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_357
timestamp 1676037725
transform 1 0 33948 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_363
timestamp 1676037725
transform 1 0 34500 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_102_365
timestamp 1676037725
transform 1 0 34684 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_102_369
timestamp 1676037725
transform 1 0 35052 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_387
timestamp 1676037725
transform 1 0 36708 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_399
timestamp 1676037725
transform 1 0 37812 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_102_411
timestamp 1676037725
transform 1 0 38916 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_102_419
timestamp 1676037725
transform 1 0 39652 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_421
timestamp 1676037725
transform 1 0 39836 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_433
timestamp 1676037725
transform 1 0 40940 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_445
timestamp 1676037725
transform 1 0 42044 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_457
timestamp 1676037725
transform 1 0 43148 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_469
timestamp 1676037725
transform 1 0 44252 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_475
timestamp 1676037725
transform 1 0 44804 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_477
timestamp 1676037725
transform 1 0 44988 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_489
timestamp 1676037725
transform 1 0 46092 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_501
timestamp 1676037725
transform 1 0 47196 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_513
timestamp 1676037725
transform 1 0 48300 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_525
timestamp 1676037725
transform 1 0 49404 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_531
timestamp 1676037725
transform 1 0 49956 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_533
timestamp 1676037725
transform 1 0 50140 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_545
timestamp 1676037725
transform 1 0 51244 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_557
timestamp 1676037725
transform 1 0 52348 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_569
timestamp 1676037725
transform 1 0 53452 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_581
timestamp 1676037725
transform 1 0 54556 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_587
timestamp 1676037725
transform 1 0 55108 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_589
timestamp 1676037725
transform 1 0 55292 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_601
timestamp 1676037725
transform 1 0 56396 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_102_613
timestamp 1676037725
transform 1 0 57500 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_102_623
timestamp 1676037725
transform 1 0 58420 0 1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_103_3
timestamp 1676037725
transform 1 0 1380 0 -1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_103_11
timestamp 1676037725
transform 1 0 2116 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_23
timestamp 1676037725
transform 1 0 3220 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_35
timestamp 1676037725
transform 1 0 4324 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_103_47
timestamp 1676037725
transform 1 0 5428 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_103_55
timestamp 1676037725
transform 1 0 6164 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_57
timestamp 1676037725
transform 1 0 6348 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_69
timestamp 1676037725
transform 1 0 7452 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_81
timestamp 1676037725
transform 1 0 8556 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_93
timestamp 1676037725
transform 1 0 9660 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_105
timestamp 1676037725
transform 1 0 10764 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_111
timestamp 1676037725
transform 1 0 11316 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_113
timestamp 1676037725
transform 1 0 11500 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_125
timestamp 1676037725
transform 1 0 12604 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_137
timestamp 1676037725
transform 1 0 13708 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_149
timestamp 1676037725
transform 1 0 14812 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_161
timestamp 1676037725
transform 1 0 15916 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_167
timestamp 1676037725
transform 1 0 16468 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_169
timestamp 1676037725
transform 1 0 16652 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_181
timestamp 1676037725
transform 1 0 17756 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_193
timestamp 1676037725
transform 1 0 18860 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_205
timestamp 1676037725
transform 1 0 19964 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_217
timestamp 1676037725
transform 1 0 21068 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_223
timestamp 1676037725
transform 1 0 21620 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_225
timestamp 1676037725
transform 1 0 21804 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_237
timestamp 1676037725
transform 1 0 22908 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_249
timestamp 1676037725
transform 1 0 24012 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_261
timestamp 1676037725
transform 1 0 25116 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_273
timestamp 1676037725
transform 1 0 26220 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_279
timestamp 1676037725
transform 1 0 26772 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_281
timestamp 1676037725
transform 1 0 26956 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_293
timestamp 1676037725
transform 1 0 28060 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_305
timestamp 1676037725
transform 1 0 29164 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_317
timestamp 1676037725
transform 1 0 30268 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_329
timestamp 1676037725
transform 1 0 31372 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_335
timestamp 1676037725
transform 1 0 31924 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_337
timestamp 1676037725
transform 1 0 32108 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_349
timestamp 1676037725
transform 1 0 33212 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_361
timestamp 1676037725
transform 1 0 34316 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_373
timestamp 1676037725
transform 1 0 35420 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_385
timestamp 1676037725
transform 1 0 36524 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_391
timestamp 1676037725
transform 1 0 37076 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_103_393
timestamp 1676037725
transform 1 0 37260 0 -1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_103_412
timestamp 1676037725
transform 1 0 39008 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_103_424
timestamp 1676037725
transform 1 0 40112 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_103_446
timestamp 1676037725
transform 1 0 42136 0 -1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_103_449
timestamp 1676037725
transform 1 0 42412 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_461
timestamp 1676037725
transform 1 0 43516 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_473
timestamp 1676037725
transform 1 0 44620 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_485
timestamp 1676037725
transform 1 0 45724 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_497
timestamp 1676037725
transform 1 0 46828 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_503
timestamp 1676037725
transform 1 0 47380 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_505
timestamp 1676037725
transform 1 0 47564 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_517
timestamp 1676037725
transform 1 0 48668 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_529
timestamp 1676037725
transform 1 0 49772 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_541
timestamp 1676037725
transform 1 0 50876 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_553
timestamp 1676037725
transform 1 0 51980 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_559
timestamp 1676037725
transform 1 0 52532 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_561
timestamp 1676037725
transform 1 0 52716 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_573
timestamp 1676037725
transform 1 0 53820 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_585
timestamp 1676037725
transform 1 0 54924 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_597
timestamp 1676037725
transform 1 0 56028 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_609
timestamp 1676037725
transform 1 0 57132 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_615
timestamp 1676037725
transform 1 0 57684 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_103_617
timestamp 1676037725
transform 1 0 57868 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_103_623
timestamp 1676037725
transform 1 0 58420 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_104_3
timestamp 1676037725
transform 1 0 1380 0 1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_104_9
timestamp 1676037725
transform 1 0 1932 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_21
timestamp 1676037725
transform 1 0 3036 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_27
timestamp 1676037725
transform 1 0 3588 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_29
timestamp 1676037725
transform 1 0 3772 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_41
timestamp 1676037725
transform 1 0 4876 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_53
timestamp 1676037725
transform 1 0 5980 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_65
timestamp 1676037725
transform 1 0 7084 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_77
timestamp 1676037725
transform 1 0 8188 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_83
timestamp 1676037725
transform 1 0 8740 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_85
timestamp 1676037725
transform 1 0 8924 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_97
timestamp 1676037725
transform 1 0 10028 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_109
timestamp 1676037725
transform 1 0 11132 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_121
timestamp 1676037725
transform 1 0 12236 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_133
timestamp 1676037725
transform 1 0 13340 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_139
timestamp 1676037725
transform 1 0 13892 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_141
timestamp 1676037725
transform 1 0 14076 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_153
timestamp 1676037725
transform 1 0 15180 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_165
timestamp 1676037725
transform 1 0 16284 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_177
timestamp 1676037725
transform 1 0 17388 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_189
timestamp 1676037725
transform 1 0 18492 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_195
timestamp 1676037725
transform 1 0 19044 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_104_197
timestamp 1676037725
transform 1 0 19228 0 1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_104_207
timestamp 1676037725
transform 1 0 20148 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_219
timestamp 1676037725
transform 1 0 21252 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_231
timestamp 1676037725
transform 1 0 22356 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_243
timestamp 1676037725
transform 1 0 23460 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_104_251
timestamp 1676037725
transform 1 0 24196 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_253
timestamp 1676037725
transform 1 0 24380 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_265
timestamp 1676037725
transform 1 0 25484 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_277
timestamp 1676037725
transform 1 0 26588 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_289
timestamp 1676037725
transform 1 0 27692 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_301
timestamp 1676037725
transform 1 0 28796 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_307
timestamp 1676037725
transform 1 0 29348 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_309
timestamp 1676037725
transform 1 0 29532 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_321
timestamp 1676037725
transform 1 0 30636 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_333
timestamp 1676037725
transform 1 0 31740 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_345
timestamp 1676037725
transform 1 0 32844 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_357
timestamp 1676037725
transform 1 0 33948 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_363
timestamp 1676037725
transform 1 0 34500 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_365
timestamp 1676037725
transform 1 0 34684 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_377
timestamp 1676037725
transform 1 0 35788 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_389
timestamp 1676037725
transform 1 0 36892 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_401
timestamp 1676037725
transform 1 0 37996 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_413
timestamp 1676037725
transform 1 0 39100 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_419
timestamp 1676037725
transform 1 0 39652 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_104_421
timestamp 1676037725
transform 1 0 39836 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_104_429
timestamp 1676037725
transform 1 0 40572 0 1 58752
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_104_446
timestamp 1676037725
transform 1 0 42136 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_458
timestamp 1676037725
transform 1 0 43240 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_470
timestamp 1676037725
transform 1 0 44344 0 1 58752
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_104_477
timestamp 1676037725
transform 1 0 44988 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_489
timestamp 1676037725
transform 1 0 46092 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_501
timestamp 1676037725
transform 1 0 47196 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_513
timestamp 1676037725
transform 1 0 48300 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_525
timestamp 1676037725
transform 1 0 49404 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_531
timestamp 1676037725
transform 1 0 49956 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_533
timestamp 1676037725
transform 1 0 50140 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_545
timestamp 1676037725
transform 1 0 51244 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_557
timestamp 1676037725
transform 1 0 52348 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_569
timestamp 1676037725
transform 1 0 53452 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_581
timestamp 1676037725
transform 1 0 54556 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_587
timestamp 1676037725
transform 1 0 55108 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_589
timestamp 1676037725
transform 1 0 55292 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_601
timestamp 1676037725
transform 1 0 56396 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_104_613
timestamp 1676037725
transform 1 0 57500 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_104_623
timestamp 1676037725
transform 1 0 58420 0 1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_105_3
timestamp 1676037725
transform 1 0 1380 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_105_11
timestamp 1676037725
transform 1 0 2116 0 -1 59840
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_105_19
timestamp 1676037725
transform 1 0 2852 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_31
timestamp 1676037725
transform 1 0 3956 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_43
timestamp 1676037725
transform 1 0 5060 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_105_55
timestamp 1676037725
transform 1 0 6164 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_57
timestamp 1676037725
transform 1 0 6348 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_69
timestamp 1676037725
transform 1 0 7452 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_81
timestamp 1676037725
transform 1 0 8556 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_93
timestamp 1676037725
transform 1 0 9660 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_105
timestamp 1676037725
transform 1 0 10764 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_111
timestamp 1676037725
transform 1 0 11316 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_113
timestamp 1676037725
transform 1 0 11500 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_125
timestamp 1676037725
transform 1 0 12604 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_137
timestamp 1676037725
transform 1 0 13708 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_149
timestamp 1676037725
transform 1 0 14812 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_161
timestamp 1676037725
transform 1 0 15916 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_167
timestamp 1676037725
transform 1 0 16468 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_169
timestamp 1676037725
transform 1 0 16652 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_181
timestamp 1676037725
transform 1 0 17756 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_105_193
timestamp 1676037725
transform 1 0 18860 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_105_197
timestamp 1676037725
transform 1 0 19228 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_105_206
timestamp 1676037725
transform 1 0 20056 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_105_221
timestamp 1676037725
transform 1 0 21436 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_105_225
timestamp 1676037725
transform 1 0 21804 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_105_236
timestamp 1676037725
transform 1 0 22816 0 -1 59840
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_105_248
timestamp 1676037725
transform 1 0 23920 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_260
timestamp 1676037725
transform 1 0 25024 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_272
timestamp 1676037725
transform 1 0 26128 0 -1 59840
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_105_281
timestamp 1676037725
transform 1 0 26956 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_105_293
timestamp 1676037725
transform 1 0 28060 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_105_302
timestamp 1676037725
transform 1 0 28888 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_105_306
timestamp 1676037725
transform 1 0 29256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_105_309
timestamp 1676037725
transform 1 0 29532 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_105_319
timestamp 1676037725
transform 1 0 30452 0 -1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_105_323
timestamp 1676037725
transform 1 0 30820 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_105_335
timestamp 1676037725
transform 1 0 31924 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_337
timestamp 1676037725
transform 1 0 32108 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_349
timestamp 1676037725
transform 1 0 33212 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_361
timestamp 1676037725
transform 1 0 34316 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_373
timestamp 1676037725
transform 1 0 35420 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_385
timestamp 1676037725
transform 1 0 36524 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_391
timestamp 1676037725
transform 1 0 37076 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_393
timestamp 1676037725
transform 1 0 37260 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_405
timestamp 1676037725
transform 1 0 38364 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_417
timestamp 1676037725
transform 1 0 39468 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_429
timestamp 1676037725
transform 1 0 40572 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_441
timestamp 1676037725
transform 1 0 41676 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_447
timestamp 1676037725
transform 1 0 42228 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_105_449
timestamp 1676037725
transform 1 0 42412 0 -1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_105_465
timestamp 1676037725
transform 1 0 43884 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_477
timestamp 1676037725
transform 1 0 44988 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_489
timestamp 1676037725
transform 1 0 46092 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_105_501
timestamp 1676037725
transform 1 0 47196 0 -1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_105_505
timestamp 1676037725
transform 1 0 47564 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_517
timestamp 1676037725
transform 1 0 48668 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_529
timestamp 1676037725
transform 1 0 49772 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_541
timestamp 1676037725
transform 1 0 50876 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_553
timestamp 1676037725
transform 1 0 51980 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_559
timestamp 1676037725
transform 1 0 52532 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_561
timestamp 1676037725
transform 1 0 52716 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_573
timestamp 1676037725
transform 1 0 53820 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_585
timestamp 1676037725
transform 1 0 54924 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_597
timestamp 1676037725
transform 1 0 56028 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_105_609
timestamp 1676037725
transform 1 0 57132 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_105_614
timestamp 1676037725
transform 1 0 57592 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_105_617
timestamp 1676037725
transform 1 0 57868 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_105_623
timestamp 1676037725
transform 1 0 58420 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_106_3
timestamp 1676037725
transform 1 0 1380 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_106_11
timestamp 1676037725
transform 1 0 2116 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_106_19
timestamp 1676037725
transform 1 0 2852 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_106_27
timestamp 1676037725
transform 1 0 3588 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_29
timestamp 1676037725
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_41
timestamp 1676037725
transform 1 0 4876 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_53
timestamp 1676037725
transform 1 0 5980 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_65
timestamp 1676037725
transform 1 0 7084 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_106_75
timestamp 1676037725
transform 1 0 8004 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_106_83
timestamp 1676037725
transform 1 0 8740 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_85
timestamp 1676037725
transform 1 0 8924 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_97
timestamp 1676037725
transform 1 0 10028 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_109
timestamp 1676037725
transform 1 0 11132 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_121
timestamp 1676037725
transform 1 0 12236 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_133
timestamp 1676037725
transform 1 0 13340 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_139
timestamp 1676037725
transform 1 0 13892 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_141
timestamp 1676037725
transform 1 0 14076 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_153
timestamp 1676037725
transform 1 0 15180 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_165
timestamp 1676037725
transform 1 0 16284 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_106_191
timestamp 1676037725
transform 1 0 18676 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_106_195
timestamp 1676037725
transform 1 0 19044 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_197
timestamp 1676037725
transform 1 0 19228 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_209
timestamp 1676037725
transform 1 0 20332 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_106_218
timestamp 1676037725
transform 1 0 21160 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_106_239
timestamp 1676037725
transform 1 0 23092 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_106_250
timestamp 1676037725
transform 1 0 24104 0 1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_106_253
timestamp 1676037725
transform 1 0 24380 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_265
timestamp 1676037725
transform 1 0 25484 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_277
timestamp 1676037725
transform 1 0 26588 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_106_289
timestamp 1676037725
transform 1 0 27692 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_106_302
timestamp 1676037725
transform 1 0 28888 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_106_309
timestamp 1676037725
transform 1 0 29532 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_106_313
timestamp 1676037725
transform 1 0 29900 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_106_316
timestamp 1676037725
transform 1 0 30176 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_106_327
timestamp 1676037725
transform 1 0 31188 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_106_335
timestamp 1676037725
transform 1 0 31924 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_350
timestamp 1676037725
transform 1 0 33304 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_106_362
timestamp 1676037725
transform 1 0 34408 0 1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_106_365
timestamp 1676037725
transform 1 0 34684 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_377
timestamp 1676037725
transform 1 0 35788 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_389
timestamp 1676037725
transform 1 0 36892 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_401
timestamp 1676037725
transform 1 0 37996 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_413
timestamp 1676037725
transform 1 0 39100 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_419
timestamp 1676037725
transform 1 0 39652 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_106_421
timestamp 1676037725
transform 1 0 39836 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_106_437
timestamp 1676037725
transform 1 0 41308 0 1 59840
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_106_455
timestamp 1676037725
transform 1 0 42964 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_467
timestamp 1676037725
transform 1 0 44068 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_106_475
timestamp 1676037725
transform 1 0 44804 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_477
timestamp 1676037725
transform 1 0 44988 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_489
timestamp 1676037725
transform 1 0 46092 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_501
timestamp 1676037725
transform 1 0 47196 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_513
timestamp 1676037725
transform 1 0 48300 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_525
timestamp 1676037725
transform 1 0 49404 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_531
timestamp 1676037725
transform 1 0 49956 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_533
timestamp 1676037725
transform 1 0 50140 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_545
timestamp 1676037725
transform 1 0 51244 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_557
timestamp 1676037725
transform 1 0 52348 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_569
timestamp 1676037725
transform 1 0 53452 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_581
timestamp 1676037725
transform 1 0 54556 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_587
timestamp 1676037725
transform 1 0 55108 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_589
timestamp 1676037725
transform 1 0 55292 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_106_605
timestamp 1676037725
transform 1 0 56764 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_106_613
timestamp 1676037725
transform 1 0 57500 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_106_623
timestamp 1676037725
transform 1 0 58420 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_107_3
timestamp 1676037725
transform 1 0 1380 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_107_11
timestamp 1676037725
transform 1 0 2116 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_107_19
timestamp 1676037725
transform 1 0 2852 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_107_26
timestamp 1676037725
transform 1 0 3496 0 -1 60928
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_107_34
timestamp 1676037725
transform 1 0 4232 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_46
timestamp 1676037725
transform 1 0 5336 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_107_54
timestamp 1676037725
transform 1 0 6072 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_107_57
timestamp 1676037725
transform 1 0 6348 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_69
timestamp 1676037725
transform 1 0 7452 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_107_77
timestamp 1676037725
transform 1 0 8188 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_107_82
timestamp 1676037725
transform 1 0 8648 0 -1 60928
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_107_90
timestamp 1676037725
transform 1 0 9384 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_102
timestamp 1676037725
transform 1 0 10488 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_107_110
timestamp 1676037725
transform 1 0 11224 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_107_113
timestamp 1676037725
transform 1 0 11500 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_125
timestamp 1676037725
transform 1 0 12604 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_107_133
timestamp 1676037725
transform 1 0 13340 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_107_138
timestamp 1676037725
transform 1 0 13800 0 -1 60928
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_107_146
timestamp 1676037725
transform 1 0 14536 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_162
timestamp 1676037725
transform 1 0 16008 0 -1 60928
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_107_169
timestamp 1676037725
transform 1 0 16652 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_181
timestamp 1676037725
transform 1 0 17756 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_107_193
timestamp 1676037725
transform 1 0 18860 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_107_197
timestamp 1676037725
transform 1 0 19228 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_202
timestamp 1676037725
transform 1 0 19688 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_214
timestamp 1676037725
transform 1 0 20792 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_107_222
timestamp 1676037725
transform 1 0 21528 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_107_225
timestamp 1676037725
transform 1 0 21804 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_107_236
timestamp 1676037725
transform 1 0 22816 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_107_244
timestamp 1676037725
transform 1 0 23552 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_107_252
timestamp 1676037725
transform 1 0 24288 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_107_258
timestamp 1676037725
transform 1 0 24840 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_270
timestamp 1676037725
transform 1 0 25944 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_107_278
timestamp 1676037725
transform 1 0 26680 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_107_281
timestamp 1676037725
transform 1 0 26956 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_107_285
timestamp 1676037725
transform 1 0 27324 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_290
timestamp 1676037725
transform 1 0 27784 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_306
timestamp 1676037725
transform 1 0 29256 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_322
timestamp 1676037725
transform 1 0 30728 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_107_334
timestamp 1676037725
transform 1 0 31832 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_107_337
timestamp 1676037725
transform 1 0 32108 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_349
timestamp 1676037725
transform 1 0 33212 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_361
timestamp 1676037725
transform 1 0 34316 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_373
timestamp 1676037725
transform 1 0 35420 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_107_381
timestamp 1676037725
transform 1 0 36156 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_107_386
timestamp 1676037725
transform 1 0 36616 0 -1 60928
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_107_393
timestamp 1676037725
transform 1 0 37260 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_405
timestamp 1676037725
transform 1 0 38364 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_417
timestamp 1676037725
transform 1 0 39468 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_429
timestamp 1676037725
transform 1 0 40572 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_107_437
timestamp 1676037725
transform 1 0 41308 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_107_442
timestamp 1676037725
transform 1 0 41768 0 -1 60928
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_107_449
timestamp 1676037725
transform 1 0 42412 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_461
timestamp 1676037725
transform 1 0 43516 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_473
timestamp 1676037725
transform 1 0 44620 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_485
timestamp 1676037725
transform 1 0 45724 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_107_493
timestamp 1676037725
transform 1 0 46460 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_107_498
timestamp 1676037725
transform 1 0 46920 0 -1 60928
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_107_505
timestamp 1676037725
transform 1 0 47564 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_517
timestamp 1676037725
transform 1 0 48668 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_107_529
timestamp 1676037725
transform 1 0 49772 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_107_533
timestamp 1676037725
transform 1 0 50140 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_538
timestamp 1676037725
transform 1 0 50600 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_550
timestamp 1676037725
transform 1 0 51704 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_107_558
timestamp 1676037725
transform 1 0 52440 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_107_561
timestamp 1676037725
transform 1 0 52716 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_107_567
timestamp 1676037725
transform 1 0 53268 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_107_579
timestamp 1676037725
transform 1 0 54372 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_107_586
timestamp 1676037725
transform 1 0 55016 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_107_594
timestamp 1676037725
transform 1 0 55752 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_107_602
timestamp 1676037725
transform 1 0 56488 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_107_610
timestamp 1676037725
transform 1 0 57224 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_107_617
timestamp 1676037725
transform 1 0 57868 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_107_623
timestamp 1676037725
transform 1 0 58420 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_108_3
timestamp 1676037725
transform 1 0 1380 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_14
timestamp 1676037725
transform 1 0 2392 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_24
timestamp 1676037725
transform 1 0 3312 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_29
timestamp 1676037725
transform 1 0 3772 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_33
timestamp 1676037725
transform 1 0 4140 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_38
timestamp 1676037725
transform 1 0 4600 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_46
timestamp 1676037725
transform 1 0 5336 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_108_54
timestamp 1676037725
transform 1 0 6072 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_108_57
timestamp 1676037725
transform 1 0 6348 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_108_66
timestamp 1676037725
transform 1 0 7176 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_108_76
timestamp 1676037725
transform 1 0 8096 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_108_85
timestamp 1676037725
transform 1 0 8924 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_89
timestamp 1676037725
transform 1 0 9292 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_94
timestamp 1676037725
transform 1 0 9752 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_102
timestamp 1676037725
transform 1 0 10488 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_108_110
timestamp 1676037725
transform 1 0 11224 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_113
timestamp 1676037725
transform 1 0 11500 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_117
timestamp 1676037725
transform 1 0 11868 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_122
timestamp 1676037725
transform 1 0 12328 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_108_132
timestamp 1676037725
transform 1 0 13248 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_108_141
timestamp 1676037725
transform 1 0 14076 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_149
timestamp 1676037725
transform 1 0 14812 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_108_156
timestamp 1676037725
transform 1 0 15456 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_108_166
timestamp 1676037725
transform 1 0 16376 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_169
timestamp 1676037725
transform 1 0 16652 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_173
timestamp 1676037725
transform 1 0 17020 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_178
timestamp 1676037725
transform 1 0 17480 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_186
timestamp 1676037725
transform 1 0 18216 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_108_194
timestamp 1676037725
transform 1 0 18952 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_197
timestamp 1676037725
transform 1 0 19228 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_201
timestamp 1676037725
transform 1 0 19596 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_206
timestamp 1676037725
transform 1 0 20056 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_214
timestamp 1676037725
transform 1 0 20792 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_108_222
timestamp 1676037725
transform 1 0 21528 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_225
timestamp 1676037725
transform 1 0 21804 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_229
timestamp 1676037725
transform 1 0 22172 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_108_236
timestamp 1676037725
transform 1 0 22816 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_108_244
timestamp 1676037725
transform 1 0 23552 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_108_250
timestamp 1676037725
transform 1 0 24104 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_108_253
timestamp 1676037725
transform 1 0 24380 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_261
timestamp 1676037725
transform 1 0 25116 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_268
timestamp 1676037725
transform 1 0 25760 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_276
timestamp 1676037725
transform 1 0 26496 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_108_281
timestamp 1676037725
transform 1 0 26956 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_289
timestamp 1676037725
transform 1 0 27692 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_293
timestamp 1676037725
transform 1 0 28060 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_108_300
timestamp 1676037725
transform 1 0 28704 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_108_309
timestamp 1676037725
transform 1 0 29532 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_108_317
timestamp 1676037725
transform 1 0 30268 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_325
timestamp 1676037725
transform 1 0 31004 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_332
timestamp 1676037725
transform 1 0 31648 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_108_337
timestamp 1676037725
transform 1 0 32108 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_345
timestamp 1676037725
transform 1 0 32844 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_353
timestamp 1676037725
transform 1 0 33580 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_108_361
timestamp 1676037725
transform 1 0 34316 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_108_365
timestamp 1676037725
transform 1 0 34684 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_371
timestamp 1676037725
transform 1 0 35236 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_379
timestamp 1676037725
transform 1 0 35972 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_387
timestamp 1676037725
transform 1 0 36708 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_391
timestamp 1676037725
transform 1 0 37076 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_108_393
timestamp 1676037725
transform 1 0 37260 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_399
timestamp 1676037725
transform 1 0 37812 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_407
timestamp 1676037725
transform 1 0 38548 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_415
timestamp 1676037725
transform 1 0 39284 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_419
timestamp 1676037725
transform 1 0 39652 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_108_421
timestamp 1676037725
transform 1 0 39836 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_427
timestamp 1676037725
transform 1 0 40388 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_435
timestamp 1676037725
transform 1 0 41124 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_443
timestamp 1676037725
transform 1 0 41860 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_447
timestamp 1676037725
transform 1 0 42228 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_108_449
timestamp 1676037725
transform 1 0 42412 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_457
timestamp 1676037725
transform 1 0 43148 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_465
timestamp 1676037725
transform 1 0 43884 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_108_473
timestamp 1676037725
transform 1 0 44620 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_108_477
timestamp 1676037725
transform 1 0 44988 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_483
timestamp 1676037725
transform 1 0 45540 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_491
timestamp 1676037725
transform 1 0 46276 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_499
timestamp 1676037725
transform 1 0 47012 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_503
timestamp 1676037725
transform 1 0 47380 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_108_505
timestamp 1676037725
transform 1 0 47564 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_511
timestamp 1676037725
transform 1 0 48116 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_519
timestamp 1676037725
transform 1 0 48852 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_527
timestamp 1676037725
transform 1 0 49588 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_531
timestamp 1676037725
transform 1 0 49956 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_108_533
timestamp 1676037725
transform 1 0 50140 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_541
timestamp 1676037725
transform 1 0 50876 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_549
timestamp 1676037725
transform 1 0 51612 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_108_557
timestamp 1676037725
transform 1 0 52348 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_108_561
timestamp 1676037725
transform 1 0 52716 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_565
timestamp 1676037725
transform 1 0 53084 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_572
timestamp 1676037725
transform 1 0 53728 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_108_580
timestamp 1676037725
transform 1 0 54464 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_108_589
timestamp 1676037725
transform 1 0 55292 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_597
timestamp 1676037725
transform 1 0 56028 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_108_607
timestamp 1676037725
transform 1 0 56948 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_615
timestamp 1676037725
transform 1 0 57684 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_108_617
timestamp 1676037725
transform 1 0 57868 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_108_623
timestamp 1676037725
transform 1 0 58420 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1676037725
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1676037725
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1676037725
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1676037725
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1676037725
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1676037725
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1676037725
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1676037725
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1676037725
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1676037725
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1676037725
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1676037725
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1676037725
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1676037725
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1676037725
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1676037725
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1676037725
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1676037725
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1676037725
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1676037725
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1676037725
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1676037725
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1676037725
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1676037725
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1676037725
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1676037725
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1676037725
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1676037725
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1676037725
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1676037725
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1676037725
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1676037725
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1676037725
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1676037725
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1676037725
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1676037725
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1676037725
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1676037725
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1676037725
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1676037725
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1676037725
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1676037725
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1676037725
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1676037725
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1676037725
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1676037725
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1676037725
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1676037725
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1676037725
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1676037725
transform -1 0 58880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1676037725
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1676037725
transform -1 0 58880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1676037725
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1676037725
transform -1 0 58880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1676037725
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1676037725
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1676037725
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1676037725
transform -1 0 58880 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1676037725
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1676037725
transform -1 0 58880 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1676037725
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1676037725
transform -1 0 58880 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1676037725
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1676037725
transform -1 0 58880 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1676037725
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1676037725
transform -1 0 58880 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1676037725
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1676037725
transform -1 0 58880 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1676037725
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1676037725
transform -1 0 58880 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1676037725
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1676037725
transform -1 0 58880 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1676037725
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1676037725
transform -1 0 58880 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1676037725
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1676037725
transform -1 0 58880 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1676037725
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1676037725
transform -1 0 58880 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1676037725
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1676037725
transform -1 0 58880 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1676037725
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1676037725
transform -1 0 58880 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1676037725
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1676037725
transform -1 0 58880 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1676037725
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1676037725
transform -1 0 58880 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1676037725
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1676037725
transform -1 0 58880 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1676037725
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1676037725
transform -1 0 58880 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1676037725
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1676037725
transform -1 0 58880 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1676037725
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1676037725
transform -1 0 58880 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1676037725
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1676037725
transform -1 0 58880 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1676037725
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1676037725
transform -1 0 58880 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1676037725
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1676037725
transform -1 0 58880 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1676037725
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1676037725
transform -1 0 58880 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1676037725
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1676037725
transform -1 0 58880 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1676037725
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1676037725
transform -1 0 58880 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1676037725
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1676037725
transform -1 0 58880 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1676037725
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1676037725
transform -1 0 58880 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1676037725
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1676037725
transform -1 0 58880 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1676037725
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1676037725
transform -1 0 58880 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1676037725
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1676037725
transform -1 0 58880 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1676037725
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1676037725
transform -1 0 58880 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1676037725
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1676037725
transform -1 0 58880 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1676037725
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1676037725
transform -1 0 58880 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1676037725
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1676037725
transform -1 0 58880 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1676037725
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1676037725
transform -1 0 58880 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1676037725
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1676037725
transform -1 0 58880 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1676037725
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1676037725
transform -1 0 58880 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1676037725
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1676037725
transform -1 0 58880 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_214
timestamp 1676037725
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_215
timestamp 1676037725
transform -1 0 58880 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_216
timestamp 1676037725
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_217
timestamp 1676037725
transform -1 0 58880 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1676037725
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1676037725
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1676037725
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1676037725
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1676037725
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1676037725
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1676037725
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1676037725
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1676037725
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1676037725
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1676037725
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1676037725
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1676037725
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1676037725
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1676037725
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1676037725
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1676037725
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1676037725
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1676037725
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1676037725
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1676037725
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1676037725
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1676037725
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1676037725
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1676037725
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1676037725
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1676037725
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1676037725
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1676037725
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1676037725
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1676037725
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1676037725
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1676037725
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1676037725
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1676037725
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1676037725
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1676037725
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1676037725
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1676037725
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1676037725
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1676037725
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1676037725
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1676037725
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1676037725
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1676037725
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1676037725
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1676037725
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1676037725
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1676037725
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1676037725
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1676037725
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1676037725
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1676037725
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1676037725
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1676037725
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1676037725
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1676037725
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1676037725
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1676037725
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1676037725
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1676037725
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1676037725
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1676037725
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1676037725
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1676037725
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1676037725
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1676037725
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1676037725
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1676037725
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1676037725
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1676037725
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1676037725
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1676037725
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1676037725
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1676037725
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1676037725
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1676037725
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1676037725
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1676037725
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1676037725
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1676037725
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1676037725
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1676037725
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1676037725
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1676037725
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1676037725
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1676037725
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1676037725
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1676037725
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1676037725
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1676037725
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1676037725
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1676037725
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1676037725
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1676037725
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1676037725
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1676037725
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1676037725
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1676037725
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1676037725
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1676037725
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1676037725
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1676037725
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1676037725
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1676037725
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1676037725
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1676037725
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1676037725
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1676037725
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1676037725
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1676037725
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1676037725
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1676037725
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1676037725
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1676037725
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1676037725
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1676037725
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1676037725
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1676037725
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1676037725
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1676037725
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1676037725
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1676037725
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1676037725
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1676037725
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1676037725
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1676037725
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1676037725
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1676037725
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1676037725
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1676037725
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1676037725
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1676037725
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1676037725
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1676037725
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1676037725
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1676037725
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1676037725
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1676037725
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1676037725
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1676037725
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1676037725
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1676037725
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1676037725
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1676037725
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1676037725
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1676037725
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1676037725
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1676037725
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1676037725
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1676037725
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1676037725
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1676037725
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1676037725
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1676037725
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1676037725
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1676037725
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1676037725
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1676037725
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1676037725
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1676037725
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1676037725
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1676037725
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1676037725
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1676037725
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1676037725
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1676037725
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1676037725
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1676037725
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1676037725
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1676037725
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1676037725
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1676037725
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1676037725
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1676037725
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1676037725
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1676037725
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1676037725
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1676037725
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1676037725
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1676037725
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1676037725
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1676037725
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1676037725
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1676037725
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1676037725
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1676037725
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1676037725
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1676037725
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1676037725
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1676037725
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1676037725
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1676037725
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1676037725
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1676037725
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1676037725
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1676037725
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1676037725
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1676037725
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1676037725
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1676037725
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1676037725
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1676037725
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1676037725
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1676037725
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1676037725
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1676037725
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1676037725
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1676037725
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1676037725
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1676037725
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1676037725
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1676037725
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1676037725
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1676037725
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1676037725
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1676037725
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1676037725
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1676037725
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1676037725
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1676037725
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1676037725
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1676037725
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1676037725
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1676037725
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1676037725
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1676037725
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1676037725
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1676037725
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1676037725
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1676037725
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1676037725
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1676037725
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1676037725
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1676037725
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1676037725
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1676037725
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1676037725
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1676037725
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1676037725
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1676037725
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1676037725
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1676037725
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1676037725
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1676037725
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1676037725
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1676037725
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1676037725
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1676037725
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1676037725
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1676037725
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1676037725
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1676037725
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1676037725
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1676037725
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1676037725
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1676037725
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1676037725
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1676037725
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1676037725
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1676037725
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1676037725
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1676037725
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1676037725
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1676037725
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1676037725
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1676037725
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1676037725
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1676037725
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1676037725
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1676037725
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1676037725
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1676037725
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1676037725
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1676037725
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1676037725
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1676037725
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1676037725
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1676037725
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1676037725
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1676037725
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1676037725
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1676037725
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1676037725
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1676037725
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1676037725
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1676037725
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1676037725
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1676037725
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1676037725
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1676037725
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1676037725
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1676037725
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1676037725
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1676037725
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1676037725
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1676037725
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1676037725
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1676037725
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1676037725
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1676037725
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1676037725
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1676037725
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1676037725
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1676037725
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1676037725
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1676037725
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1676037725
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1676037725
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1676037725
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1676037725
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1676037725
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1676037725
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1676037725
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1676037725
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1676037725
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1676037725
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1676037725
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1676037725
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1676037725
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1676037725
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1676037725
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1676037725
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1676037725
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1676037725
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1676037725
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1676037725
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1676037725
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1676037725
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1676037725
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1676037725
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1676037725
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1676037725
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1676037725
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1676037725
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1676037725
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1676037725
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1676037725
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1676037725
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1676037725
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1676037725
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1676037725
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1676037725
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1676037725
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1676037725
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1676037725
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1676037725
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1676037725
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1676037725
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1676037725
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1676037725
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1676037725
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1676037725
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1676037725
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1676037725
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1676037725
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1676037725
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1676037725
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1676037725
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1676037725
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1676037725
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1676037725
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1676037725
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1676037725
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1676037725
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1676037725
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1676037725
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1676037725
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1676037725
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1676037725
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1676037725
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1676037725
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1676037725
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1676037725
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1676037725
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1676037725
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1676037725
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1676037725
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1676037725
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1676037725
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1676037725
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1676037725
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1676037725
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1676037725
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1676037725
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1676037725
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1676037725
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1676037725
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1676037725
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1676037725
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1676037725
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1676037725
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1676037725
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1676037725
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1676037725
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1676037725
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1676037725
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1676037725
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1676037725
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1676037725
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1676037725
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1676037725
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1676037725
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1676037725
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1676037725
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1676037725
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1676037725
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1676037725
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1676037725
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1676037725
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1676037725
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1676037725
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1676037725
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1676037725
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1676037725
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1676037725
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1676037725
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1676037725
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1676037725
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1676037725
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1676037725
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1676037725
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1676037725
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1676037725
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1676037725
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1676037725
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1676037725
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1676037725
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1676037725
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1676037725
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1676037725
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1676037725
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1676037725
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1676037725
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1676037725
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1676037725
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1676037725
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1676037725
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1676037725
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1676037725
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1676037725
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1676037725
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1676037725
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1676037725
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1676037725
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1676037725
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1676037725
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1676037725
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1676037725
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1676037725
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1676037725
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1676037725
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1676037725
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1676037725
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1676037725
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1676037725
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1676037725
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1676037725
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1676037725
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1676037725
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1676037725
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1676037725
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1676037725
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1676037725
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1676037725
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1676037725
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1676037725
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1676037725
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1676037725
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1676037725
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1676037725
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1676037725
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1676037725
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1676037725
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1676037725
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1676037725
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1676037725
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1676037725
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1676037725
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1676037725
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1676037725
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1676037725
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1676037725
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1676037725
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1676037725
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1676037725
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1676037725
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1676037725
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1676037725
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1676037725
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1676037725
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1676037725
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1676037725
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1676037725
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1676037725
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1676037725
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1676037725
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1676037725
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1676037725
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1676037725
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1676037725
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1676037725
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1676037725
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1676037725
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1676037725
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1676037725
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1676037725
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1676037725
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1676037725
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1676037725
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1676037725
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1676037725
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1676037725
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1676037725
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1676037725
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1676037725
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1676037725
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1676037725
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1676037725
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1676037725
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1676037725
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1676037725
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1676037725
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1676037725
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1676037725
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1676037725
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1676037725
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1676037725
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1676037725
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1676037725
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1676037725
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1676037725
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1676037725
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1676037725
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1676037725
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1676037725
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1676037725
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1676037725
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1676037725
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1676037725
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1676037725
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1676037725
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1676037725
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1676037725
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1676037725
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1676037725
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1676037725
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1676037725
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1676037725
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1676037725
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1676037725
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1676037725
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1676037725
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1676037725
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1676037725
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1676037725
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1676037725
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1676037725
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1676037725
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1676037725
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1676037725
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1676037725
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1676037725
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1676037725
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1676037725
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1676037725
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1676037725
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1676037725
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1676037725
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1676037725
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1676037725
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1676037725
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1676037725
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1676037725
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1676037725
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1676037725
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1676037725
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1676037725
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1676037725
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1676037725
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1676037725
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1676037725
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1676037725
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1676037725
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1676037725
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1676037725
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1676037725
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1676037725
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1676037725
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1676037725
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1676037725
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1676037725
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1676037725
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1676037725
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1676037725
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1676037725
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1676037725
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1676037725
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1676037725
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1676037725
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1676037725
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1676037725
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1676037725
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1676037725
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1676037725
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1676037725
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1676037725
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1676037725
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1676037725
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1676037725
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1676037725
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1676037725
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1676037725
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1676037725
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1676037725
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1676037725
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1676037725
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1676037725
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1676037725
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1676037725
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1676037725
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1676037725
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1676037725
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1676037725
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1676037725
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1676037725
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1676037725
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1676037725
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1676037725
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1676037725
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1676037725
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1676037725
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1676037725
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1676037725
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1676037725
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1676037725
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1676037725
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1676037725
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1676037725
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1676037725
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1676037725
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1676037725
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1676037725
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1676037725
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1676037725
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1676037725
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1676037725
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1676037725
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1676037725
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1676037725
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1676037725
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1676037725
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1676037725
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1676037725
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1676037725
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1676037725
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1676037725
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1676037725
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1676037725
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1676037725
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1676037725
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1676037725
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1676037725
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1676037725
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1676037725
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1676037725
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1676037725
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1676037725
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1676037725
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1676037725
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1676037725
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1676037725
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1676037725
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1676037725
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1676037725
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1676037725
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1676037725
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1676037725
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1676037725
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1676037725
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1676037725
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1676037725
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1676037725
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1676037725
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1676037725
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1676037725
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1676037725
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1676037725
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1676037725
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1676037725
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1676037725
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1676037725
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1676037725
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1676037725
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1676037725
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1676037725
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1676037725
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1676037725
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1676037725
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1676037725
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1676037725
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1676037725
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1676037725
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1676037725
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1676037725
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1676037725
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1676037725
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1676037725
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1676037725
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1676037725
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1676037725
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1676037725
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1676037725
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1676037725
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1676037725
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1676037725
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1676037725
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1676037725
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1676037725
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1676037725
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1676037725
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1676037725
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1676037725
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1676037725
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1676037725
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1676037725
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1676037725
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1676037725
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1676037725
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1676037725
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1676037725
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1676037725
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1676037725
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1676037725
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1676037725
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1676037725
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1676037725
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1676037725
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1676037725
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1676037725
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1676037725
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1676037725
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1676037725
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1676037725
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1676037725
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1676037725
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1676037725
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1676037725
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1676037725
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1676037725
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1676037725
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1676037725
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1676037725
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1676037725
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1676037725
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1676037725
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1676037725
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1676037725
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1676037725
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1676037725
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1676037725
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1676037725
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1676037725
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1676037725
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1676037725
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1676037725
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1676037725
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1676037725
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1676037725
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1676037725
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1676037725
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1676037725
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1676037725
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1676037725
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1676037725
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1676037725
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1676037725
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1676037725
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1676037725
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1676037725
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1676037725
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1676037725
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1676037725
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1676037725
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1676037725
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1676037725
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1676037725
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1676037725
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1676037725
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1676037725
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1348
timestamp 1676037725
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1349
timestamp 1676037725
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1350
timestamp 1676037725
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1351
timestamp 1676037725
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1352
timestamp 1676037725
transform 1 0 8832 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1353
timestamp 1676037725
transform 1 0 13984 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1354
timestamp 1676037725
transform 1 0 19136 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1355
timestamp 1676037725
transform 1 0 24288 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1356
timestamp 1676037725
transform 1 0 29440 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1357
timestamp 1676037725
transform 1 0 34592 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1358
timestamp 1676037725
transform 1 0 39744 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1359
timestamp 1676037725
transform 1 0 44896 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1360
timestamp 1676037725
transform 1 0 50048 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1361
timestamp 1676037725
transform 1 0 55200 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1362
timestamp 1676037725
transform 1 0 6256 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1363
timestamp 1676037725
transform 1 0 11408 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1364
timestamp 1676037725
transform 1 0 16560 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1365
timestamp 1676037725
transform 1 0 21712 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1366
timestamp 1676037725
transform 1 0 26864 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1367
timestamp 1676037725
transform 1 0 32016 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1368
timestamp 1676037725
transform 1 0 37168 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1369
timestamp 1676037725
transform 1 0 42320 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1370
timestamp 1676037725
transform 1 0 47472 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1371
timestamp 1676037725
transform 1 0 52624 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1372
timestamp 1676037725
transform 1 0 57776 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1373
timestamp 1676037725
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1374
timestamp 1676037725
transform 1 0 8832 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1375
timestamp 1676037725
transform 1 0 13984 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1376
timestamp 1676037725
transform 1 0 19136 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1377
timestamp 1676037725
transform 1 0 24288 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1378
timestamp 1676037725
transform 1 0 29440 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1379
timestamp 1676037725
transform 1 0 34592 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1380
timestamp 1676037725
transform 1 0 39744 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1381
timestamp 1676037725
transform 1 0 44896 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1382
timestamp 1676037725
transform 1 0 50048 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1383
timestamp 1676037725
transform 1 0 55200 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1384
timestamp 1676037725
transform 1 0 6256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1385
timestamp 1676037725
transform 1 0 11408 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1386
timestamp 1676037725
transform 1 0 16560 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1387
timestamp 1676037725
transform 1 0 21712 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1388
timestamp 1676037725
transform 1 0 26864 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1389
timestamp 1676037725
transform 1 0 32016 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1390
timestamp 1676037725
transform 1 0 37168 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1391
timestamp 1676037725
transform 1 0 42320 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1392
timestamp 1676037725
transform 1 0 47472 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1393
timestamp 1676037725
transform 1 0 52624 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1394
timestamp 1676037725
transform 1 0 57776 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1395
timestamp 1676037725
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1396
timestamp 1676037725
transform 1 0 8832 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1397
timestamp 1676037725
transform 1 0 13984 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1398
timestamp 1676037725
transform 1 0 19136 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1399
timestamp 1676037725
transform 1 0 24288 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1400
timestamp 1676037725
transform 1 0 29440 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1401
timestamp 1676037725
transform 1 0 34592 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1402
timestamp 1676037725
transform 1 0 39744 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1403
timestamp 1676037725
transform 1 0 44896 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1404
timestamp 1676037725
transform 1 0 50048 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1405
timestamp 1676037725
transform 1 0 55200 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1406
timestamp 1676037725
transform 1 0 6256 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1407
timestamp 1676037725
transform 1 0 11408 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1408
timestamp 1676037725
transform 1 0 16560 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1409
timestamp 1676037725
transform 1 0 21712 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1410
timestamp 1676037725
transform 1 0 26864 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1411
timestamp 1676037725
transform 1 0 32016 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1412
timestamp 1676037725
transform 1 0 37168 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1413
timestamp 1676037725
transform 1 0 42320 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1414
timestamp 1676037725
transform 1 0 47472 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1415
timestamp 1676037725
transform 1 0 52624 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1416
timestamp 1676037725
transform 1 0 57776 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1417
timestamp 1676037725
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1418
timestamp 1676037725
transform 1 0 6256 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1419
timestamp 1676037725
transform 1 0 8832 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1420
timestamp 1676037725
transform 1 0 11408 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1421
timestamp 1676037725
transform 1 0 13984 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1422
timestamp 1676037725
transform 1 0 16560 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1423
timestamp 1676037725
transform 1 0 19136 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1424
timestamp 1676037725
transform 1 0 21712 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1425
timestamp 1676037725
transform 1 0 24288 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1426
timestamp 1676037725
transform 1 0 26864 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1427
timestamp 1676037725
transform 1 0 29440 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1428
timestamp 1676037725
transform 1 0 32016 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1429
timestamp 1676037725
transform 1 0 34592 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1430
timestamp 1676037725
transform 1 0 37168 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1431
timestamp 1676037725
transform 1 0 39744 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1432
timestamp 1676037725
transform 1 0 42320 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1433
timestamp 1676037725
transform 1 0 44896 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1434
timestamp 1676037725
transform 1 0 47472 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1435
timestamp 1676037725
transform 1 0 50048 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1436
timestamp 1676037725
transform 1 0 52624 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1437
timestamp 1676037725
transform 1 0 55200 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1438
timestamp 1676037725
transform 1 0 57776 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0449_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 40756 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0450_
timestamp 1676037725
transform 1 0 23828 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0451_
timestamp 1676037725
transform 1 0 23828 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0452_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 38824 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0453_
timestamp 1676037725
transform 1 0 44344 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0454_
timestamp 1676037725
transform 1 0 41768 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0455_
timestamp 1676037725
transform 1 0 42780 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0456_
timestamp 1676037725
transform 1 0 14168 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0457_
timestamp 1676037725
transform 1 0 13984 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0458_
timestamp 1676037725
transform 1 0 16100 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor4b_4  _0459_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15640 0 1 9792
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_4  _0460_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7544 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2b_1  _0461_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2852 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _0462_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15180 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor4b_4  _0463_
timestamp 1676037725
transform 1 0 18216 0 -1 8704
box -38 -48 1786 592
use sky130_fd_sc_hd__or3_4  _0464_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12880 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_4  _0465_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15180 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_1  _0466_
timestamp 1676037725
transform 1 0 9476 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_2  _0467_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24932 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor4b_4  _0468_
timestamp 1676037725
transform 1 0 16376 0 1 7616
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2b_1  _0469_
timestamp 1676037725
transform 1 0 2484 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_4  _0470_
timestamp 1676037725
transform 1 0 16836 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_1  _0471_
timestamp 1676037725
transform 1 0 10672 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_4  _0472_
timestamp 1676037725
transform 1 0 16836 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_1  _0473_
timestamp 1676037725
transform 1 0 2484 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_2  _0474_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_1  _0475_
timestamp 1676037725
transform 1 0 11960 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0476_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13156 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor4b_4  _0477_
timestamp 1676037725
transform 1 0 16928 0 1 5440
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2b_1  _0478_
timestamp 1676037725
transform 1 0 11684 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0479_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27140 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_4  _0480_
timestamp 1676037725
transform 1 0 15180 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_1  _0481_
timestamp 1676037725
transform 1 0 10856 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_2  _0482_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23460 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__or3_4  _0483_
timestamp 1676037725
transform 1 0 12788 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_4  _0484_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__nand2b_2  _0485_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2024 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _0486_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18400 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__nand2b_1  _0487_
timestamp 1676037725
transform 1 0 2484 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_4  _0488_
timestamp 1676037725
transform 1 0 15548 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__nand2b_1  _0489_
timestamp 1676037725
transform 1 0 9292 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2_4  _0490_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24656 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_4  _0491_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32384 0 1 56576
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _0492_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 37260 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_4  _0493_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32568 0 1 42432
box -38 -48 1602 592
use sky130_fd_sc_hd__a221o_1  _0494_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33304 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0495_
timestamp 1676037725
transform 1 0 32936 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _0496_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29716 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0497_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29716 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0498_
timestamp 1676037725
transform 1 0 28152 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _0499_
timestamp 1676037725
transform 1 0 31372 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _0500_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 30912 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _0501_
timestamp 1676037725
transform 1 0 27140 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0502_
timestamp 1676037725
transform 1 0 32292 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0503_
timestamp 1676037725
transform 1 0 43608 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_4  _0504_
timestamp 1676037725
transform 1 0 32016 0 1 59840
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _0505_
timestamp 1676037725
transform 1 0 31832 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0506_
timestamp 1676037725
transform 1 0 35328 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0507_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32384 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_4  _0508_
timestamp 1676037725
transform 1 0 32660 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0509_
timestamp 1676037725
transform 1 0 38088 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0510_
timestamp 1676037725
transform 1 0 38548 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_4  _0511_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24748 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_1  _0512_
timestamp 1676037725
transform 1 0 53084 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0513_
timestamp 1676037725
transform 1 0 33672 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0514_
timestamp 1676037725
transform 1 0 33764 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0515_
timestamp 1676037725
transform 1 0 34776 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0516_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 34960 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0517_
timestamp 1676037725
transform 1 0 37076 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_4  _0518_
timestamp 1676037725
transform 1 0 17388 0 1 59840
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_1  _0519_
timestamp 1676037725
transform 1 0 36248 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0520_
timestamp 1676037725
transform 1 0 37444 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _0521_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35696 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _0522_
timestamp 1676037725
transform 1 0 37444 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _0523_
timestamp 1676037725
transform 1 0 37996 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0524_
timestamp 1676037725
transform 1 0 34040 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _0525_
timestamp 1676037725
transform 1 0 17020 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0526_
timestamp 1676037725
transform 1 0 18676 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_4  _0527_
timestamp 1676037725
transform 1 0 35144 0 1 57664
box -38 -48 1602 592
use sky130_fd_sc_hd__or3_4  _0528_
timestamp 1676037725
transform 1 0 19412 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_2  _0529_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14720 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _0530_
timestamp 1676037725
transform 1 0 27416 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _0531_
timestamp 1676037725
transform 1 0 29716 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_2  _0532_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9660 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0533_
timestamp 1676037725
transform 1 0 36340 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_4  _0534_
timestamp 1676037725
transform 1 0 37444 0 -1 58752
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_2  _0535_
timestamp 1676037725
transform 1 0 23184 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0536_
timestamp 1676037725
transform 1 0 24564 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0537_
timestamp 1676037725
transform 1 0 24104 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0538_
timestamp 1676037725
transform 1 0 24748 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0539_
timestamp 1676037725
transform 1 0 22724 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0540_
timestamp 1676037725
transform 1 0 21528 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0541_
timestamp 1676037725
transform 1 0 20792 0 -1 59840
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_4  _0542_
timestamp 1676037725
transform 1 0 21528 0 1 59840
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_1  _0543_
timestamp 1676037725
transform 1 0 22540 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _0544_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22816 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _0545_
timestamp 1676037725
transform 1 0 22264 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _0546_
timestamp 1676037725
transform 1 0 19412 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0547_
timestamp 1676037725
transform 1 0 19320 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0548_
timestamp 1676037725
transform 1 0 53636 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0549_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20608 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0550_
timestamp 1676037725
transform 1 0 18400 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0551_
timestamp 1676037725
transform 1 0 19044 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0552_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20056 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _0553_
timestamp 1676037725
transform 1 0 20148 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0554_
timestamp 1676037725
transform 1 0 20884 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0555_
timestamp 1676037725
transform 1 0 21988 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0556_
timestamp 1676037725
transform 1 0 53820 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0557_
timestamp 1676037725
transform 1 0 2024 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0558_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2576 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_4  _0559_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15640 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_2  _0560_
timestamp 1676037725
transform 1 0 19320 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0561_
timestamp 1676037725
transform 1 0 20148 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__or3_4  _0562_
timestamp 1676037725
transform 1 0 21804 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_4  _0563_
timestamp 1676037725
transform 1 0 14812 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_2  _0564_
timestamp 1676037725
transform 1 0 20424 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0565_
timestamp 1676037725
transform 1 0 22172 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _0566_
timestamp 1676037725
transform 1 0 21344 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0567_
timestamp 1676037725
transform 1 0 40020 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0568_
timestamp 1676037725
transform 1 0 2300 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _0569_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22540 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _0570_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22540 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0571_
timestamp 1676037725
transform 1 0 21712 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_4  _0572_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25024 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_2  _0573_
timestamp 1676037725
transform 1 0 22080 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0574_
timestamp 1676037725
transform 1 0 22908 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0575_
timestamp 1676037725
transform 1 0 2484 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0576_
timestamp 1676037725
transform 1 0 23276 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0577_
timestamp 1676037725
transform 1 0 40204 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0578_
timestamp 1676037725
transform 1 0 23736 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _0579_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_4  _0580_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26496 0 1 6528
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _0581_
timestamp 1676037725
transform 1 0 20884 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_4  _0582_
timestamp 1676037725
transform 1 0 40112 0 1 3264
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_2  _0583_
timestamp 1676037725
transform 1 0 2024 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0584_
timestamp 1676037725
transform 1 0 40572 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _0585_
timestamp 1676037725
transform 1 0 20516 0 1 51136
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _0586_
timestamp 1676037725
transform 1 0 21436 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0587_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31740 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0588_
timestamp 1676037725
transform 1 0 30452 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0589_
timestamp 1676037725
transform 1 0 32108 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0590_
timestamp 1676037725
transform 1 0 3680 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_4  _0591_
timestamp 1676037725
transform 1 0 5428 0 1 36992
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_1  _0592_
timestamp 1676037725
transform 1 0 27508 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0593_
timestamp 1676037725
transform 1 0 28520 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0594_
timestamp 1676037725
transform 1 0 29716 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0595_
timestamp 1676037725
transform 1 0 31096 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0596_
timestamp 1676037725
transform 1 0 32108 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0597_
timestamp 1676037725
transform 1 0 23092 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0598_
timestamp 1676037725
transform 1 0 23092 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0599_
timestamp 1676037725
transform 1 0 7360 0 1 59840
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _0600_
timestamp 1676037725
transform 1 0 7728 0 -1 52224
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _0601_
timestamp 1676037725
transform 1 0 22724 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _0602_
timestamp 1676037725
transform 1 0 27324 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_4  _0603_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25668 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_1  _0604_
timestamp 1676037725
transform 1 0 23460 0 1 59840
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_4  _0605_
timestamp 1676037725
transform 1 0 23736 0 -1 56576
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _0606_
timestamp 1676037725
transform 1 0 26220 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_2  _0607_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25024 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _0608_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0609_
timestamp 1676037725
transform 1 0 23828 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0610_
timestamp 1676037725
transform 1 0 23552 0 -1 53312
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0611_
timestamp 1676037725
transform 1 0 24932 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0612_
timestamp 1676037725
transform 1 0 22724 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _0613_
timestamp 1676037725
transform 1 0 23736 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _0614_
timestamp 1676037725
transform 1 0 40296 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0615_
timestamp 1676037725
transform 1 0 39836 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0616_
timestamp 1676037725
transform 1 0 40480 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0617_
timestamp 1676037725
transform 1 0 38456 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _0618_
timestamp 1676037725
transform 1 0 23828 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_4  _0619_
timestamp 1676037725
transform 1 0 41676 0 1 4352
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_2  _0620_
timestamp 1676037725
transform 1 0 28060 0 1 59840
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _0621_
timestamp 1676037725
transform 1 0 22816 0 1 54400
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _0622_
timestamp 1676037725
transform 1 0 42596 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0623_
timestamp 1676037725
transform 1 0 40848 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0624_
timestamp 1676037725
transform 1 0 41492 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0625_
timestamp 1676037725
transform 1 0 37444 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_4  _0626_
timestamp 1676037725
transform 1 0 42596 0 -1 3264
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_2  _0627_
timestamp 1676037725
transform 1 0 30360 0 1 59840
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _0628_
timestamp 1676037725
transform 1 0 24564 0 1 55488
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _0629_
timestamp 1676037725
transform 1 0 40848 0 -1 56576
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_1  _0630_
timestamp 1676037725
transform 1 0 41032 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0631_
timestamp 1676037725
transform 1 0 40848 0 -1 16320
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _0632_
timestamp 1676037725
transform 1 0 42688 0 -1 4352
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_1  _0633_
timestamp 1676037725
transform 1 0 29716 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0634_
timestamp 1676037725
transform 1 0 28796 0 -1 56576
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_4  _0635_
timestamp 1676037725
transform 1 0 32292 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_4  _0636_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31740 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0637_
timestamp 1676037725
transform 1 0 41492 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0638_
timestamp 1676037725
transform 1 0 42596 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_2  _0639_
timestamp 1676037725
transform 1 0 29440 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_4  _0640_
timestamp 1676037725
transform 1 0 41676 0 1 59840
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_2  _0641_
timestamp 1676037725
transform 1 0 42596 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_2  _0642_
timestamp 1676037725
transform 1 0 32292 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_4  _0643_
timestamp 1676037725
transform 1 0 40848 0 1 58752
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_1  _0644_
timestamp 1676037725
transform 1 0 42412 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0645_
timestamp 1676037725
transform 1 0 41124 0 1 11968
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _0646_
timestamp 1676037725
transform 1 0 40848 0 -1 58752
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_1  _0647_
timestamp 1676037725
transform 1 0 40020 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0648_
timestamp 1676037725
transform 1 0 42596 0 -1 11968
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _0649_
timestamp 1676037725
transform 1 0 42596 0 -1 59840
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_4  _0650_
timestamp 1676037725
transform 1 0 42780 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__a211o_4  _0651_
timestamp 1676037725
transform 1 0 30452 0 -1 14144
box -38 -48 1326 592
use sky130_fd_sc_hd__a211o_4  _0652_
timestamp 1676037725
transform 1 0 15088 0 -1 10880
box -38 -48 1326 592
use sky130_fd_sc_hd__a211o_2  _0653_
timestamp 1676037725
transform 1 0 13064 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_2  _0654_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0655_
timestamp 1676037725
transform 1 0 17296 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0656_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10396 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0657_
timestamp 1676037725
transform 1 0 26680 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0658_
timestamp 1676037725
transform 1 0 8004 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0659_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9384 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0660_
timestamp 1676037725
transform 1 0 8464 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0661_
timestamp 1676037725
transform 1 0 9384 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0662_
timestamp 1676037725
transform 1 0 7176 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0663_
timestamp 1676037725
transform 1 0 8924 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0664_
timestamp 1676037725
transform 1 0 8096 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0665_
timestamp 1676037725
transform 1 0 9568 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0666_
timestamp 1676037725
transform 1 0 10396 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0667_
timestamp 1676037725
transform 1 0 10120 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0668_
timestamp 1676037725
transform 1 0 8924 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0669_
timestamp 1676037725
transform 1 0 9108 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0670_
timestamp 1676037725
transform 1 0 9936 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0671_
timestamp 1676037725
transform 1 0 9108 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0672_
timestamp 1676037725
transform 1 0 10580 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0673_
timestamp 1676037725
transform 1 0 10764 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0674_
timestamp 1676037725
transform 1 0 10396 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0675_
timestamp 1676037725
transform 1 0 10580 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0676_
timestamp 1676037725
transform 1 0 12420 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0677_
timestamp 1676037725
transform 1 0 23460 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0678_
timestamp 1676037725
transform 1 0 12880 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0679_
timestamp 1676037725
transform 1 0 28612 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0680_
timestamp 1676037725
transform 1 0 14260 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0681_
timestamp 1676037725
transform 1 0 27140 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0682_
timestamp 1676037725
transform 1 0 12512 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0683_
timestamp 1676037725
transform 1 0 24564 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0684_
timestamp 1676037725
transform 1 0 11040 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0685_
timestamp 1676037725
transform 1 0 10948 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0686_
timestamp 1676037725
transform 1 0 11684 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0687_
timestamp 1676037725
transform 1 0 11684 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0688_
timestamp 1676037725
transform 1 0 12880 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0689_
timestamp 1676037725
transform 1 0 31372 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0690_
timestamp 1676037725
transform 1 0 12420 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0691_
timestamp 1676037725
transform 1 0 23092 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0692_
timestamp 1676037725
transform 1 0 13248 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0693_
timestamp 1676037725
transform 1 0 32568 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0694_
timestamp 1676037725
transform 1 0 13340 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0695_
timestamp 1676037725
transform 1 0 23460 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0696_
timestamp 1676037725
transform 1 0 14260 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0697_
timestamp 1676037725
transform 1 0 30820 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0698_
timestamp 1676037725
transform 1 0 13248 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0699_
timestamp 1676037725
transform 1 0 13156 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0700_
timestamp 1676037725
transform 1 0 14260 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0701_
timestamp 1676037725
transform 1 0 29164 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0702_
timestamp 1676037725
transform 1 0 12328 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0703_
timestamp 1676037725
transform 1 0 13156 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_2  _0704_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15364 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_4  _0705_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29716 0 1 7616
box -38 -48 1326 592
use sky130_fd_sc_hd__and2b_2  _0706_
timestamp 1676037725
transform 1 0 15640 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_4  _0707_
timestamp 1676037725
transform 1 0 29716 0 1 6528
box -38 -48 1326 592
use sky130_fd_sc_hd__and2b_1  _0708_
timestamp 1676037725
transform 1 0 13248 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0709_
timestamp 1676037725
transform 1 0 15088 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0710_
timestamp 1676037725
transform 1 0 8740 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0711_
timestamp 1676037725
transform 1 0 9200 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _0712_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 57040 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _0713_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 43700 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0714_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 36156 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0715_
timestamp 1676037725
transform 1 0 36524 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0716_
timestamp 1676037725
transform 1 0 46368 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0717_
timestamp 1676037725
transform 1 0 23644 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0718_
timestamp 1676037725
transform 1 0 19964 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0719_
timestamp 1676037725
transform 1 0 34868 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0720_
timestamp 1676037725
transform 1 0 33948 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0721_
timestamp 1676037725
transform 1 0 35972 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0722_
timestamp 1676037725
transform 1 0 37444 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0723_
timestamp 1676037725
transform 1 0 38732 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0724_
timestamp 1676037725
transform 1 0 38732 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0725_
timestamp 1676037725
transform 1 0 31372 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0726_
timestamp 1676037725
transform 1 0 32568 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0727_
timestamp 1676037725
transform 1 0 27140 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0728_
timestamp 1676037725
transform 1 0 26220 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0729_
timestamp 1676037725
transform 1 0 18492 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0730_
timestamp 1676037725
transform 1 0 45172 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0731_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 43792 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0732_
timestamp 1676037725
transform 1 0 28428 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0733_
timestamp 1676037725
transform 1 0 27784 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0734_
timestamp 1676037725
transform 1 0 32292 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0735_
timestamp 1676037725
transform 1 0 31464 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0736_
timestamp 1676037725
transform 1 0 32108 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0737_
timestamp 1676037725
transform 1 0 33304 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0738_
timestamp 1676037725
transform 1 0 37812 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0739_
timestamp 1676037725
transform 1 0 37444 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0740_
timestamp 1676037725
transform 1 0 27692 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0741_
timestamp 1676037725
transform 1 0 26312 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0742_
timestamp 1676037725
transform 1 0 29256 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0743_
timestamp 1676037725
transform 1 0 28796 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0744_
timestamp 1676037725
transform 1 0 25024 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0745_
timestamp 1676037725
transform 1 0 27232 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0746_
timestamp 1676037725
transform 1 0 23000 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0747_
timestamp 1676037725
transform 1 0 21988 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0748_
timestamp 1676037725
transform 1 0 23828 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0749_
timestamp 1676037725
transform 1 0 20792 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0750_
timestamp 1676037725
transform 1 0 20700 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0751_
timestamp 1676037725
transform 1 0 16836 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0752_
timestamp 1676037725
transform 1 0 27232 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0753_
timestamp 1676037725
transform 1 0 28704 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0754_
timestamp 1676037725
transform 1 0 41492 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0755_
timestamp 1676037725
transform 1 0 41216 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0756_
timestamp 1676037725
transform 1 0 38272 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0757_
timestamp 1676037725
transform 1 0 38272 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0758_
timestamp 1676037725
transform 1 0 27324 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0759_
timestamp 1676037725
transform 1 0 26312 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0760_
timestamp 1676037725
transform 1 0 27416 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0761_
timestamp 1676037725
transform 1 0 28520 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0762_
timestamp 1676037725
transform 1 0 21988 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0763_
timestamp 1676037725
transform 1 0 20976 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0764_
timestamp 1676037725
transform 1 0 35972 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0765_
timestamp 1676037725
transform 1 0 37444 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0766_
timestamp 1676037725
transform 1 0 24564 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0767_
timestamp 1676037725
transform 1 0 25760 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0768_
timestamp 1676037725
transform 1 0 35604 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0769_
timestamp 1676037725
transform 1 0 34960 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0770_
timestamp 1676037725
transform 1 0 25576 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0771_
timestamp 1676037725
transform 1 0 23644 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0772_
timestamp 1676037725
transform 1 0 38732 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0773_
timestamp 1676037725
transform 1 0 38640 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0774_
timestamp 1676037725
transform 1 0 30636 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0775_
timestamp 1676037725
transform 1 0 29808 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0776_
timestamp 1676037725
transform 1 0 30820 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0777_
timestamp 1676037725
transform 1 0 29716 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0778_
timestamp 1676037725
transform 1 0 34592 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0779_
timestamp 1676037725
transform 1 0 33304 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0780_
timestamp 1676037725
transform 1 0 51244 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _0781_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 45264 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0782_
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0783_
timestamp 1676037725
transform 1 0 23184 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0784_
timestamp 1676037725
transform 1 0 21436 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0785_
timestamp 1676037725
transform 1 0 18768 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0786_
timestamp 1676037725
transform 1 0 20516 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0787_
timestamp 1676037725
transform 1 0 18124 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0788_
timestamp 1676037725
transform 1 0 21160 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0789_
timestamp 1676037725
transform 1 0 18124 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0790_
timestamp 1676037725
transform 1 0 21988 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0791_
timestamp 1676037725
transform 1 0 21620 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0792_
timestamp 1676037725
transform 1 0 27508 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0793_
timestamp 1676037725
transform 1 0 41124 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0794_
timestamp 1676037725
transform 1 0 35328 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0795_
timestamp 1676037725
transform 1 0 25300 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0796_
timestamp 1676037725
transform 1 0 25392 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0797_
timestamp 1676037725
transform 1 0 21988 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0798_
timestamp 1676037725
transform 1 0 34500 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0799_
timestamp 1676037725
transform 1 0 36156 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0800_
timestamp 1676037725
transform 1 0 34868 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0801_
timestamp 1676037725
transform 1 0 33304 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0802_
timestamp 1676037725
transform 1 0 38180 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0803_
timestamp 1676037725
transform 1 0 29716 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0804_
timestamp 1676037725
transform 1 0 40572 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0805_
timestamp 1676037725
transform 1 0 35052 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0806_
timestamp 1676037725
transform 1 0 45816 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0807_
timestamp 1676037725
transform 1 0 47748 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0808_
timestamp 1676037725
transform 1 0 46368 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0809_
timestamp 1676037725
transform 1 0 46092 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0810_
timestamp 1676037725
transform 1 0 20608 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0811_
timestamp 1676037725
transform 1 0 19228 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0812_
timestamp 1676037725
transform 1 0 24564 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0813_
timestamp 1676037725
transform 1 0 23276 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0814_
timestamp 1676037725
transform 1 0 25852 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0815_
timestamp 1676037725
transform 1 0 25576 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0816_
timestamp 1676037725
transform 1 0 23000 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0817_
timestamp 1676037725
transform 1 0 22632 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _0818_
timestamp 1676037725
transform 1 0 44252 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0819_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 46092 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0820_
timestamp 1676037725
transform 1 0 58052 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0821_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27140 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0822_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33212 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _0823_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32844 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _0824_
timestamp 1676037725
transform 1 0 32292 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0825_
timestamp 1676037725
transform 1 0 55660 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0826_
timestamp 1676037725
transform 1 0 55476 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0827_
timestamp 1676037725
transform 1 0 30452 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0828_
timestamp 1676037725
transform 1 0 32752 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0829_
timestamp 1676037725
transform 1 0 35972 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_4  _0830_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35788 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0831_
timestamp 1676037725
transform 1 0 56120 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0832_
timestamp 1676037725
transform 1 0 56948 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0833_
timestamp 1676037725
transform 1 0 33856 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0834_
timestamp 1676037725
transform 1 0 34132 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_4  _0835_
timestamp 1676037725
transform 1 0 35328 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0836_
timestamp 1676037725
transform 1 0 56120 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0837_
timestamp 1676037725
transform 1 0 36432 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0838_
timestamp 1676037725
transform 1 0 52900 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _0839_
timestamp 1676037725
transform 1 0 38272 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0840_
timestamp 1676037725
transform 1 0 37720 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0841_
timestamp 1676037725
transform 1 0 40020 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _0842_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 38640 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0843_
timestamp 1676037725
transform 1 0 57132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _0844_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23276 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0845_
timestamp 1676037725
transform 1 0 31372 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _0846_
timestamp 1676037725
transform 1 0 32292 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _0847_
timestamp 1676037725
transform 1 0 31832 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0848_
timestamp 1676037725
transform 1 0 56120 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _0849_
timestamp 1676037725
transform 1 0 27600 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0850_
timestamp 1676037725
transform 1 0 23000 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0851_
timestamp 1676037725
transform 1 0 30912 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _0852_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31096 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0853_
timestamp 1676037725
transform 1 0 45724 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0854_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 43792 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0855_
timestamp 1676037725
transform 1 0 25668 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0856_
timestamp 1676037725
transform 1 0 50968 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0857_
timestamp 1676037725
transform 1 0 51336 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0858_
timestamp 1676037725
transform 1 0 24564 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0859_
timestamp 1676037725
transform 1 0 53544 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0860_
timestamp 1676037725
transform 1 0 53912 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0861_
timestamp 1676037725
transform 1 0 23828 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0862_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 30268 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0863_
timestamp 1676037725
transform 1 0 22724 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _0864_
timestamp 1676037725
transform 1 0 37904 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0865_
timestamp 1676037725
transform 1 0 37352 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0866_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _0867_
timestamp 1676037725
transform 1 0 38456 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0868_
timestamp 1676037725
transform 1 0 39008 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0869_
timestamp 1676037725
transform 1 0 28244 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0870_
timestamp 1676037725
transform 1 0 27876 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0871_
timestamp 1676037725
transform 1 0 54740 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0872_
timestamp 1676037725
transform 1 0 55752 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0873_
timestamp 1676037725
transform 1 0 29900 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0874_
timestamp 1676037725
transform 1 0 43516 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0875_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 42688 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0876_
timestamp 1676037725
transform 1 0 42688 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0877_
timestamp 1676037725
transform 1 0 30820 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0878_
timestamp 1676037725
transform 1 0 40296 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0879_
timestamp 1676037725
transform 1 0 42596 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0880_
timestamp 1676037725
transform 1 0 41676 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0881_
timestamp 1676037725
transform 1 0 27324 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0882_
timestamp 1676037725
transform 1 0 28060 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0883_
timestamp 1676037725
transform 1 0 53820 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0884_
timestamp 1676037725
transform 1 0 54556 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0885_
timestamp 1676037725
transform 1 0 23460 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_2  _0886_
timestamp 1676037725
transform 1 0 25944 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0887_
timestamp 1676037725
transform 1 0 50416 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0888_
timestamp 1676037725
transform 1 0 51336 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0889_
timestamp 1676037725
transform 1 0 23184 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_2  _0890_
timestamp 1676037725
transform 1 0 24564 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0891_
timestamp 1676037725
transform 1 0 54372 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0892_
timestamp 1676037725
transform 1 0 55476 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0893_
timestamp 1676037725
transform 1 0 37720 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0894_
timestamp 1676037725
transform 1 0 47472 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0895_
timestamp 1676037725
transform 1 0 48024 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_4  _0896_
timestamp 1676037725
transform 1 0 24564 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _0897_
timestamp 1676037725
transform 1 0 55476 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0898_
timestamp 1676037725
transform 1 0 55568 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0899_
timestamp 1676037725
transform 1 0 36800 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0900_
timestamp 1676037725
transform 1 0 50324 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0901_
timestamp 1676037725
transform 1 0 50048 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _0902_
timestamp 1676037725
transform 1 0 24748 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0903_
timestamp 1676037725
transform 1 0 52716 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0904_
timestamp 1676037725
transform 1 0 53728 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0905_
timestamp 1676037725
transform 1 0 40572 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0906_
timestamp 1676037725
transform 1 0 45816 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0907_
timestamp 1676037725
transform 1 0 45172 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0908_
timestamp 1676037725
transform 1 0 32200 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0909_
timestamp 1676037725
transform 1 0 32108 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0910_
timestamp 1676037725
transform 1 0 46000 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0911_
timestamp 1676037725
transform 1 0 46828 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _0912_
timestamp 1676037725
transform 1 0 30176 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0913_
timestamp 1676037725
transform 1 0 50876 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0914_
timestamp 1676037725
transform 1 0 51888 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0915_
timestamp 1676037725
transform 1 0 34868 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0916_
timestamp 1676037725
transform 1 0 32292 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0917_
timestamp 1676037725
transform 1 0 47840 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0918_
timestamp 1676037725
transform 1 0 48300 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _0919_
timestamp 1676037725
transform 1 0 38088 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0920_
timestamp 1676037725
transform 1 0 42228 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0921_
timestamp 1676037725
transform 1 0 43240 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0922_
timestamp 1676037725
transform 1 0 41492 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0923_
timestamp 1676037725
transform 1 0 42780 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a32oi_4  _0924_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32384 0 1 14144
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _0925_
timestamp 1676037725
transform 1 0 31740 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0926_
timestamp 1676037725
transform 1 0 35788 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0927_
timestamp 1676037725
transform 1 0 36248 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0928_
timestamp 1676037725
transform 1 0 16008 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0929_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13156 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0930_
timestamp 1676037725
transform 1 0 13984 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_2  _0931_
timestamp 1676037725
transform 1 0 14536 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0932_
timestamp 1676037725
transform 1 0 14996 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0933_
timestamp 1676037725
transform 1 0 13064 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0934_
timestamp 1676037725
transform 1 0 10488 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0935_
timestamp 1676037725
transform 1 0 10488 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0936_
timestamp 1676037725
transform 1 0 9936 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0937_
timestamp 1676037725
transform 1 0 9384 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and4_4  _0938_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11868 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0939_
timestamp 1676037725
transform 1 0 11684 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0940_
timestamp 1676037725
transform 1 0 10672 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0941_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11684 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0942_
timestamp 1676037725
transform 1 0 19412 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0943_
timestamp 1676037725
transform 1 0 18676 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0944_
timestamp 1676037725
transform 1 0 16836 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0945_
timestamp 1676037725
transform 1 0 14812 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0946_
timestamp 1676037725
transform 1 0 17572 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0947_
timestamp 1676037725
transform 1 0 21252 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0948_
timestamp 1676037725
transform 1 0 18768 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0949_
timestamp 1676037725
transform 1 0 15732 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0950_
timestamp 1676037725
transform 1 0 15824 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and4_2  _0951_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0952_
timestamp 1676037725
transform 1 0 16100 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0953_
timestamp 1676037725
transform 1 0 14628 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0954_
timestamp 1676037725
transform 1 0 18032 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0955_
timestamp 1676037725
transform 1 0 15916 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0956_
timestamp 1676037725
transform 1 0 15272 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0957_
timestamp 1676037725
transform 1 0 16836 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0958_
timestamp 1676037725
transform 1 0 18216 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0959_
timestamp 1676037725
transform 1 0 19412 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0960_
timestamp 1676037725
transform 1 0 19412 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0961_
timestamp 1676037725
transform 1 0 21252 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0962_
timestamp 1676037725
transform 1 0 15916 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0963_
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0964_
timestamp 1676037725
transform 1 0 19596 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0965_
timestamp 1676037725
transform 1 0 15272 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0966_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17388 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and4_2  _0967_
timestamp 1676037725
transform 1 0 19412 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0968_
timestamp 1676037725
transform 1 0 16100 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0969_
timestamp 1676037725
transform 1 0 15180 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0970_
timestamp 1676037725
transform 1 0 10948 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0971_
timestamp 1676037725
transform 1 0 11592 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0972_
timestamp 1676037725
transform 1 0 11776 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and4_2  _0973_
timestamp 1676037725
transform 1 0 12604 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0974_
timestamp 1676037725
transform 1 0 12788 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0975_
timestamp 1676037725
transform 1 0 12880 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0976_
timestamp 1676037725
transform 1 0 9108 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0977_
timestamp 1676037725
transform 1 0 6992 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0978_
timestamp 1676037725
transform 1 0 10120 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0979_
timestamp 1676037725
transform 1 0 9108 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0980_
timestamp 1676037725
transform 1 0 8004 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0981_
timestamp 1676037725
transform 1 0 9108 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0982_
timestamp 1676037725
transform 1 0 6532 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_2  _0983_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 36248 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0984_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19596 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0985_
timestamp 1676037725
transform 1 0 34040 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0986_
timestamp 1676037725
transform 1 0 35512 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0987_
timestamp 1676037725
transform 1 0 38548 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0988_
timestamp 1676037725
transform 1 0 31188 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0989_
timestamp 1676037725
transform 1 0 27048 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0990_
timestamp 1676037725
transform 1 0 19688 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0991_
timestamp 1676037725
transform 1 0 48760 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _0992_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28704 0 -1 10880
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _0993_
timestamp 1676037725
transform 1 0 32292 0 1 3264
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _0994_
timestamp 1676037725
transform 1 0 33212 0 -1 3264
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _0995_
timestamp 1676037725
transform 1 0 37260 0 1 3264
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _0996_
timestamp 1676037725
transform 1 0 28428 0 -1 3264
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _0997_
timestamp 1676037725
transform 1 0 29716 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0998_
timestamp 1676037725
transform 1 0 24748 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0999_
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1000_
timestamp 1676037725
transform 1 0 19688 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1001_
timestamp 1676037725
transform 1 0 21988 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1002_
timestamp 1676037725
transform 1 0 27324 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1003_
timestamp 1676037725
transform 1 0 41124 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1004_
timestamp 1676037725
transform 1 0 38364 0 -1 20672
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1005_
timestamp 1676037725
transform 1 0 27140 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1006_
timestamp 1676037725
transform 1 0 27508 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1007_
timestamp 1676037725
transform 1 0 21988 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1008_
timestamp 1676037725
transform 1 0 35788 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1009_
timestamp 1676037725
transform 1 0 22356 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1010_
timestamp 1676037725
transform 1 0 35144 0 -1 20672
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1011_
timestamp 1676037725
transform 1 0 24564 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1012_
timestamp 1676037725
transform 1 0 38732 0 -1 18496
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1013_
timestamp 1676037725
transform 1 0 30268 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1014_
timestamp 1676037725
transform 1 0 30268 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1015_
timestamp 1676037725
transform 1 0 32476 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1016_
timestamp 1676037725
transform 1 0 56856 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1017_
timestamp 1676037725
transform 1 0 27324 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1018_
timestamp 1676037725
transform 1 0 22632 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1019_
timestamp 1676037725
transform 1 0 19596 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1020_
timestamp 1676037725
transform 1 0 19596 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1021_
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1022_
timestamp 1676037725
transform 1 0 19596 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1023_
timestamp 1676037725
transform 1 0 20056 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1024_
timestamp 1676037725
transform 1 0 19412 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1025_
timestamp 1676037725
transform 1 0 19780 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1026_
timestamp 1676037725
transform 1 0 19780 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1027_
timestamp 1676037725
transform 1 0 25668 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1028_
timestamp 1676037725
transform 1 0 40572 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1029_
timestamp 1676037725
transform 1 0 34684 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1030_
timestamp 1676037725
transform 1 0 26128 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1031_
timestamp 1676037725
transform 1 0 24748 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1032_
timestamp 1676037725
transform 1 0 19412 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1033_
timestamp 1676037725
transform 1 0 33856 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1034_
timestamp 1676037725
transform 1 0 36340 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1035_
timestamp 1676037725
transform 1 0 34408 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1036_
timestamp 1676037725
transform 1 0 32936 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1037_
timestamp 1676037725
transform 1 0 37352 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1038_
timestamp 1676037725
transform 1 0 28428 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1039_
timestamp 1676037725
transform 1 0 40296 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1040_
timestamp 1676037725
transform 1 0 33672 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1041_
timestamp 1676037725
transform 1 0 44988 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1042_
timestamp 1676037725
transform 1 0 46736 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1043_
timestamp 1676037725
transform 1 0 45172 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1044_
timestamp 1676037725
transform 1 0 45448 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1045_
timestamp 1676037725
transform 1 0 19412 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1046_
timestamp 1676037725
transform 1 0 23276 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1047_
timestamp 1676037725
transform 1 0 24656 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1048_
timestamp 1676037725
transform 1 0 22448 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1049_
timestamp 1676037725
transform 1 0 56856 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1050_
timestamp 1676037725
transform 1 0 56856 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1051_
timestamp 1676037725
transform 1 0 56856 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1052_
timestamp 1676037725
transform 1 0 39100 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1053_
timestamp 1676037725
transform 1 0 56856 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1054_
timestamp 1676037725
transform 1 0 45172 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1055_
timestamp 1676037725
transform 1 0 50968 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1056_
timestamp 1676037725
transform 1 0 53544 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1057_
timestamp 1676037725
transform 1 0 37996 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1058_
timestamp 1676037725
transform 1 0 40020 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1059_
timestamp 1676037725
transform 1 0 56856 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1060_
timestamp 1676037725
transform 1 0 42688 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1061_
timestamp 1676037725
transform 1 0 43056 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1062_
timestamp 1676037725
transform 1 0 54924 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1063_
timestamp 1676037725
transform 1 0 51428 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1064_
timestamp 1676037725
transform 1 0 55752 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1065_
timestamp 1676037725
transform 1 0 48116 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1066_
timestamp 1676037725
transform 1 0 56580 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1067_
timestamp 1676037725
transform 1 0 50232 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1068_
timestamp 1676037725
transform 1 0 53084 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1069_
timestamp 1676037725
transform 1 0 45356 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1070_
timestamp 1676037725
transform 1 0 46092 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1071_
timestamp 1676037725
transform 1 0 51428 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1072_
timestamp 1676037725
transform 1 0 48484 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1073_
timestamp 1676037725
transform 1 0 42964 0 1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1074_
timestamp 1676037725
transform 1 0 43056 0 -1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1075_
timestamp 1676037725
transform 1 0 32292 0 -1 15232
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1076_
timestamp 1676037725
transform 1 0 36340 0 1 11968
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1077_
timestamp 1676037725
transform 1 0 14260 0 1 15232
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1078_
timestamp 1676037725
transform 1 0 14260 0 1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1079_
timestamp 1676037725
transform 1 0 14260 0 1 13056
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1080_
timestamp 1676037725
transform 1 0 9292 0 1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1081_
timestamp 1676037725
transform 1 0 9292 0 1 13056
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1082_
timestamp 1676037725
transform 1 0 11684 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1083_
timestamp 1676037725
transform 1 0 11040 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1084_
timestamp 1676037725
transform 1 0 16836 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1085_
timestamp 1676037725
transform 1 0 16836 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1086_
timestamp 1676037725
transform 1 0 14720 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1087_
timestamp 1676037725
transform 1 0 16836 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1088_
timestamp 1676037725
transform 1 0 14628 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1089_
timestamp 1676037725
transform 1 0 16836 0 -1 19584
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1090_
timestamp 1676037725
transform 1 0 19412 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1091_
timestamp 1676037725
transform 1 0 17112 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1092_
timestamp 1676037725
transform 1 0 16928 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1093_
timestamp 1676037725
transform 1 0 14444 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1094_
timestamp 1676037725
transform 1 0 13156 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1095_
timestamp 1676037725
transform 1 0 11868 0 -1 19584
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1096_
timestamp 1676037725
transform 1 0 12144 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1097_
timestamp 1676037725
transform 1 0 8188 0 -1 17408
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1098_
timestamp 1676037725
transform 1 0 9108 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1099_
timestamp 1676037725
transform 1 0 6808 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1100_
timestamp 1676037725
transform 1 0 6532 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_2  _1121_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29716 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1122_
timestamp 1676037725
transform 1 0 28888 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1123_
timestamp 1676037725
transform 1 0 30636 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1124_
timestamp 1676037725
transform 1 0 31464 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1125_
timestamp 1676037725
transform 1 0 32752 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1126_
timestamp 1676037725
transform 1 0 33488 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1127_
timestamp 1676037725
transform 1 0 34224 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1128_
timestamp 1676037725
transform 1 0 34040 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1129_
timestamp 1676037725
transform 1 0 33304 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1130_
timestamp 1676037725
transform 1 0 34868 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1131_
timestamp 1676037725
transform 1 0 33764 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1132_
timestamp 1676037725
transform 1 0 37444 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1133_
timestamp 1676037725
transform 1 0 36340 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 38732 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_wb_clk_i
timestamp 1676037725
transform 1 0 23368 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_wb_clk_i
timestamp 1676037725
transform 1 0 28612 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_wb_clk_i
timestamp 1676037725
transform 1 0 26036 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_wb_clk_i
timestamp 1676037725
transform 1 0 28612 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_wb_clk_i
timestamp 1676037725
transform 1 0 44160 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_wb_clk_i
timestamp 1676037725
transform 1 0 46828 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_wb_clk_i
timestamp 1676037725
transform 1 0 44160 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_wb_clk_i
timestamp 1676037725
transform 1 0 46828 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_4  fanout411 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 55476 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout412 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 54556 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout413 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 30912 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout414
timestamp 1676037725
transform 1 0 30176 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout415
timestamp 1676037725
transform 1 0 45172 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout416
timestamp 1676037725
transform 1 0 44160 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout417
timestamp 1676037725
transform 1 0 47748 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout418
timestamp 1676037725
transform 1 0 52164 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout419
timestamp 1676037725
transform 1 0 47012 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout420 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28428 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout421
timestamp 1676037725
transform 1 0 33764 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout422
timestamp 1676037725
transform 1 0 46184 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout423
timestamp 1676037725
transform 1 0 46368 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout424
timestamp 1676037725
transform 1 0 29808 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout425
timestamp 1676037725
transform 1 0 30728 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout426
timestamp 1676037725
transform 1 0 38180 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout427 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33304 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout429
timestamp 1676037725
transform 1 0 14260 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout430
timestamp 1676037725
transform 1 0 37444 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  fanout431 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  fanout432
timestamp 1676037725
transform 1 0 22632 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  fanout433
timestamp 1676037725
transform 1 0 24564 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout434
timestamp 1676037725
transform 1 0 20700 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout435
timestamp 1676037725
transform 1 0 17940 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout436
timestamp 1676037725
transform 1 0 36064 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout437
timestamp 1676037725
transform 1 0 28428 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout438
timestamp 1676037725
transform 1 0 28152 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout439
timestamp 1676037725
transform 1 0 28244 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout440
timestamp 1676037725
transform 1 0 30820 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  fanout441
timestamp 1676037725
transform 1 0 15732 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_6  fanout442
timestamp 1676037725
transform 1 0 12144 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout443
timestamp 1676037725
transform 1 0 19504 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout444
timestamp 1676037725
transform 1 0 28336 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout445
timestamp 1676037725
transform 1 0 29440 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout446
timestamp 1676037725
transform 1 0 24564 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_12  fanout447
timestamp 1676037725
transform 1 0 27508 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  fanout448
timestamp 1676037725
transform 1 0 21988 0 -1 59840
box -38 -48 866 592
use sky130_fd_sc_hd__buf_12  fanout449
timestamp 1676037725
transform 1 0 10672 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  fanout450
timestamp 1676037725
transform 1 0 27140 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  fanout451
timestamp 1676037725
transform 1 0 25576 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_4  fanout452
timestamp 1676037725
transform 1 0 12972 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout453
timestamp 1676037725
transform 1 0 35604 0 -1 57664
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout454
timestamp 1676037725
transform 1 0 24564 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  fanout455
timestamp 1676037725
transform 1 0 19412 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_8  fanout456
timestamp 1676037725
transform 1 0 29900 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout457
timestamp 1676037725
transform 1 0 19412 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout458
timestamp 1676037725
transform 1 0 18860 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout459
timestamp 1676037725
transform 1 0 22356 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_8  fanout460 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16560 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout461
timestamp 1676037725
transform 1 0 17020 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout462
timestamp 1676037725
transform 1 0 25116 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  fanout463
timestamp 1676037725
transform 1 0 17940 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout464
timestamp 1676037725
transform 1 0 24564 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_8  fanout465
timestamp 1676037725
transform 1 0 17480 0 -1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout466
timestamp 1676037725
transform 1 0 21436 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout467
timestamp 1676037725
transform 1 0 9476 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout468
timestamp 1676037725
transform 1 0 9568 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout469
timestamp 1676037725
transform 1 0 11684 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout470
timestamp 1676037725
transform 1 0 13984 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout471
timestamp 1676037725
transform 1 0 13432 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout472
timestamp 1676037725
transform 1 0 14168 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout473
timestamp 1676037725
transform 1 0 22356 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_8  fanout474
timestamp 1676037725
transform 1 0 29992 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  fanout475
timestamp 1676037725
transform 1 0 35420 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout476
timestamp 1676037725
transform 1 0 31372 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout477
timestamp 1676037725
transform 1 0 33764 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout478
timestamp 1676037725
transform 1 0 43700 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout479
timestamp 1676037725
transform 1 0 26128 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout480
timestamp 1676037725
transform 1 0 34500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout481
timestamp 1676037725
transform 1 0 29072 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout482
timestamp 1676037725
transform 1 0 34868 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout483
timestamp 1676037725
transform 1 0 42872 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout484
timestamp 1676037725
transform 1 0 37076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout485
timestamp 1676037725
transform 1 0 45172 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout486
timestamp 1676037725
transform 1 0 45908 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout487
timestamp 1676037725
transform 1 0 45264 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout488
timestamp 1676037725
transform 1 0 42780 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout489
timestamp 1676037725
transform 1 0 43700 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout490
timestamp 1676037725
transform 1 0 56396 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__bufbuf_16  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19136 0 -1 18496
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold2
timestamp 1676037725
transform 1 0 6256 0 1 18496
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold3
timestamp 1676037725
transform 1 0 21252 0 1 18496
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold4
timestamp 1676037725
transform 1 0 10120 0 1 17408
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold5
timestamp 1676037725
transform 1 0 28612 0 -1 21760
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold6
timestamp 1676037725
transform 1 0 16560 0 1 20672
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold7
timestamp 1676037725
transform 1 0 24288 0 -1 20672
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold8
timestamp 1676037725
transform 1 0 11408 0 1 18496
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold9
timestamp 1676037725
transform 1 0 24288 0 -1 18496
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold10
timestamp 1676037725
transform 1 0 8556 0 -1 18496
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold11
timestamp 1676037725
transform 1 0 21988 0 -1 13056
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold12
timestamp 1676037725
transform 1 0 13708 0 -1 14144
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold13
timestamp 1676037725
transform 1 0 19136 0 -1 14144
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold14
timestamp 1676037725
transform 1 0 16560 0 1 14144
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold15
timestamp 1676037725
transform 1 0 19872 0 1 8704
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold16
timestamp 1676037725
transform 1 0 8832 0 -1 15232
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold17
timestamp 1676037725
transform 1 0 16560 0 1 15232
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold18
timestamp 1676037725
transform 1 0 12236 0 -1 15232
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold19
timestamp 1676037725
transform 1 0 24288 0 -1 7616
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold20
timestamp 1676037725
transform 1 0 13984 0 -1 13056
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold21
timestamp 1676037725
transform 1 0 17664 0 -1 17408
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold22
timestamp 1676037725
transform 1 0 12788 0 -1 18496
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold23
timestamp 1676037725
transform 1 0 29440 0 -1 20672
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold24
timestamp 1676037725
transform 1 0 16560 0 1 21760
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold25
timestamp 1676037725
transform 1 0 13984 0 -1 20672
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold26
timestamp 1676037725
transform 1 0 26312 0 1 19584
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold27
timestamp 1676037725
transform 1 0 16100 0 1 17408
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold28
timestamp 1676037725
transform 1 0 13984 0 -1 19584
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold29
timestamp 1676037725
transform 1 0 23828 0 -1 16320
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold30
timestamp 1676037725
transform 1 0 21988 0 -1 17408
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold31
timestamp 1676037725
transform 1 0 16560 0 1 16320
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold32
timestamp 1676037725
transform 1 0 24288 0 -1 19584
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold33
timestamp 1676037725
transform 1 0 19964 0 1 16320
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold34
timestamp 1676037725
transform 1 0 18492 0 -1 16320
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold35
timestamp 1676037725
transform 1 0 20884 0 1 20672
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold36
timestamp 1676037725
transform 1 0 16560 0 1 18496
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold37
timestamp 1676037725
transform 1 0 23552 0 -1 21760
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold38
timestamp 1676037725
transform 1 0 18768 0 -1 21760
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold39
timestamp 1676037725
transform 1 0 16560 0 1 19584
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold40
timestamp 1676037725
transform 1 0 21620 0 1 14144
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold41
timestamp 1676037725
transform 1 0 11408 0 1 13056
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold42
timestamp 1676037725
transform 1 0 11408 0 1 14144
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold43
timestamp 1676037725
transform 1 0 20056 0 1 17408
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold44
timestamp 1676037725
transform 1 0 8004 0 -1 20672
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold45
timestamp 1676037725
transform 1 0 6256 0 1 19584
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold46
timestamp 1676037725
transform 1 0 20056 0 1 11968
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold47
timestamp 1676037725
transform 1 0 17756 0 -1 13056
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold48
timestamp 1676037725
transform 1 0 16560 0 1 13056
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold49
timestamp 1676037725
transform 1 0 24932 0 1 7616
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold50
timestamp 1676037725
transform 1 0 15916 0 1 11968
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold51
timestamp 1676037725
transform 1 0 24104 0 -1 8704
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold52
timestamp 1676037725
transform 1 0 8832 0 -1 14144
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold53
timestamp 1676037725
transform 1 0 9844 0 1 15232
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold54
timestamp 1676037725
transform 1 0 21068 0 1 15232
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold55
timestamp 1676037725
transform 1 0 18952 0 -1 15232
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold56
timestamp 1676037725
transform 1 0 18492 0 -1 20672
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold57
timestamp 1676037725
transform 1 0 11408 0 1 19584
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold58
timestamp 1676037725
transform 1 0 26496 0 1 18496
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold59
timestamp 1676037725
transform 1 0 27140 0 -1 19584
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold60
timestamp 1676037725
transform 1 0 8832 0 -1 19584
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold61
timestamp 1676037725
transform 1 0 34868 0 1 20672
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold62
timestamp 1676037725
transform 1 0 30636 0 1 19584
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold63
timestamp 1676037725
transform 1 0 12512 0 -1 17408
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold64
timestamp 1676037725
transform 1 0 26036 0 1 10880
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold65
timestamp 1676037725
transform 1 0 20976 0 1 13056
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold66
timestamp 1676037725
transform 1 0 32108 0 -1 18496
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold67
timestamp 1676037725
transform 1 0 21988 0 -1 15232
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold68
timestamp 1676037725
transform 1 0 29072 0 -1 6528
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold69
timestamp 1676037725
transform 1 0 24932 0 1 5440
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold70
timestamp 1676037725
transform 1 0 19136 0 -1 19584
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold71
timestamp 1676037725
transform 1 0 21528 0 1 19584
box -38 -48 2430 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1676037725
transform 1 0 41768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp 1676037725
transform 1 0 40940 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1676037725
transform 1 0 41032 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1676037725
transform 1 0 44988 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1676037725
transform 1 0 41768 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1676037725
transform 1 0 41308 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input7
timestamp 1676037725
transform 1 0 41584 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1676037725
transform 1 0 42596 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1676037725
transform 1 0 44344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1676037725
transform 1 0 46920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1676037725
transform 1 0 45172 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1676037725
transform 1 0 41216 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1676037725
transform 1 0 43332 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1676037725
transform 1 0 45908 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1676037725
transform 1 0 45080 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1676037725
transform 1 0 44068 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1676037725
transform 1 0 45816 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1676037725
transform 1 0 45172 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1676037725
transform 1 0 44804 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1676037725
transform 1 0 43792 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1676037725
transform 1 0 40756 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input22
timestamp 1676037725
transform 1 0 40296 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input23
timestamp 1676037725
transform 1 0 44252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input24
timestamp 1676037725
transform 1 0 45172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input25
timestamp 1676037725
transform 1 0 40020 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input26
timestamp 1676037725
transform 1 0 39928 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1676037725
transform 1 0 40020 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input28
timestamp 1676037725
transform 1 0 54096 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input29
timestamp 1676037725
transform 1 0 54648 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input30
timestamp 1676037725
transform 1 0 55476 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input31
timestamp 1676037725
transform 1 0 56396 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input32
timestamp 1676037725
transform 1 0 56856 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1676037725
transform 1 0 58052 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input34
timestamp 1676037725
transform 1 0 57868 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input35
timestamp 1676037725
transform 1 0 57132 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1676037725
transform 1 0 46552 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input37
timestamp 1676037725
transform 1 0 48484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1676037725
transform 1 0 50324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1676037725
transform 1 0 48208 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input40
timestamp 1676037725
transform 1 0 48668 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input41
timestamp 1676037725
transform 1 0 49220 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input42
timestamp 1676037725
transform 1 0 49588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1676037725
transform 1 0 51060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1676037725
transform 1 0 50508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1676037725
transform 1 0 50324 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1676037725
transform 1 0 51796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1676037725
transform 1 0 45908 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1676037725
transform 1 0 51244 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1676037725
transform 1 0 51060 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1676037725
transform 1 0 51980 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1676037725
transform 1 0 51796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1676037725
transform 1 0 52900 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input53
timestamp 1676037725
transform 1 0 52532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 1676037725
transform 1 0 52072 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1676037725
transform 1 0 47748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input56
timestamp 1676037725
transform 1 0 45724 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input57
timestamp 1676037725
transform 1 0 46000 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input58
timestamp 1676037725
transform 1 0 46276 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input59
timestamp 1676037725
transform 1 0 47748 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input60
timestamp 1676037725
transform 1 0 46828 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input61
timestamp 1676037725
transform 1 0 47748 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input62
timestamp 1676037725
transform 1 0 48668 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1676037725
transform 1 0 13432 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1676037725
transform 1 0 20424 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1676037725
transform 1 0 21160 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input66
timestamp 1676037725
transform 1 0 22264 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input67
timestamp 1676037725
transform 1 0 23184 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1676037725
transform 1 0 23736 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1676037725
transform 1 0 24472 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input70
timestamp 1676037725
transform 1 0 25208 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input71
timestamp 1676037725
transform 1 0 26128 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input72
timestamp 1676037725
transform 1 0 27140 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 1676037725
transform 1 0 27416 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1676037725
transform 1 0 14168 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input75
timestamp 1676037725
transform 1 0 28152 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input76
timestamp 1676037725
transform 1 0 28888 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input77
timestamp 1676037725
transform 1 0 29716 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input78
timestamp 1676037725
transform 1 0 30360 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input79
timestamp 1676037725
transform 1 0 31096 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input80
timestamp 1676037725
transform 1 0 32292 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input81
timestamp 1676037725
transform 1 0 33212 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input82
timestamp 1676037725
transform 1 0 14904 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input83
timestamp 1676037725
transform 1 0 15640 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input84
timestamp 1676037725
transform 1 0 16008 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input85
timestamp 1676037725
transform 1 0 17112 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input86
timestamp 1676037725
transform 1 0 17848 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input87
timestamp 1676037725
transform 1 0 18584 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input88
timestamp 1676037725
transform 1 0 19320 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input89
timestamp 1676037725
transform 1 0 19688 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input90
timestamp 1676037725
transform 1 0 1564 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input91
timestamp 1676037725
transform 1 0 1564 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input92
timestamp 1676037725
transform 1 0 1564 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input93
timestamp 1676037725
transform 1 0 1564 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input94
timestamp 1676037725
transform 1 0 1564 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input95
timestamp 1676037725
transform 1 0 1564 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input96
timestamp 1676037725
transform 1 0 1564 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input97
timestamp 1676037725
transform 1 0 1564 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input98
timestamp 1676037725
transform 1 0 1564 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input99
timestamp 1676037725
transform 1 0 1564 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input100
timestamp 1676037725
transform 1 0 1564 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input101
timestamp 1676037725
transform 1 0 1564 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input102
timestamp 1676037725
transform 1 0 1564 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input103
timestamp 1676037725
transform 1 0 1564 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input104
timestamp 1676037725
transform 1 0 1564 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input105
timestamp 1676037725
transform 1 0 1564 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input106
timestamp 1676037725
transform 1 0 1564 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input107
timestamp 1676037725
transform 1 0 1564 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input108
timestamp 1676037725
transform 1 0 1564 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input109
timestamp 1676037725
transform 1 0 2760 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input110
timestamp 1676037725
transform 1 0 1564 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input111
timestamp 1676037725
transform 1 0 1564 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input112
timestamp 1676037725
transform 1 0 1564 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input113
timestamp 1676037725
transform 1 0 1564 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input114
timestamp 1676037725
transform 1 0 1564 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input115
timestamp 1676037725
transform 1 0 1564 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input116
timestamp 1676037725
transform 1 0 1564 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input117
timestamp 1676037725
transform 1 0 1564 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input118
timestamp 1676037725
transform 1 0 33948 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input119
timestamp 1676037725
transform 1 0 41492 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input120
timestamp 1676037725
transform 1 0 41400 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input121
timestamp 1676037725
transform 1 0 42596 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input122
timestamp 1676037725
transform 1 0 43516 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input123
timestamp 1676037725
transform 1 0 44252 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input124
timestamp 1676037725
transform 1 0 45172 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input125
timestamp 1676037725
transform 1 0 45908 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input126
timestamp 1676037725
transform 1 0 46644 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input127
timestamp 1676037725
transform 1 0 46552 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input128
timestamp 1676037725
transform 1 0 47748 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input129
timestamp 1676037725
transform 1 0 34868 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input130
timestamp 1676037725
transform 1 0 48484 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input131
timestamp 1676037725
transform 1 0 49220 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input132
timestamp 1676037725
transform 1 0 50324 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input133
timestamp 1676037725
transform 1 0 50232 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input134
timestamp 1676037725
transform 1 0 51244 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input135
timestamp 1676037725
transform 1 0 51980 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input136
timestamp 1676037725
transform 1 0 52900 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input137
timestamp 1676037725
transform 1 0 35604 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input138
timestamp 1676037725
transform 1 0 36340 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input139
timestamp 1676037725
transform 1 0 36248 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input140
timestamp 1676037725
transform 1 0 37444 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input141
timestamp 1676037725
transform 1 0 38180 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input142
timestamp 1676037725
transform 1 0 38916 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input143
timestamp 1676037725
transform 1 0 40020 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input144
timestamp 1676037725
transform 1 0 40756 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input145
timestamp 1676037725
transform 1 0 58052 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input146
timestamp 1676037725
transform 1 0 56120 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input147
timestamp 1676037725
transform 1 0 57224 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input148
timestamp 1676037725
transform 1 0 57868 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input149
timestamp 1676037725
transform 1 0 57868 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input150
timestamp 1676037725
transform 1 0 57868 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input151
timestamp 1676037725
transform 1 0 58052 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input152
timestamp 1676037725
transform 1 0 58052 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input153
timestamp 1676037725
transform 1 0 58052 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input154
timestamp 1676037725
transform 1 0 57132 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input155
timestamp 1676037725
transform 1 0 56396 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input156
timestamp 1676037725
transform 1 0 55384 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input157
timestamp 1676037725
transform 1 0 6624 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input158
timestamp 1676037725
transform 1 0 7544 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input159
timestamp 1676037725
transform 1 0 8280 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input160
timestamp 1676037725
transform 1 0 9016 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input161
timestamp 1676037725
transform 1 0 9384 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input162
timestamp 1676037725
transform 1 0 10120 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input163
timestamp 1676037725
transform 1 0 10856 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input164
timestamp 1676037725
transform 1 0 11960 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input165
timestamp 1676037725
transform 1 0 1564 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input166
timestamp 1676037725
transform 1 0 1564 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input167
timestamp 1676037725
transform 1 0 1564 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input168
timestamp 1676037725
transform 1 0 1564 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input169
timestamp 1676037725
transform 1 0 1564 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input170
timestamp 1676037725
transform 1 0 1564 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input171
timestamp 1676037725
transform 1 0 1564 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input172
timestamp 1676037725
transform 1 0 1564 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input173
timestamp 1676037725
transform 1 0 1564 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input174
timestamp 1676037725
transform 1 0 1564 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input175
timestamp 1676037725
transform 1 0 2484 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input176
timestamp 1676037725
transform 1 0 2484 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input177
timestamp 1676037725
transform 1 0 3128 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input178
timestamp 1676037725
transform 1 0 3864 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input179
timestamp 1676037725
transform 1 0 4232 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input180
timestamp 1676037725
transform 1 0 4968 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input181
timestamp 1676037725
transform 1 0 5704 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input182
timestamp 1676037725
transform 1 0 40848 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input183
timestamp 1676037725
transform 1 0 40480 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input184
timestamp 1676037725
transform 1 0 37444 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input185
timestamp 1676037725
transform 1 0 40020 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input186
timestamp 1676037725
transform 1 0 1564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input187
timestamp 1676037725
transform 1 0 1564 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input188
timestamp 1676037725
transform 1 0 1564 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input189
timestamp 1676037725
transform 1 0 1564 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input190
timestamp 1676037725
transform 1 0 1564 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input191
timestamp 1676037725
transform 1 0 1564 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input192
timestamp 1676037725
transform 1 0 1564 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input193
timestamp 1676037725
transform 1 0 1564 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input194
timestamp 1676037725
transform 1 0 52900 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input195
timestamp 1676037725
transform 1 0 52900 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input196
timestamp 1676037725
transform 1 0 54004 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input197
timestamp 1676037725
transform 1 0 53636 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input198
timestamp 1676037725
transform 1 0 53820 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input199
timestamp 1676037725
transform 1 0 54004 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input200
timestamp 1676037725
transform 1 0 54924 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input201
timestamp 1676037725
transform 1 0 54556 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input202
timestamp 1676037725
transform 1 0 55476 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input203
timestamp 1676037725
transform 1 0 55476 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input204
timestamp 1676037725
transform 1 0 55844 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input205
timestamp 1676037725
transform 1 0 3128 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input206
timestamp 1676037725
transform 1 0 6532 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input207
timestamp 1676037725
transform 1 0 4968 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input208
timestamp 1676037725
transform 1 0 4232 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input209
timestamp 1676037725
transform 1 0 8188 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input210
timestamp 1676037725
transform 1 0 7544 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input211
timestamp 1676037725
transform 1 0 6440 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input212
timestamp 1676037725
transform 1 0 7268 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input213
timestamp 1676037725
transform 1 0 5704 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input214
timestamp 1676037725
transform 1 0 4968 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input215
timestamp 1676037725
transform 1 0 8280 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input216
timestamp 1676037725
transform 1 0 5704 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input217
timestamp 1676037725
transform 1 0 6992 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input218
timestamp 1676037725
transform 1 0 6808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input219
timestamp 1676037725
transform 1 0 7728 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input220
timestamp 1676037725
transform 1 0 7544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input221
timestamp 1676037725
transform 1 0 8280 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input222
timestamp 1676037725
transform 1 0 10856 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input223
timestamp 1676037725
transform 1 0 12052 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input224
timestamp 1676037725
transform 1 0 11776 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input225
timestamp 1676037725
transform 1 0 11684 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input226
timestamp 1676037725
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input227
timestamp 1676037725
transform 1 0 12512 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input228
timestamp 1676037725
transform 1 0 11592 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input229
timestamp 1676037725
transform 1 0 10120 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input230
timestamp 1676037725
transform 1 0 10856 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input231
timestamp 1676037725
transform 1 0 12052 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input232
timestamp 1676037725
transform 1 0 12788 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input233
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input234
timestamp 1676037725
transform 1 0 4232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input235
timestamp 1676037725
transform 1 0 4968 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input236
timestamp 1676037725
transform 1 0 5704 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input237
timestamp 1676037725
transform 1 0 6808 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input238
timestamp 1676037725
transform 1 0 5704 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input239
timestamp 1676037725
transform 1 0 39560 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input240
timestamp 1676037725
transform 1 0 53268 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input241
timestamp 1676037725
transform 1 0 12696 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  input242
timestamp 1676037725
transform 1 0 1564 0 1 60928
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  input243
timestamp 1676037725
transform 1 0 53176 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input244
timestamp 1676037725
transform 1 0 1564 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input245
timestamp 1676037725
transform 1 0 58052 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input246
timestamp 1676037725
transform 1 0 57868 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input247
timestamp 1676037725
transform 1 0 56948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input248
timestamp 1676037725
transform 1 0 57868 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input249
timestamp 1676037725
transform 1 0 58052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input250
timestamp 1676037725
transform 1 0 58052 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input251
timestamp 1676037725
transform 1 0 58052 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input252
timestamp 1676037725
transform 1 0 58052 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input253
timestamp 1676037725
transform 1 0 58052 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input254
timestamp 1676037725
transform 1 0 58052 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input255
timestamp 1676037725
transform 1 0 57868 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input256
timestamp 1676037725
transform 1 0 56948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input257
timestamp 1676037725
transform 1 0 58052 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input258
timestamp 1676037725
transform 1 0 56948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input259
timestamp 1676037725
transform 1 0 58052 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input260
timestamp 1676037725
transform 1 0 57868 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input261
timestamp 1676037725
transform 1 0 57040 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input262
timestamp 1676037725
transform 1 0 58052 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input263
timestamp 1676037725
transform 1 0 56948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input264
timestamp 1676037725
transform 1 0 57868 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input265
timestamp 1676037725
transform 1 0 56948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input266
timestamp 1676037725
transform 1 0 57868 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input267
timestamp 1676037725
transform 1 0 58052 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input268
timestamp 1676037725
transform 1 0 58052 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input269
timestamp 1676037725
transform 1 0 57868 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input270
timestamp 1676037725
transform 1 0 56120 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input271
timestamp 1676037725
transform 1 0 56948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input272
timestamp 1676037725
transform 1 0 57040 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input273
timestamp 1676037725
transform 1 0 56948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input274
timestamp 1676037725
transform 1 0 57868 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input275
timestamp 1676037725
transform 1 0 56948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input276
timestamp 1676037725
transform 1 0 57868 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input277
timestamp 1676037725
transform 1 0 57868 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input278
timestamp 1676037725
transform 1 0 58052 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input279
timestamp 1676037725
transform 1 0 58052 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  max_cap428
timestamp 1676037725
transform 1 0 23000 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  multiplexer_491 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23828 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_492
timestamp 1676037725
transform 1 0 22356 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_493
timestamp 1676037725
transform 1 0 24472 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_494
timestamp 1676037725
transform 1 0 27692 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_495
timestamp 1676037725
transform 1 0 15916 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_496
timestamp 1676037725
transform 1 0 16100 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_497
timestamp 1676037725
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_498
timestamp 1676037725
transform 1 0 16836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_499
timestamp 1676037725
transform 1 0 14260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_500
timestamp 1676037725
transform 1 0 16836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_501
timestamp 1676037725
transform 1 0 58144 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_502
timestamp 1676037725
transform 1 0 58144 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_503
timestamp 1676037725
transform 1 0 58144 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_504
timestamp 1676037725
transform 1 0 58144 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_505
timestamp 1676037725
transform 1 0 27140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_506
timestamp 1676037725
transform 1 0 21988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_507
timestamp 1676037725
transform 1 0 24564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_508
timestamp 1676037725
transform 1 0 26404 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_509
timestamp 1676037725
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_510
timestamp 1676037725
transform 1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output280
timestamp 1676037725
transform 1 0 1564 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  output281
timestamp 1676037725
transform 1 0 1564 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output282
timestamp 1676037725
transform 1 0 1564 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output283
timestamp 1676037725
transform 1 0 1564 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output284
timestamp 1676037725
transform 1 0 1564 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output285
timestamp 1676037725
transform 1 0 1564 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output286
timestamp 1676037725
transform 1 0 1564 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output287
timestamp 1676037725
transform 1 0 1564 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output288
timestamp 1676037725
transform 1 0 1564 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output289
timestamp 1676037725
transform 1 0 1564 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output290
timestamp 1676037725
transform 1 0 1564 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output291
timestamp 1676037725
transform 1 0 1564 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output292
timestamp 1676037725
transform 1 0 1564 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output293
timestamp 1676037725
transform 1 0 1564 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output294
timestamp 1676037725
transform 1 0 1564 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output295
timestamp 1676037725
transform 1 0 1564 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output296
timestamp 1676037725
transform 1 0 1564 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output297
timestamp 1676037725
transform 1 0 1564 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output298
timestamp 1676037725
transform 1 0 1564 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output299
timestamp 1676037725
transform 1 0 1564 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output300
timestamp 1676037725
transform 1 0 1564 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output301
timestamp 1676037725
transform 1 0 1564 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output302
timestamp 1676037725
transform 1 0 1564 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output303
timestamp 1676037725
transform 1 0 1564 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output304
timestamp 1676037725
transform 1 0 1564 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output305
timestamp 1676037725
transform 1 0 1564 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output306
timestamp 1676037725
transform 1 0 1564 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output307
timestamp 1676037725
transform 1 0 1564 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output308
timestamp 1676037725
transform 1 0 1564 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output309
timestamp 1676037725
transform 1 0 25208 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output310
timestamp 1676037725
transform 1 0 26128 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output311
timestamp 1676037725
transform 1 0 26128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output312
timestamp 1676037725
transform 1 0 27508 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output313
timestamp 1676037725
transform 1 0 27784 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output314
timestamp 1676037725
transform 1 0 29716 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output315
timestamp 1676037725
transform 1 0 28704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output316
timestamp 1676037725
transform 1 0 30268 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output317
timestamp 1676037725
transform 1 0 30176 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output318
timestamp 1676037725
transform 1 0 30820 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output319
timestamp 1676037725
transform 1 0 31096 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output320
timestamp 1676037725
transform 1 0 32292 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output321
timestamp 1676037725
transform 1 0 32292 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output322
timestamp 1676037725
transform 1 0 33212 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output323
timestamp 1676037725
transform 1 0 34868 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output324
timestamp 1676037725
transform 1 0 35788 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output325
timestamp 1676037725
transform 1 0 33488 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output326
timestamp 1676037725
transform 1 0 35328 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output327
timestamp 1676037725
transform 1 0 34868 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output328
timestamp 1676037725
transform 1 0 34408 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output329
timestamp 1676037725
transform 1 0 37444 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output330
timestamp 1676037725
transform 1 0 35328 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output331
timestamp 1676037725
transform 1 0 38364 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output332
timestamp 1676037725
transform 1 0 36248 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output333
timestamp 1676037725
transform 1 0 34960 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output334
timestamp 1676037725
transform 1 0 35880 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output335
timestamp 1676037725
transform 1 0 39008 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output336
timestamp 1676037725
transform 1 0 37444 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output337
timestamp 1676037725
transform 1 0 12328 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output338
timestamp 1676037725
transform 1 0 14444 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output339
timestamp 1676037725
transform 1 0 16560 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output340
timestamp 1676037725
transform 1 0 16928 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output341
timestamp 1676037725
transform 1 0 17480 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output342
timestamp 1676037725
transform 1 0 14904 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output343
timestamp 1676037725
transform 1 0 17848 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output344
timestamp 1676037725
transform 1 0 18400 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output345
timestamp 1676037725
transform 1 0 15824 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output346
timestamp 1676037725
transform 1 0 16836 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output347
timestamp 1676037725
transform 1 0 13524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output348
timestamp 1676037725
transform 1 0 17480 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output349
timestamp 1676037725
transform 1 0 19596 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output350
timestamp 1676037725
transform 1 0 18400 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output351
timestamp 1676037725
transform 1 0 17756 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output352
timestamp 1676037725
transform 1 0 17480 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output353
timestamp 1676037725
transform 1 0 18676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output354
timestamp 1676037725
transform 1 0 18400 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output355
timestamp 1676037725
transform 1 0 22540 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output356
timestamp 1676037725
transform 1 0 22356 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output357
timestamp 1676037725
transform 1 0 22356 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output358
timestamp 1676037725
transform 1 0 14720 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output359
timestamp 1676037725
transform 1 0 19872 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output360
timestamp 1676037725
transform 1 0 20976 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output361
timestamp 1676037725
transform 1 0 22264 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output362
timestamp 1676037725
transform 1 0 25760 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output363
timestamp 1676037725
transform 1 0 22632 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output364
timestamp 1676037725
transform 1 0 25116 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output365
timestamp 1676037725
transform 1 0 23552 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output366
timestamp 1676037725
transform 1 0 25208 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output367
timestamp 1676037725
transform 1 0 13248 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output368
timestamp 1676037725
transform 1 0 15824 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output369
timestamp 1676037725
transform 1 0 1564 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output370
timestamp 1676037725
transform 1 0 1564 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output371
timestamp 1676037725
transform 1 0 1564 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output372
timestamp 1676037725
transform 1 0 1564 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output373
timestamp 1676037725
transform 1 0 1564 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output374
timestamp 1676037725
transform 1 0 1564 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output375
timestamp 1676037725
transform 1 0 1564 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output376
timestamp 1676037725
transform 1 0 1564 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output377
timestamp 1676037725
transform 1 0 1564 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output378
timestamp 1676037725
transform 1 0 1564 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output379
timestamp 1676037725
transform 1 0 1564 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output380
timestamp 1676037725
transform 1 0 1564 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output381
timestamp 1676037725
transform 1 0 1564 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output382
timestamp 1676037725
transform 1 0 57040 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output383
timestamp 1676037725
transform 1 0 56948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output384
timestamp 1676037725
transform 1 0 57868 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output385
timestamp 1676037725
transform 1 0 57868 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output386
timestamp 1676037725
transform 1 0 57868 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output387
timestamp 1676037725
transform 1 0 57868 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output388
timestamp 1676037725
transform 1 0 57868 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output389
timestamp 1676037725
transform 1 0 57868 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output390
timestamp 1676037725
transform 1 0 57868 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output391
timestamp 1676037725
transform 1 0 57868 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output392
timestamp 1676037725
transform 1 0 57868 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output393
timestamp 1676037725
transform 1 0 57868 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output394
timestamp 1676037725
transform 1 0 57868 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output395
timestamp 1676037725
transform 1 0 57868 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output396
timestamp 1676037725
transform 1 0 57868 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output397
timestamp 1676037725
transform 1 0 56948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output398
timestamp 1676037725
transform 1 0 57868 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output399
timestamp 1676037725
transform 1 0 56948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output400
timestamp 1676037725
transform 1 0 57868 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output401
timestamp 1676037725
transform 1 0 57868 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output402
timestamp 1676037725
transform 1 0 57868 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output403
timestamp 1676037725
transform 1 0 57040 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output404
timestamp 1676037725
transform 1 0 57868 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output405
timestamp 1676037725
transform 1 0 57868 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output406
timestamp 1676037725
transform 1 0 57868 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output407
timestamp 1676037725
transform 1 0 57868 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output408
timestamp 1676037725
transform 1 0 57040 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output409
timestamp 1676037725
transform 1 0 56948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output410
timestamp 1676037725
transform 1 0 57868 0 1 20672
box -38 -48 590 592
<< labels >>
flabel metal3 s 0 20952 800 21072 0 FreeSans 480 0 0 0 design_clk_o
port 0 nsew signal tristate
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 dsi_all[0]
port 1 nsew signal tristate
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 dsi_all[10]
port 2 nsew signal tristate
flabel metal3 s 0 9392 800 9512 0 FreeSans 480 0 0 0 dsi_all[11]
port 3 nsew signal tristate
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 dsi_all[12]
port 4 nsew signal tristate
flabel metal3 s 0 10752 800 10872 0 FreeSans 480 0 0 0 dsi_all[13]
port 5 nsew signal tristate
flabel metal3 s 0 11432 800 11552 0 FreeSans 480 0 0 0 dsi_all[14]
port 6 nsew signal tristate
flabel metal3 s 0 12112 800 12232 0 FreeSans 480 0 0 0 dsi_all[15]
port 7 nsew signal tristate
flabel metal3 s 0 12792 800 12912 0 FreeSans 480 0 0 0 dsi_all[16]
port 8 nsew signal tristate
flabel metal3 s 0 13472 800 13592 0 FreeSans 480 0 0 0 dsi_all[17]
port 9 nsew signal tristate
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 dsi_all[18]
port 10 nsew signal tristate
flabel metal3 s 0 14832 800 14952 0 FreeSans 480 0 0 0 dsi_all[19]
port 11 nsew signal tristate
flabel metal3 s 0 2592 800 2712 0 FreeSans 480 0 0 0 dsi_all[1]
port 12 nsew signal tristate
flabel metal3 s 0 15512 800 15632 0 FreeSans 480 0 0 0 dsi_all[20]
port 13 nsew signal tristate
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 dsi_all[21]
port 14 nsew signal tristate
flabel metal3 s 0 16872 800 16992 0 FreeSans 480 0 0 0 dsi_all[22]
port 15 nsew signal tristate
flabel metal3 s 0 17552 800 17672 0 FreeSans 480 0 0 0 dsi_all[23]
port 16 nsew signal tristate
flabel metal3 s 0 18232 800 18352 0 FreeSans 480 0 0 0 dsi_all[24]
port 17 nsew signal tristate
flabel metal3 s 0 18912 800 19032 0 FreeSans 480 0 0 0 dsi_all[25]
port 18 nsew signal tristate
flabel metal3 s 0 19592 800 19712 0 FreeSans 480 0 0 0 dsi_all[26]
port 19 nsew signal tristate
flabel metal3 s 0 20272 800 20392 0 FreeSans 480 0 0 0 dsi_all[27]
port 20 nsew signal tristate
flabel metal3 s 0 3272 800 3392 0 FreeSans 480 0 0 0 dsi_all[2]
port 21 nsew signal tristate
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 dsi_all[3]
port 22 nsew signal tristate
flabel metal3 s 0 4632 800 4752 0 FreeSans 480 0 0 0 dsi_all[4]
port 23 nsew signal tristate
flabel metal3 s 0 5312 800 5432 0 FreeSans 480 0 0 0 dsi_all[5]
port 24 nsew signal tristate
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 dsi_all[6]
port 25 nsew signal tristate
flabel metal3 s 0 6672 800 6792 0 FreeSans 480 0 0 0 dsi_all[7]
port 26 nsew signal tristate
flabel metal3 s 0 7352 800 7472 0 FreeSans 480 0 0 0 dsi_all[8]
port 27 nsew signal tristate
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 dsi_all[9]
port 28 nsew signal tristate
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 dso_6502[0]
port 29 nsew signal input
flabel metal2 s 40130 0 40186 800 0 FreeSans 224 90 0 0 dso_6502[10]
port 30 nsew signal input
flabel metal2 s 40406 0 40462 800 0 FreeSans 224 90 0 0 dso_6502[11]
port 31 nsew signal input
flabel metal2 s 40682 0 40738 800 0 FreeSans 224 90 0 0 dso_6502[12]
port 32 nsew signal input
flabel metal2 s 40958 0 41014 800 0 FreeSans 224 90 0 0 dso_6502[13]
port 33 nsew signal input
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 dso_6502[14]
port 34 nsew signal input
flabel metal2 s 41510 0 41566 800 0 FreeSans 224 90 0 0 dso_6502[15]
port 35 nsew signal input
flabel metal2 s 41786 0 41842 800 0 FreeSans 224 90 0 0 dso_6502[16]
port 36 nsew signal input
flabel metal2 s 42062 0 42118 800 0 FreeSans 224 90 0 0 dso_6502[17]
port 37 nsew signal input
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 dso_6502[18]
port 38 nsew signal input
flabel metal2 s 42614 0 42670 800 0 FreeSans 224 90 0 0 dso_6502[19]
port 39 nsew signal input
flabel metal2 s 37646 0 37702 800 0 FreeSans 224 90 0 0 dso_6502[1]
port 40 nsew signal input
flabel metal2 s 42890 0 42946 800 0 FreeSans 224 90 0 0 dso_6502[20]
port 41 nsew signal input
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 dso_6502[21]
port 42 nsew signal input
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 dso_6502[22]
port 43 nsew signal input
flabel metal2 s 43718 0 43774 800 0 FreeSans 224 90 0 0 dso_6502[23]
port 44 nsew signal input
flabel metal2 s 43994 0 44050 800 0 FreeSans 224 90 0 0 dso_6502[24]
port 45 nsew signal input
flabel metal2 s 44270 0 44326 800 0 FreeSans 224 90 0 0 dso_6502[25]
port 46 nsew signal input
flabel metal2 s 44546 0 44602 800 0 FreeSans 224 90 0 0 dso_6502[26]
port 47 nsew signal input
flabel metal2 s 37922 0 37978 800 0 FreeSans 224 90 0 0 dso_6502[2]
port 48 nsew signal input
flabel metal2 s 38198 0 38254 800 0 FreeSans 224 90 0 0 dso_6502[3]
port 49 nsew signal input
flabel metal2 s 38474 0 38530 800 0 FreeSans 224 90 0 0 dso_6502[4]
port 50 nsew signal input
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 dso_6502[5]
port 51 nsew signal input
flabel metal2 s 39026 0 39082 800 0 FreeSans 224 90 0 0 dso_6502[6]
port 52 nsew signal input
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 dso_6502[7]
port 53 nsew signal input
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 dso_6502[8]
port 54 nsew signal input
flabel metal2 s 39854 0 39910 800 0 FreeSans 224 90 0 0 dso_6502[9]
port 55 nsew signal input
flabel metal2 s 53838 63200 53894 64000 0 FreeSans 224 90 0 0 dso_LCD[0]
port 56 nsew signal input
flabel metal2 s 54574 63200 54630 64000 0 FreeSans 224 90 0 0 dso_LCD[1]
port 57 nsew signal input
flabel metal2 s 55310 63200 55366 64000 0 FreeSans 224 90 0 0 dso_LCD[2]
port 58 nsew signal input
flabel metal2 s 56046 63200 56102 64000 0 FreeSans 224 90 0 0 dso_LCD[3]
port 59 nsew signal input
flabel metal2 s 56782 63200 56838 64000 0 FreeSans 224 90 0 0 dso_LCD[4]
port 60 nsew signal input
flabel metal2 s 57518 63200 57574 64000 0 FreeSans 224 90 0 0 dso_LCD[5]
port 61 nsew signal input
flabel metal2 s 58254 63200 58310 64000 0 FreeSans 224 90 0 0 dso_LCD[6]
port 62 nsew signal input
flabel metal2 s 58990 63200 59046 64000 0 FreeSans 224 90 0 0 dso_LCD[7]
port 63 nsew signal input
flabel metal2 s 44822 0 44878 800 0 FreeSans 224 90 0 0 dso_as1802[0]
port 64 nsew signal input
flabel metal2 s 47582 0 47638 800 0 FreeSans 224 90 0 0 dso_as1802[10]
port 65 nsew signal input
flabel metal2 s 47858 0 47914 800 0 FreeSans 224 90 0 0 dso_as1802[11]
port 66 nsew signal input
flabel metal2 s 48134 0 48190 800 0 FreeSans 224 90 0 0 dso_as1802[12]
port 67 nsew signal input
flabel metal2 s 48410 0 48466 800 0 FreeSans 224 90 0 0 dso_as1802[13]
port 68 nsew signal input
flabel metal2 s 48686 0 48742 800 0 FreeSans 224 90 0 0 dso_as1802[14]
port 69 nsew signal input
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 dso_as1802[15]
port 70 nsew signal input
flabel metal2 s 49238 0 49294 800 0 FreeSans 224 90 0 0 dso_as1802[16]
port 71 nsew signal input
flabel metal2 s 49514 0 49570 800 0 FreeSans 224 90 0 0 dso_as1802[17]
port 72 nsew signal input
flabel metal2 s 49790 0 49846 800 0 FreeSans 224 90 0 0 dso_as1802[18]
port 73 nsew signal input
flabel metal2 s 50066 0 50122 800 0 FreeSans 224 90 0 0 dso_as1802[19]
port 74 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 dso_as1802[1]
port 75 nsew signal input
flabel metal2 s 50342 0 50398 800 0 FreeSans 224 90 0 0 dso_as1802[20]
port 76 nsew signal input
flabel metal2 s 50618 0 50674 800 0 FreeSans 224 90 0 0 dso_as1802[21]
port 77 nsew signal input
flabel metal2 s 50894 0 50950 800 0 FreeSans 224 90 0 0 dso_as1802[22]
port 78 nsew signal input
flabel metal2 s 51170 0 51226 800 0 FreeSans 224 90 0 0 dso_as1802[23]
port 79 nsew signal input
flabel metal2 s 51446 0 51502 800 0 FreeSans 224 90 0 0 dso_as1802[24]
port 80 nsew signal input
flabel metal2 s 51722 0 51778 800 0 FreeSans 224 90 0 0 dso_as1802[25]
port 81 nsew signal input
flabel metal2 s 51998 0 52054 800 0 FreeSans 224 90 0 0 dso_as1802[26]
port 82 nsew signal input
flabel metal2 s 45374 0 45430 800 0 FreeSans 224 90 0 0 dso_as1802[2]
port 83 nsew signal input
flabel metal2 s 45650 0 45706 800 0 FreeSans 224 90 0 0 dso_as1802[3]
port 84 nsew signal input
flabel metal2 s 45926 0 45982 800 0 FreeSans 224 90 0 0 dso_as1802[4]
port 85 nsew signal input
flabel metal2 s 46202 0 46258 800 0 FreeSans 224 90 0 0 dso_as1802[5]
port 86 nsew signal input
flabel metal2 s 46478 0 46534 800 0 FreeSans 224 90 0 0 dso_as1802[6]
port 87 nsew signal input
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 dso_as1802[7]
port 88 nsew signal input
flabel metal2 s 47030 0 47086 800 0 FreeSans 224 90 0 0 dso_as1802[8]
port 89 nsew signal input
flabel metal2 s 47306 0 47362 800 0 FreeSans 224 90 0 0 dso_as1802[9]
port 90 nsew signal input
flabel metal2 s 13358 63200 13414 64000 0 FreeSans 224 90 0 0 dso_as2650[0]
port 91 nsew signal input
flabel metal2 s 20718 63200 20774 64000 0 FreeSans 224 90 0 0 dso_as2650[10]
port 92 nsew signal input
flabel metal2 s 21454 63200 21510 64000 0 FreeSans 224 90 0 0 dso_as2650[11]
port 93 nsew signal input
flabel metal2 s 22190 63200 22246 64000 0 FreeSans 224 90 0 0 dso_as2650[12]
port 94 nsew signal input
flabel metal2 s 22926 63200 22982 64000 0 FreeSans 224 90 0 0 dso_as2650[13]
port 95 nsew signal input
flabel metal2 s 23662 63200 23718 64000 0 FreeSans 224 90 0 0 dso_as2650[14]
port 96 nsew signal input
flabel metal2 s 24398 63200 24454 64000 0 FreeSans 224 90 0 0 dso_as2650[15]
port 97 nsew signal input
flabel metal2 s 25134 63200 25190 64000 0 FreeSans 224 90 0 0 dso_as2650[16]
port 98 nsew signal input
flabel metal2 s 25870 63200 25926 64000 0 FreeSans 224 90 0 0 dso_as2650[17]
port 99 nsew signal input
flabel metal2 s 26606 63200 26662 64000 0 FreeSans 224 90 0 0 dso_as2650[18]
port 100 nsew signal input
flabel metal2 s 27342 63200 27398 64000 0 FreeSans 224 90 0 0 dso_as2650[19]
port 101 nsew signal input
flabel metal2 s 14094 63200 14150 64000 0 FreeSans 224 90 0 0 dso_as2650[1]
port 102 nsew signal input
flabel metal2 s 28078 63200 28134 64000 0 FreeSans 224 90 0 0 dso_as2650[20]
port 103 nsew signal input
flabel metal2 s 28814 63200 28870 64000 0 FreeSans 224 90 0 0 dso_as2650[21]
port 104 nsew signal input
flabel metal2 s 29550 63200 29606 64000 0 FreeSans 224 90 0 0 dso_as2650[22]
port 105 nsew signal input
flabel metal2 s 30286 63200 30342 64000 0 FreeSans 224 90 0 0 dso_as2650[23]
port 106 nsew signal input
flabel metal2 s 31022 63200 31078 64000 0 FreeSans 224 90 0 0 dso_as2650[24]
port 107 nsew signal input
flabel metal2 s 31758 63200 31814 64000 0 FreeSans 224 90 0 0 dso_as2650[25]
port 108 nsew signal input
flabel metal2 s 32494 63200 32550 64000 0 FreeSans 224 90 0 0 dso_as2650[26]
port 109 nsew signal input
flabel metal2 s 14830 63200 14886 64000 0 FreeSans 224 90 0 0 dso_as2650[2]
port 110 nsew signal input
flabel metal2 s 15566 63200 15622 64000 0 FreeSans 224 90 0 0 dso_as2650[3]
port 111 nsew signal input
flabel metal2 s 16302 63200 16358 64000 0 FreeSans 224 90 0 0 dso_as2650[4]
port 112 nsew signal input
flabel metal2 s 17038 63200 17094 64000 0 FreeSans 224 90 0 0 dso_as2650[5]
port 113 nsew signal input
flabel metal2 s 17774 63200 17830 64000 0 FreeSans 224 90 0 0 dso_as2650[6]
port 114 nsew signal input
flabel metal2 s 18510 63200 18566 64000 0 FreeSans 224 90 0 0 dso_as2650[7]
port 115 nsew signal input
flabel metal2 s 19246 63200 19302 64000 0 FreeSans 224 90 0 0 dso_as2650[8]
port 116 nsew signal input
flabel metal2 s 19982 63200 20038 64000 0 FreeSans 224 90 0 0 dso_as2650[9]
port 117 nsew signal input
flabel metal3 s 0 42712 800 42832 0 FreeSans 480 0 0 0 dso_as512512512[0]
port 118 nsew signal input
flabel metal3 s 0 49512 800 49632 0 FreeSans 480 0 0 0 dso_as512512512[10]
port 119 nsew signal input
flabel metal3 s 0 50192 800 50312 0 FreeSans 480 0 0 0 dso_as512512512[11]
port 120 nsew signal input
flabel metal3 s 0 50872 800 50992 0 FreeSans 480 0 0 0 dso_as512512512[12]
port 121 nsew signal input
flabel metal3 s 0 51552 800 51672 0 FreeSans 480 0 0 0 dso_as512512512[13]
port 122 nsew signal input
flabel metal3 s 0 52232 800 52352 0 FreeSans 480 0 0 0 dso_as512512512[14]
port 123 nsew signal input
flabel metal3 s 0 52912 800 53032 0 FreeSans 480 0 0 0 dso_as512512512[15]
port 124 nsew signal input
flabel metal3 s 0 53592 800 53712 0 FreeSans 480 0 0 0 dso_as512512512[16]
port 125 nsew signal input
flabel metal3 s 0 54272 800 54392 0 FreeSans 480 0 0 0 dso_as512512512[17]
port 126 nsew signal input
flabel metal3 s 0 54952 800 55072 0 FreeSans 480 0 0 0 dso_as512512512[18]
port 127 nsew signal input
flabel metal3 s 0 55632 800 55752 0 FreeSans 480 0 0 0 dso_as512512512[19]
port 128 nsew signal input
flabel metal3 s 0 43392 800 43512 0 FreeSans 480 0 0 0 dso_as512512512[1]
port 129 nsew signal input
flabel metal3 s 0 56312 800 56432 0 FreeSans 480 0 0 0 dso_as512512512[20]
port 130 nsew signal input
flabel metal3 s 0 56992 800 57112 0 FreeSans 480 0 0 0 dso_as512512512[21]
port 131 nsew signal input
flabel metal3 s 0 57672 800 57792 0 FreeSans 480 0 0 0 dso_as512512512[22]
port 132 nsew signal input
flabel metal3 s 0 58352 800 58472 0 FreeSans 480 0 0 0 dso_as512512512[23]
port 133 nsew signal input
flabel metal3 s 0 59032 800 59152 0 FreeSans 480 0 0 0 dso_as512512512[24]
port 134 nsew signal input
flabel metal3 s 0 59712 800 59832 0 FreeSans 480 0 0 0 dso_as512512512[25]
port 135 nsew signal input
flabel metal3 s 0 60392 800 60512 0 FreeSans 480 0 0 0 dso_as512512512[26]
port 136 nsew signal input
flabel metal3 s 0 61072 800 61192 0 FreeSans 480 0 0 0 dso_as512512512[27]
port 137 nsew signal input
flabel metal3 s 0 44072 800 44192 0 FreeSans 480 0 0 0 dso_as512512512[2]
port 138 nsew signal input
flabel metal3 s 0 44752 800 44872 0 FreeSans 480 0 0 0 dso_as512512512[3]
port 139 nsew signal input
flabel metal3 s 0 45432 800 45552 0 FreeSans 480 0 0 0 dso_as512512512[4]
port 140 nsew signal input
flabel metal3 s 0 46112 800 46232 0 FreeSans 480 0 0 0 dso_as512512512[5]
port 141 nsew signal input
flabel metal3 s 0 46792 800 46912 0 FreeSans 480 0 0 0 dso_as512512512[6]
port 142 nsew signal input
flabel metal3 s 0 47472 800 47592 0 FreeSans 480 0 0 0 dso_as512512512[7]
port 143 nsew signal input
flabel metal3 s 0 48152 800 48272 0 FreeSans 480 0 0 0 dso_as512512512[8]
port 144 nsew signal input
flabel metal3 s 0 48832 800 48952 0 FreeSans 480 0 0 0 dso_as512512512[9]
port 145 nsew signal input
flabel metal2 s 33230 63200 33286 64000 0 FreeSans 224 90 0 0 dso_as5401[0]
port 146 nsew signal input
flabel metal2 s 40590 63200 40646 64000 0 FreeSans 224 90 0 0 dso_as5401[10]
port 147 nsew signal input
flabel metal2 s 41326 63200 41382 64000 0 FreeSans 224 90 0 0 dso_as5401[11]
port 148 nsew signal input
flabel metal2 s 42062 63200 42118 64000 0 FreeSans 224 90 0 0 dso_as5401[12]
port 149 nsew signal input
flabel metal2 s 42798 63200 42854 64000 0 FreeSans 224 90 0 0 dso_as5401[13]
port 150 nsew signal input
flabel metal2 s 43534 63200 43590 64000 0 FreeSans 224 90 0 0 dso_as5401[14]
port 151 nsew signal input
flabel metal2 s 44270 63200 44326 64000 0 FreeSans 224 90 0 0 dso_as5401[15]
port 152 nsew signal input
flabel metal2 s 45006 63200 45062 64000 0 FreeSans 224 90 0 0 dso_as5401[16]
port 153 nsew signal input
flabel metal2 s 45742 63200 45798 64000 0 FreeSans 224 90 0 0 dso_as5401[17]
port 154 nsew signal input
flabel metal2 s 46478 63200 46534 64000 0 FreeSans 224 90 0 0 dso_as5401[18]
port 155 nsew signal input
flabel metal2 s 47214 63200 47270 64000 0 FreeSans 224 90 0 0 dso_as5401[19]
port 156 nsew signal input
flabel metal2 s 33966 63200 34022 64000 0 FreeSans 224 90 0 0 dso_as5401[1]
port 157 nsew signal input
flabel metal2 s 47950 63200 48006 64000 0 FreeSans 224 90 0 0 dso_as5401[20]
port 158 nsew signal input
flabel metal2 s 48686 63200 48742 64000 0 FreeSans 224 90 0 0 dso_as5401[21]
port 159 nsew signal input
flabel metal2 s 49422 63200 49478 64000 0 FreeSans 224 90 0 0 dso_as5401[22]
port 160 nsew signal input
flabel metal2 s 50158 63200 50214 64000 0 FreeSans 224 90 0 0 dso_as5401[23]
port 161 nsew signal input
flabel metal2 s 50894 63200 50950 64000 0 FreeSans 224 90 0 0 dso_as5401[24]
port 162 nsew signal input
flabel metal2 s 51630 63200 51686 64000 0 FreeSans 224 90 0 0 dso_as5401[25]
port 163 nsew signal input
flabel metal2 s 52366 63200 52422 64000 0 FreeSans 224 90 0 0 dso_as5401[26]
port 164 nsew signal input
flabel metal2 s 34702 63200 34758 64000 0 FreeSans 224 90 0 0 dso_as5401[2]
port 165 nsew signal input
flabel metal2 s 35438 63200 35494 64000 0 FreeSans 224 90 0 0 dso_as5401[3]
port 166 nsew signal input
flabel metal2 s 36174 63200 36230 64000 0 FreeSans 224 90 0 0 dso_as5401[4]
port 167 nsew signal input
flabel metal2 s 36910 63200 36966 64000 0 FreeSans 224 90 0 0 dso_as5401[5]
port 168 nsew signal input
flabel metal2 s 37646 63200 37702 64000 0 FreeSans 224 90 0 0 dso_as5401[6]
port 169 nsew signal input
flabel metal2 s 38382 63200 38438 64000 0 FreeSans 224 90 0 0 dso_as5401[7]
port 170 nsew signal input
flabel metal2 s 39118 63200 39174 64000 0 FreeSans 224 90 0 0 dso_as5401[8]
port 171 nsew signal input
flabel metal2 s 39854 63200 39910 64000 0 FreeSans 224 90 0 0 dso_as5401[9]
port 172 nsew signal input
flabel metal3 s 59200 56584 60000 56704 0 FreeSans 480 0 0 0 dso_counter[0]
port 173 nsew signal input
flabel metal3 s 59200 62024 60000 62144 0 FreeSans 480 0 0 0 dso_counter[10]
port 174 nsew signal input
flabel metal3 s 59200 62568 60000 62688 0 FreeSans 480 0 0 0 dso_counter[11]
port 175 nsew signal input
flabel metal3 s 59200 57128 60000 57248 0 FreeSans 480 0 0 0 dso_counter[1]
port 176 nsew signal input
flabel metal3 s 59200 57672 60000 57792 0 FreeSans 480 0 0 0 dso_counter[2]
port 177 nsew signal input
flabel metal3 s 59200 58216 60000 58336 0 FreeSans 480 0 0 0 dso_counter[3]
port 178 nsew signal input
flabel metal3 s 59200 58760 60000 58880 0 FreeSans 480 0 0 0 dso_counter[4]
port 179 nsew signal input
flabel metal3 s 59200 59304 60000 59424 0 FreeSans 480 0 0 0 dso_counter[5]
port 180 nsew signal input
flabel metal3 s 59200 59848 60000 59968 0 FreeSans 480 0 0 0 dso_counter[6]
port 181 nsew signal input
flabel metal3 s 59200 60392 60000 60512 0 FreeSans 480 0 0 0 dso_counter[7]
port 182 nsew signal input
flabel metal3 s 59200 60936 60000 61056 0 FreeSans 480 0 0 0 dso_counter[8]
port 183 nsew signal input
flabel metal3 s 59200 61480 60000 61600 0 FreeSans 480 0 0 0 dso_counter[9]
port 184 nsew signal input
flabel metal2 s 6734 63200 6790 64000 0 FreeSans 224 90 0 0 dso_diceroll[0]
port 185 nsew signal input
flabel metal2 s 7470 63200 7526 64000 0 FreeSans 224 90 0 0 dso_diceroll[1]
port 186 nsew signal input
flabel metal2 s 8206 63200 8262 64000 0 FreeSans 224 90 0 0 dso_diceroll[2]
port 187 nsew signal input
flabel metal2 s 8942 63200 8998 64000 0 FreeSans 224 90 0 0 dso_diceroll[3]
port 188 nsew signal input
flabel metal2 s 9678 63200 9734 64000 0 FreeSans 224 90 0 0 dso_diceroll[4]
port 189 nsew signal input
flabel metal2 s 10414 63200 10470 64000 0 FreeSans 224 90 0 0 dso_diceroll[5]
port 190 nsew signal input
flabel metal2 s 11150 63200 11206 64000 0 FreeSans 224 90 0 0 dso_diceroll[6]
port 191 nsew signal input
flabel metal2 s 11886 63200 11942 64000 0 FreeSans 224 90 0 0 dso_diceroll[7]
port 192 nsew signal input
flabel metal3 s 0 30472 800 30592 0 FreeSans 480 0 0 0 dso_mc14500[0]
port 193 nsew signal input
flabel metal3 s 0 31152 800 31272 0 FreeSans 480 0 0 0 dso_mc14500[1]
port 194 nsew signal input
flabel metal3 s 0 31832 800 31952 0 FreeSans 480 0 0 0 dso_mc14500[2]
port 195 nsew signal input
flabel metal3 s 0 32512 800 32632 0 FreeSans 480 0 0 0 dso_mc14500[3]
port 196 nsew signal input
flabel metal3 s 0 33192 800 33312 0 FreeSans 480 0 0 0 dso_mc14500[4]
port 197 nsew signal input
flabel metal3 s 0 33872 800 33992 0 FreeSans 480 0 0 0 dso_mc14500[5]
port 198 nsew signal input
flabel metal3 s 0 34552 800 34672 0 FreeSans 480 0 0 0 dso_mc14500[6]
port 199 nsew signal input
flabel metal3 s 0 35232 800 35352 0 FreeSans 480 0 0 0 dso_mc14500[7]
port 200 nsew signal input
flabel metal3 s 0 35912 800 36032 0 FreeSans 480 0 0 0 dso_mc14500[8]
port 201 nsew signal input
flabel metal2 s 846 63200 902 64000 0 FreeSans 224 90 0 0 dso_multiplier[0]
port 202 nsew signal input
flabel metal2 s 1582 63200 1638 64000 0 FreeSans 224 90 0 0 dso_multiplier[1]
port 203 nsew signal input
flabel metal2 s 2318 63200 2374 64000 0 FreeSans 224 90 0 0 dso_multiplier[2]
port 204 nsew signal input
flabel metal2 s 3054 63200 3110 64000 0 FreeSans 224 90 0 0 dso_multiplier[3]
port 205 nsew signal input
flabel metal2 s 3790 63200 3846 64000 0 FreeSans 224 90 0 0 dso_multiplier[4]
port 206 nsew signal input
flabel metal2 s 4526 63200 4582 64000 0 FreeSans 224 90 0 0 dso_multiplier[5]
port 207 nsew signal input
flabel metal2 s 5262 63200 5318 64000 0 FreeSans 224 90 0 0 dso_multiplier[6]
port 208 nsew signal input
flabel metal2 s 5998 63200 6054 64000 0 FreeSans 224 90 0 0 dso_multiplier[7]
port 209 nsew signal input
flabel metal2 s 35990 0 36046 800 0 FreeSans 224 90 0 0 dso_posit[0]
port 210 nsew signal input
flabel metal2 s 36266 0 36322 800 0 FreeSans 224 90 0 0 dso_posit[1]
port 211 nsew signal input
flabel metal2 s 36542 0 36598 800 0 FreeSans 224 90 0 0 dso_posit[2]
port 212 nsew signal input
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 dso_posit[3]
port 213 nsew signal input
flabel metal3 s 0 37272 800 37392 0 FreeSans 480 0 0 0 dso_tbb1143[0]
port 214 nsew signal input
flabel metal3 s 0 37952 800 38072 0 FreeSans 480 0 0 0 dso_tbb1143[1]
port 215 nsew signal input
flabel metal3 s 0 38632 800 38752 0 FreeSans 480 0 0 0 dso_tbb1143[2]
port 216 nsew signal input
flabel metal3 s 0 39312 800 39432 0 FreeSans 480 0 0 0 dso_tbb1143[3]
port 217 nsew signal input
flabel metal3 s 0 39992 800 40112 0 FreeSans 480 0 0 0 dso_tbb1143[4]
port 218 nsew signal input
flabel metal3 s 0 40672 800 40792 0 FreeSans 480 0 0 0 dso_tbb1143[5]
port 219 nsew signal input
flabel metal3 s 0 41352 800 41472 0 FreeSans 480 0 0 0 dso_tbb1143[6]
port 220 nsew signal input
flabel metal3 s 0 42032 800 42152 0 FreeSans 480 0 0 0 dso_tbb1143[7]
port 221 nsew signal input
flabel metal2 s 52550 0 52606 800 0 FreeSans 224 90 0 0 dso_tune
port 222 nsew signal input
flabel metal2 s 52826 0 52882 800 0 FreeSans 224 90 0 0 dso_vgatest[0]
port 223 nsew signal input
flabel metal2 s 53102 0 53158 800 0 FreeSans 224 90 0 0 dso_vgatest[1]
port 224 nsew signal input
flabel metal2 s 53378 0 53434 800 0 FreeSans 224 90 0 0 dso_vgatest[2]
port 225 nsew signal input
flabel metal2 s 53654 0 53710 800 0 FreeSans 224 90 0 0 dso_vgatest[3]
port 226 nsew signal input
flabel metal2 s 53930 0 53986 800 0 FreeSans 224 90 0 0 dso_vgatest[4]
port 227 nsew signal input
flabel metal2 s 54206 0 54262 800 0 FreeSans 224 90 0 0 dso_vgatest[5]
port 228 nsew signal input
flabel metal2 s 54482 0 54538 800 0 FreeSans 224 90 0 0 dso_vgatest[6]
port 229 nsew signal input
flabel metal2 s 54758 0 54814 800 0 FreeSans 224 90 0 0 dso_vgatest[7]
port 230 nsew signal input
flabel metal2 s 55034 0 55090 800 0 FreeSans 224 90 0 0 dso_vgatest[8]
port 231 nsew signal input
flabel metal2 s 55310 0 55366 800 0 FreeSans 224 90 0 0 dso_vgatest[9]
port 232 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 io_in[0]
port 233 nsew signal input
flabel metal2 s 7286 0 7342 800 0 FreeSans 224 90 0 0 io_in[10]
port 234 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 io_in[11]
port 235 nsew signal input
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 io_in[12]
port 236 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 io_in[13]
port 237 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 io_in[14]
port 238 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 io_in[15]
port 239 nsew signal input
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 io_in[16]
port 240 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 io_in[17]
port 241 nsew signal input
flabel metal2 s 9494 0 9550 800 0 FreeSans 224 90 0 0 io_in[18]
port 242 nsew signal input
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 io_in[19]
port 243 nsew signal input
flabel metal2 s 4802 0 4858 800 0 FreeSans 224 90 0 0 io_in[1]
port 244 nsew signal input
flabel metal2 s 10046 0 10102 800 0 FreeSans 224 90 0 0 io_in[20]
port 245 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 io_in[21]
port 246 nsew signal input
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 io_in[22]
port 247 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 io_in[23]
port 248 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 io_in[24]
port 249 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 io_in[25]
port 250 nsew signal input
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 io_in[26]
port 251 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 io_in[27]
port 252 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 io_in[28]
port 253 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 io_in[29]
port 254 nsew signal input
flabel metal2 s 5078 0 5134 800 0 FreeSans 224 90 0 0 io_in[2]
port 255 nsew signal input
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 io_in[30]
port 256 nsew signal input
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 io_in[31]
port 257 nsew signal input
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 io_in[32]
port 258 nsew signal input
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 io_in[33]
port 259 nsew signal input
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 io_in[34]
port 260 nsew signal input
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 io_in[35]
port 261 nsew signal input
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 io_in[36]
port 262 nsew signal input
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 io_in[37]
port 263 nsew signal input
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 io_in[3]
port 264 nsew signal input
flabel metal2 s 5630 0 5686 800 0 FreeSans 224 90 0 0 io_in[4]
port 265 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 io_in[5]
port 266 nsew signal input
flabel metal2 s 6182 0 6238 800 0 FreeSans 224 90 0 0 io_in[6]
port 267 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 io_in[7]
port 268 nsew signal input
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 io_in[8]
port 269 nsew signal input
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 io_in[9]
port 270 nsew signal input
flabel metal2 s 25502 0 25558 800 0 FreeSans 224 90 0 0 io_oeb[0]
port 271 nsew signal tristate
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 io_oeb[10]
port 272 nsew signal tristate
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 io_oeb[11]
port 273 nsew signal tristate
flabel metal2 s 28814 0 28870 800 0 FreeSans 224 90 0 0 io_oeb[12]
port 274 nsew signal tristate
flabel metal2 s 29090 0 29146 800 0 FreeSans 224 90 0 0 io_oeb[13]
port 275 nsew signal tristate
flabel metal2 s 29366 0 29422 800 0 FreeSans 224 90 0 0 io_oeb[14]
port 276 nsew signal tristate
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 io_oeb[15]
port 277 nsew signal tristate
flabel metal2 s 29918 0 29974 800 0 FreeSans 224 90 0 0 io_oeb[16]
port 278 nsew signal tristate
flabel metal2 s 30194 0 30250 800 0 FreeSans 224 90 0 0 io_oeb[17]
port 279 nsew signal tristate
flabel metal2 s 30470 0 30526 800 0 FreeSans 224 90 0 0 io_oeb[18]
port 280 nsew signal tristate
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 io_oeb[19]
port 281 nsew signal tristate
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 io_oeb[1]
port 282 nsew signal tristate
flabel metal2 s 31022 0 31078 800 0 FreeSans 224 90 0 0 io_oeb[20]
port 283 nsew signal tristate
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 io_oeb[21]
port 284 nsew signal tristate
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 io_oeb[22]
port 285 nsew signal tristate
flabel metal2 s 31850 0 31906 800 0 FreeSans 224 90 0 0 io_oeb[23]
port 286 nsew signal tristate
flabel metal2 s 32126 0 32182 800 0 FreeSans 224 90 0 0 io_oeb[24]
port 287 nsew signal tristate
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 io_oeb[25]
port 288 nsew signal tristate
flabel metal2 s 32678 0 32734 800 0 FreeSans 224 90 0 0 io_oeb[26]
port 289 nsew signal tristate
flabel metal2 s 32954 0 33010 800 0 FreeSans 224 90 0 0 io_oeb[27]
port 290 nsew signal tristate
flabel metal2 s 33230 0 33286 800 0 FreeSans 224 90 0 0 io_oeb[28]
port 291 nsew signal tristate
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 io_oeb[29]
port 292 nsew signal tristate
flabel metal2 s 26054 0 26110 800 0 FreeSans 224 90 0 0 io_oeb[2]
port 293 nsew signal tristate
flabel metal2 s 33782 0 33838 800 0 FreeSans 224 90 0 0 io_oeb[30]
port 294 nsew signal tristate
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 io_oeb[31]
port 295 nsew signal tristate
flabel metal2 s 34334 0 34390 800 0 FreeSans 224 90 0 0 io_oeb[32]
port 296 nsew signal tristate
flabel metal2 s 34610 0 34666 800 0 FreeSans 224 90 0 0 io_oeb[33]
port 297 nsew signal tristate
flabel metal2 s 34886 0 34942 800 0 FreeSans 224 90 0 0 io_oeb[34]
port 298 nsew signal tristate
flabel metal2 s 35162 0 35218 800 0 FreeSans 224 90 0 0 io_oeb[35]
port 299 nsew signal tristate
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 io_oeb[36]
port 300 nsew signal tristate
flabel metal2 s 35714 0 35770 800 0 FreeSans 224 90 0 0 io_oeb[37]
port 301 nsew signal tristate
flabel metal2 s 26330 0 26386 800 0 FreeSans 224 90 0 0 io_oeb[3]
port 302 nsew signal tristate
flabel metal2 s 26606 0 26662 800 0 FreeSans 224 90 0 0 io_oeb[4]
port 303 nsew signal tristate
flabel metal2 s 26882 0 26938 800 0 FreeSans 224 90 0 0 io_oeb[5]
port 304 nsew signal tristate
flabel metal2 s 27158 0 27214 800 0 FreeSans 224 90 0 0 io_oeb[6]
port 305 nsew signal tristate
flabel metal2 s 27434 0 27490 800 0 FreeSans 224 90 0 0 io_oeb[7]
port 306 nsew signal tristate
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 io_oeb[8]
port 307 nsew signal tristate
flabel metal2 s 27986 0 28042 800 0 FreeSans 224 90 0 0 io_oeb[9]
port 308 nsew signal tristate
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 io_out[0]
port 309 nsew signal tristate
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 io_out[10]
port 310 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 io_out[11]
port 311 nsew signal tristate
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 io_out[12]
port 312 nsew signal tristate
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 io_out[13]
port 313 nsew signal tristate
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 io_out[14]
port 314 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 io_out[15]
port 315 nsew signal tristate
flabel metal2 s 19430 0 19486 800 0 FreeSans 224 90 0 0 io_out[16]
port 316 nsew signal tristate
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 io_out[17]
port 317 nsew signal tristate
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 io_out[18]
port 318 nsew signal tristate
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 io_out[19]
port 319 nsew signal tristate
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 io_out[1]
port 320 nsew signal tristate
flabel metal2 s 20534 0 20590 800 0 FreeSans 224 90 0 0 io_out[20]
port 321 nsew signal tristate
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 io_out[21]
port 322 nsew signal tristate
flabel metal2 s 21086 0 21142 800 0 FreeSans 224 90 0 0 io_out[22]
port 323 nsew signal tristate
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 io_out[23]
port 324 nsew signal tristate
flabel metal2 s 21638 0 21694 800 0 FreeSans 224 90 0 0 io_out[24]
port 325 nsew signal tristate
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 io_out[25]
port 326 nsew signal tristate
flabel metal2 s 22190 0 22246 800 0 FreeSans 224 90 0 0 io_out[26]
port 327 nsew signal tristate
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 io_out[27]
port 328 nsew signal tristate
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 io_out[28]
port 329 nsew signal tristate
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 io_out[29]
port 330 nsew signal tristate
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 io_out[2]
port 331 nsew signal tristate
flabel metal2 s 23294 0 23350 800 0 FreeSans 224 90 0 0 io_out[30]
port 332 nsew signal tristate
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 io_out[31]
port 333 nsew signal tristate
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 io_out[32]
port 334 nsew signal tristate
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 io_out[33]
port 335 nsew signal tristate
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 io_out[34]
port 336 nsew signal tristate
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 io_out[35]
port 337 nsew signal tristate
flabel metal2 s 24950 0 25006 800 0 FreeSans 224 90 0 0 io_out[36]
port 338 nsew signal tristate
flabel metal2 s 25226 0 25282 800 0 FreeSans 224 90 0 0 io_out[37]
port 339 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 io_out[3]
port 340 nsew signal tristate
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 io_out[4]
port 341 nsew signal tristate
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 io_out[5]
port 342 nsew signal tristate
flabel metal2 s 16670 0 16726 800 0 FreeSans 224 90 0 0 io_out[6]
port 343 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 io_out[7]
port 344 nsew signal tristate
flabel metal2 s 17222 0 17278 800 0 FreeSans 224 90 0 0 io_out[8]
port 345 nsew signal tristate
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 io_out[9]
port 346 nsew signal tristate
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 oeb_6502
port 347 nsew signal input
flabel metal2 s 52274 0 52330 800 0 FreeSans 224 90 0 0 oeb_as1802
port 348 nsew signal input
flabel metal2 s 12622 63200 12678 64000 0 FreeSans 224 90 0 0 oeb_as2650
port 349 nsew signal input
flabel metal3 s 0 61752 800 61872 0 FreeSans 480 0 0 0 oeb_as512512512
port 350 nsew signal input
flabel metal2 s 53102 63200 53158 64000 0 FreeSans 224 90 0 0 oeb_as5401
port 351 nsew signal input
flabel metal3 s 0 36592 800 36712 0 FreeSans 480 0 0 0 oeb_mc14500
port 352 nsew signal input
flabel metal3 s 0 21632 800 21752 0 FreeSans 480 0 0 0 rst_6502
port 353 nsew signal tristate
flabel metal3 s 0 22312 800 22432 0 FreeSans 480 0 0 0 rst_LCD
port 354 nsew signal tristate
flabel metal3 s 0 22992 800 23112 0 FreeSans 480 0 0 0 rst_as1802
port 355 nsew signal tristate
flabel metal3 s 0 23672 800 23792 0 FreeSans 480 0 0 0 rst_as2650
port 356 nsew signal tristate
flabel metal3 s 0 25032 800 25152 0 FreeSans 480 0 0 0 rst_as512512512
port 357 nsew signal tristate
flabel metal3 s 0 24352 800 24472 0 FreeSans 480 0 0 0 rst_as5401
port 358 nsew signal tristate
flabel metal3 s 0 25712 800 25832 0 FreeSans 480 0 0 0 rst_counter
port 359 nsew signal tristate
flabel metal3 s 0 26392 800 26512 0 FreeSans 480 0 0 0 rst_diceroll
port 360 nsew signal tristate
flabel metal3 s 0 27072 800 27192 0 FreeSans 480 0 0 0 rst_mc14500
port 361 nsew signal tristate
flabel metal3 s 0 27752 800 27872 0 FreeSans 480 0 0 0 rst_posit
port 362 nsew signal tristate
flabel metal3 s 0 28432 800 28552 0 FreeSans 480 0 0 0 rst_tbb1143
port 363 nsew signal tristate
flabel metal3 s 0 29112 800 29232 0 FreeSans 480 0 0 0 rst_tune
port 364 nsew signal tristate
flabel metal3 s 0 29792 800 29912 0 FreeSans 480 0 0 0 rst_vgatest
port 365 nsew signal tristate
flabel metal4 s 4208 2128 4528 61520 0 FreeSans 1920 90 0 0 vccd1
port 366 nsew power bidirectional
flabel metal4 s 34928 2128 35248 61520 0 FreeSans 1920 90 0 0 vccd1
port 366 nsew power bidirectional
flabel metal4 s 19568 2128 19888 61520 0 FreeSans 1920 90 0 0 vssd1
port 367 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 61520 0 FreeSans 1920 90 0 0 vssd1
port 367 nsew ground bidirectional
flabel metal3 s 59200 1096 60000 1216 0 FreeSans 480 0 0 0 wb_clk_i
port 368 nsew signal input
flabel metal3 s 59200 1640 60000 1760 0 FreeSans 480 0 0 0 wb_rst_i
port 369 nsew signal input
flabel metal3 s 59200 2184 60000 2304 0 FreeSans 480 0 0 0 wbs_ack_o
port 370 nsew signal tristate
flabel metal3 s 59200 4360 60000 4480 0 FreeSans 480 0 0 0 wbs_adr_i[0]
port 371 nsew signal input
flabel metal3 s 59200 20680 60000 20800 0 FreeSans 480 0 0 0 wbs_adr_i[10]
port 372 nsew signal input
flabel metal3 s 59200 22312 60000 22432 0 FreeSans 480 0 0 0 wbs_adr_i[11]
port 373 nsew signal input
flabel metal3 s 59200 23944 60000 24064 0 FreeSans 480 0 0 0 wbs_adr_i[12]
port 374 nsew signal input
flabel metal3 s 59200 25576 60000 25696 0 FreeSans 480 0 0 0 wbs_adr_i[13]
port 375 nsew signal input
flabel metal3 s 59200 27208 60000 27328 0 FreeSans 480 0 0 0 wbs_adr_i[14]
port 376 nsew signal input
flabel metal3 s 59200 28840 60000 28960 0 FreeSans 480 0 0 0 wbs_adr_i[15]
port 377 nsew signal input
flabel metal3 s 59200 30472 60000 30592 0 FreeSans 480 0 0 0 wbs_adr_i[16]
port 378 nsew signal input
flabel metal3 s 59200 32104 60000 32224 0 FreeSans 480 0 0 0 wbs_adr_i[17]
port 379 nsew signal input
flabel metal3 s 59200 33736 60000 33856 0 FreeSans 480 0 0 0 wbs_adr_i[18]
port 380 nsew signal input
flabel metal3 s 59200 35368 60000 35488 0 FreeSans 480 0 0 0 wbs_adr_i[19]
port 381 nsew signal input
flabel metal3 s 59200 5992 60000 6112 0 FreeSans 480 0 0 0 wbs_adr_i[1]
port 382 nsew signal input
flabel metal3 s 59200 37000 60000 37120 0 FreeSans 480 0 0 0 wbs_adr_i[20]
port 383 nsew signal input
flabel metal3 s 59200 38632 60000 38752 0 FreeSans 480 0 0 0 wbs_adr_i[21]
port 384 nsew signal input
flabel metal3 s 59200 40264 60000 40384 0 FreeSans 480 0 0 0 wbs_adr_i[22]
port 385 nsew signal input
flabel metal3 s 59200 41896 60000 42016 0 FreeSans 480 0 0 0 wbs_adr_i[23]
port 386 nsew signal input
flabel metal3 s 59200 43528 60000 43648 0 FreeSans 480 0 0 0 wbs_adr_i[24]
port 387 nsew signal input
flabel metal3 s 59200 45160 60000 45280 0 FreeSans 480 0 0 0 wbs_adr_i[25]
port 388 nsew signal input
flabel metal3 s 59200 46792 60000 46912 0 FreeSans 480 0 0 0 wbs_adr_i[26]
port 389 nsew signal input
flabel metal3 s 59200 48424 60000 48544 0 FreeSans 480 0 0 0 wbs_adr_i[27]
port 390 nsew signal input
flabel metal3 s 59200 50056 60000 50176 0 FreeSans 480 0 0 0 wbs_adr_i[28]
port 391 nsew signal input
flabel metal3 s 59200 51688 60000 51808 0 FreeSans 480 0 0 0 wbs_adr_i[29]
port 392 nsew signal input
flabel metal3 s 59200 7624 60000 7744 0 FreeSans 480 0 0 0 wbs_adr_i[2]
port 393 nsew signal input
flabel metal3 s 59200 53320 60000 53440 0 FreeSans 480 0 0 0 wbs_adr_i[30]
port 394 nsew signal input
flabel metal3 s 59200 54952 60000 55072 0 FreeSans 480 0 0 0 wbs_adr_i[31]
port 395 nsew signal input
flabel metal3 s 59200 9256 60000 9376 0 FreeSans 480 0 0 0 wbs_adr_i[3]
port 396 nsew signal input
flabel metal3 s 59200 10888 60000 11008 0 FreeSans 480 0 0 0 wbs_adr_i[4]
port 397 nsew signal input
flabel metal3 s 59200 12520 60000 12640 0 FreeSans 480 0 0 0 wbs_adr_i[5]
port 398 nsew signal input
flabel metal3 s 59200 14152 60000 14272 0 FreeSans 480 0 0 0 wbs_adr_i[6]
port 399 nsew signal input
flabel metal3 s 59200 15784 60000 15904 0 FreeSans 480 0 0 0 wbs_adr_i[7]
port 400 nsew signal input
flabel metal3 s 59200 17416 60000 17536 0 FreeSans 480 0 0 0 wbs_adr_i[8]
port 401 nsew signal input
flabel metal3 s 59200 19048 60000 19168 0 FreeSans 480 0 0 0 wbs_adr_i[9]
port 402 nsew signal input
flabel metal3 s 59200 2728 60000 2848 0 FreeSans 480 0 0 0 wbs_cyc_i
port 403 nsew signal input
flabel metal3 s 59200 4904 60000 5024 0 FreeSans 480 0 0 0 wbs_dat_i[0]
port 404 nsew signal input
flabel metal3 s 59200 21224 60000 21344 0 FreeSans 480 0 0 0 wbs_dat_i[10]
port 405 nsew signal input
flabel metal3 s 59200 22856 60000 22976 0 FreeSans 480 0 0 0 wbs_dat_i[11]
port 406 nsew signal input
flabel metal3 s 59200 24488 60000 24608 0 FreeSans 480 0 0 0 wbs_dat_i[12]
port 407 nsew signal input
flabel metal3 s 59200 26120 60000 26240 0 FreeSans 480 0 0 0 wbs_dat_i[13]
port 408 nsew signal input
flabel metal3 s 59200 27752 60000 27872 0 FreeSans 480 0 0 0 wbs_dat_i[14]
port 409 nsew signal input
flabel metal3 s 59200 29384 60000 29504 0 FreeSans 480 0 0 0 wbs_dat_i[15]
port 410 nsew signal input
flabel metal3 s 59200 31016 60000 31136 0 FreeSans 480 0 0 0 wbs_dat_i[16]
port 411 nsew signal input
flabel metal3 s 59200 32648 60000 32768 0 FreeSans 480 0 0 0 wbs_dat_i[17]
port 412 nsew signal input
flabel metal3 s 59200 34280 60000 34400 0 FreeSans 480 0 0 0 wbs_dat_i[18]
port 413 nsew signal input
flabel metal3 s 59200 35912 60000 36032 0 FreeSans 480 0 0 0 wbs_dat_i[19]
port 414 nsew signal input
flabel metal3 s 59200 6536 60000 6656 0 FreeSans 480 0 0 0 wbs_dat_i[1]
port 415 nsew signal input
flabel metal3 s 59200 37544 60000 37664 0 FreeSans 480 0 0 0 wbs_dat_i[20]
port 416 nsew signal input
flabel metal3 s 59200 39176 60000 39296 0 FreeSans 480 0 0 0 wbs_dat_i[21]
port 417 nsew signal input
flabel metal3 s 59200 40808 60000 40928 0 FreeSans 480 0 0 0 wbs_dat_i[22]
port 418 nsew signal input
flabel metal3 s 59200 42440 60000 42560 0 FreeSans 480 0 0 0 wbs_dat_i[23]
port 419 nsew signal input
flabel metal3 s 59200 44072 60000 44192 0 FreeSans 480 0 0 0 wbs_dat_i[24]
port 420 nsew signal input
flabel metal3 s 59200 45704 60000 45824 0 FreeSans 480 0 0 0 wbs_dat_i[25]
port 421 nsew signal input
flabel metal3 s 59200 47336 60000 47456 0 FreeSans 480 0 0 0 wbs_dat_i[26]
port 422 nsew signal input
flabel metal3 s 59200 48968 60000 49088 0 FreeSans 480 0 0 0 wbs_dat_i[27]
port 423 nsew signal input
flabel metal3 s 59200 50600 60000 50720 0 FreeSans 480 0 0 0 wbs_dat_i[28]
port 424 nsew signal input
flabel metal3 s 59200 52232 60000 52352 0 FreeSans 480 0 0 0 wbs_dat_i[29]
port 425 nsew signal input
flabel metal3 s 59200 8168 60000 8288 0 FreeSans 480 0 0 0 wbs_dat_i[2]
port 426 nsew signal input
flabel metal3 s 59200 53864 60000 53984 0 FreeSans 480 0 0 0 wbs_dat_i[30]
port 427 nsew signal input
flabel metal3 s 59200 55496 60000 55616 0 FreeSans 480 0 0 0 wbs_dat_i[31]
port 428 nsew signal input
flabel metal3 s 59200 9800 60000 9920 0 FreeSans 480 0 0 0 wbs_dat_i[3]
port 429 nsew signal input
flabel metal3 s 59200 11432 60000 11552 0 FreeSans 480 0 0 0 wbs_dat_i[4]
port 430 nsew signal input
flabel metal3 s 59200 13064 60000 13184 0 FreeSans 480 0 0 0 wbs_dat_i[5]
port 431 nsew signal input
flabel metal3 s 59200 14696 60000 14816 0 FreeSans 480 0 0 0 wbs_dat_i[6]
port 432 nsew signal input
flabel metal3 s 59200 16328 60000 16448 0 FreeSans 480 0 0 0 wbs_dat_i[7]
port 433 nsew signal input
flabel metal3 s 59200 17960 60000 18080 0 FreeSans 480 0 0 0 wbs_dat_i[8]
port 434 nsew signal input
flabel metal3 s 59200 19592 60000 19712 0 FreeSans 480 0 0 0 wbs_dat_i[9]
port 435 nsew signal input
flabel metal3 s 59200 5448 60000 5568 0 FreeSans 480 0 0 0 wbs_dat_o[0]
port 436 nsew signal tristate
flabel metal3 s 59200 21768 60000 21888 0 FreeSans 480 0 0 0 wbs_dat_o[10]
port 437 nsew signal tristate
flabel metal3 s 59200 23400 60000 23520 0 FreeSans 480 0 0 0 wbs_dat_o[11]
port 438 nsew signal tristate
flabel metal3 s 59200 25032 60000 25152 0 FreeSans 480 0 0 0 wbs_dat_o[12]
port 439 nsew signal tristate
flabel metal3 s 59200 26664 60000 26784 0 FreeSans 480 0 0 0 wbs_dat_o[13]
port 440 nsew signal tristate
flabel metal3 s 59200 28296 60000 28416 0 FreeSans 480 0 0 0 wbs_dat_o[14]
port 441 nsew signal tristate
flabel metal3 s 59200 29928 60000 30048 0 FreeSans 480 0 0 0 wbs_dat_o[15]
port 442 nsew signal tristate
flabel metal3 s 59200 31560 60000 31680 0 FreeSans 480 0 0 0 wbs_dat_o[16]
port 443 nsew signal tristate
flabel metal3 s 59200 33192 60000 33312 0 FreeSans 480 0 0 0 wbs_dat_o[17]
port 444 nsew signal tristate
flabel metal3 s 59200 34824 60000 34944 0 FreeSans 480 0 0 0 wbs_dat_o[18]
port 445 nsew signal tristate
flabel metal3 s 59200 36456 60000 36576 0 FreeSans 480 0 0 0 wbs_dat_o[19]
port 446 nsew signal tristate
flabel metal3 s 59200 7080 60000 7200 0 FreeSans 480 0 0 0 wbs_dat_o[1]
port 447 nsew signal tristate
flabel metal3 s 59200 38088 60000 38208 0 FreeSans 480 0 0 0 wbs_dat_o[20]
port 448 nsew signal tristate
flabel metal3 s 59200 39720 60000 39840 0 FreeSans 480 0 0 0 wbs_dat_o[21]
port 449 nsew signal tristate
flabel metal3 s 59200 41352 60000 41472 0 FreeSans 480 0 0 0 wbs_dat_o[22]
port 450 nsew signal tristate
flabel metal3 s 59200 42984 60000 43104 0 FreeSans 480 0 0 0 wbs_dat_o[23]
port 451 nsew signal tristate
flabel metal3 s 59200 44616 60000 44736 0 FreeSans 480 0 0 0 wbs_dat_o[24]
port 452 nsew signal tristate
flabel metal3 s 59200 46248 60000 46368 0 FreeSans 480 0 0 0 wbs_dat_o[25]
port 453 nsew signal tristate
flabel metal3 s 59200 47880 60000 48000 0 FreeSans 480 0 0 0 wbs_dat_o[26]
port 454 nsew signal tristate
flabel metal3 s 59200 49512 60000 49632 0 FreeSans 480 0 0 0 wbs_dat_o[27]
port 455 nsew signal tristate
flabel metal3 s 59200 51144 60000 51264 0 FreeSans 480 0 0 0 wbs_dat_o[28]
port 456 nsew signal tristate
flabel metal3 s 59200 52776 60000 52896 0 FreeSans 480 0 0 0 wbs_dat_o[29]
port 457 nsew signal tristate
flabel metal3 s 59200 8712 60000 8832 0 FreeSans 480 0 0 0 wbs_dat_o[2]
port 458 nsew signal tristate
flabel metal3 s 59200 54408 60000 54528 0 FreeSans 480 0 0 0 wbs_dat_o[30]
port 459 nsew signal tristate
flabel metal3 s 59200 56040 60000 56160 0 FreeSans 480 0 0 0 wbs_dat_o[31]
port 460 nsew signal tristate
flabel metal3 s 59200 10344 60000 10464 0 FreeSans 480 0 0 0 wbs_dat_o[3]
port 461 nsew signal tristate
flabel metal3 s 59200 11976 60000 12096 0 FreeSans 480 0 0 0 wbs_dat_o[4]
port 462 nsew signal tristate
flabel metal3 s 59200 13608 60000 13728 0 FreeSans 480 0 0 0 wbs_dat_o[5]
port 463 nsew signal tristate
flabel metal3 s 59200 15240 60000 15360 0 FreeSans 480 0 0 0 wbs_dat_o[6]
port 464 nsew signal tristate
flabel metal3 s 59200 16872 60000 16992 0 FreeSans 480 0 0 0 wbs_dat_o[7]
port 465 nsew signal tristate
flabel metal3 s 59200 18504 60000 18624 0 FreeSans 480 0 0 0 wbs_dat_o[8]
port 466 nsew signal tristate
flabel metal3 s 59200 20136 60000 20256 0 FreeSans 480 0 0 0 wbs_dat_o[9]
port 467 nsew signal tristate
flabel metal3 s 59200 3272 60000 3392 0 FreeSans 480 0 0 0 wbs_stb_i
port 468 nsew signal input
flabel metal3 s 59200 3816 60000 3936 0 FreeSans 480 0 0 0 wbs_we_i
port 469 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 64000
<< end >>
