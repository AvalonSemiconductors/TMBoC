magic
tech sky130B
magscale 1 2
timestamp 1683723347
<< nwell >>
rect 1066 636741 338874 637307
rect 1066 635653 338874 636219
rect 1066 634565 338874 635131
rect 1066 633477 338874 634043
rect 1066 632389 338874 632955
rect 1066 631301 338874 631867
rect 1066 630213 338874 630779
rect 1066 629125 338874 629691
rect 1066 628037 338874 628603
rect 1066 626949 338874 627515
rect 1066 625861 338874 626427
rect 1066 624773 338874 625339
rect 1066 623685 338874 624251
rect 1066 622597 338874 623163
rect 1066 621509 338874 622075
rect 1066 620421 338874 620987
rect 1066 619333 338874 619899
rect 1066 618245 338874 618811
rect 1066 617157 338874 617723
rect 1066 616069 338874 616635
rect 1066 614981 338874 615547
rect 1066 613893 338874 614459
rect 1066 612805 338874 613371
rect 1066 611717 338874 612283
rect 1066 610629 338874 611195
rect 1066 609541 338874 610107
rect 1066 608453 338874 609019
rect 1066 607365 338874 607931
rect 1066 606277 338874 606843
rect 1066 605189 338874 605755
rect 1066 604101 338874 604667
rect 1066 603013 338874 603579
rect 1066 601925 338874 602491
rect 1066 600837 338874 601403
rect 1066 599749 338874 600315
rect 1066 598661 338874 599227
rect 1066 597573 338874 598139
rect 1066 596485 338874 597051
rect 1066 595397 338874 595963
rect 1066 594309 338874 594875
rect 1066 593221 338874 593787
rect 1066 592133 338874 592699
rect 1066 591045 338874 591611
rect 1066 589957 338874 590523
rect 1066 588869 338874 589435
rect 1066 587781 338874 588347
rect 1066 586693 338874 587259
rect 1066 585605 338874 586171
rect 1066 584517 338874 585083
rect 1066 583429 338874 583995
rect 1066 582341 338874 582907
rect 1066 581253 338874 581819
rect 1066 580165 338874 580731
rect 1066 579077 338874 579643
rect 1066 577989 338874 578555
rect 1066 576901 338874 577467
rect 1066 575813 338874 576379
rect 1066 574725 338874 575291
rect 1066 573637 338874 574203
rect 1066 572549 338874 573115
rect 1066 571461 338874 572027
rect 1066 570373 338874 570939
rect 1066 569285 338874 569851
rect 1066 568197 338874 568763
rect 1066 567109 338874 567675
rect 1066 566021 338874 566587
rect 1066 564933 338874 565499
rect 1066 563845 338874 564411
rect 1066 562757 338874 563323
rect 1066 561669 338874 562235
rect 1066 560581 338874 561147
rect 1066 559493 338874 560059
rect 1066 558405 338874 558971
rect 1066 557317 338874 557883
rect 1066 556229 338874 556795
rect 1066 555141 338874 555707
rect 1066 554053 338874 554619
rect 1066 552965 338874 553531
rect 1066 551877 338874 552443
rect 1066 550789 338874 551355
rect 1066 549701 338874 550267
rect 1066 548613 338874 549179
rect 1066 547525 338874 548091
rect 1066 546437 338874 547003
rect 1066 545349 338874 545915
rect 1066 544261 338874 544827
rect 1066 543173 338874 543739
rect 1066 542085 338874 542651
rect 1066 540997 338874 541563
rect 1066 539909 338874 540475
rect 1066 538821 338874 539387
rect 1066 537733 338874 538299
rect 1066 536645 338874 537211
rect 1066 535557 338874 536123
rect 1066 534469 338874 535035
rect 1066 533381 338874 533947
rect 1066 532293 338874 532859
rect 1066 531205 338874 531771
rect 1066 530117 338874 530683
rect 1066 529029 338874 529595
rect 1066 527941 338874 528507
rect 1066 526853 338874 527419
rect 1066 525765 338874 526331
rect 1066 524677 338874 525243
rect 1066 523589 338874 524155
rect 1066 522501 338874 523067
rect 1066 521413 338874 521979
rect 1066 520325 338874 520891
rect 1066 519237 338874 519803
rect 1066 518149 338874 518715
rect 1066 517061 338874 517627
rect 1066 515973 338874 516539
rect 1066 514885 338874 515451
rect 1066 513797 338874 514363
rect 1066 512709 338874 513275
rect 1066 511621 338874 512187
rect 1066 510533 338874 511099
rect 1066 509445 338874 510011
rect 1066 508357 338874 508923
rect 1066 507269 338874 507835
rect 1066 506181 338874 506747
rect 1066 505093 338874 505659
rect 1066 504005 338874 504571
rect 1066 502917 338874 503483
rect 1066 501829 338874 502395
rect 1066 500741 338874 501307
rect 1066 499653 338874 500219
rect 1066 498565 338874 499131
rect 1066 497477 338874 498043
rect 1066 496389 338874 496955
rect 1066 495301 338874 495867
rect 1066 494213 338874 494779
rect 1066 493125 338874 493691
rect 1066 492037 338874 492603
rect 1066 490949 338874 491515
rect 1066 489861 338874 490427
rect 1066 488773 338874 489339
rect 1066 487685 338874 488251
rect 1066 486597 338874 487163
rect 1066 485509 338874 486075
rect 1066 484421 338874 484987
rect 1066 483333 338874 483899
rect 1066 482245 338874 482811
rect 1066 481157 338874 481723
rect 1066 480069 338874 480635
rect 1066 478981 338874 479547
rect 1066 477893 338874 478459
rect 1066 476805 338874 477371
rect 1066 475717 338874 476283
rect 1066 474629 338874 475195
rect 1066 473541 338874 474107
rect 1066 472453 338874 473019
rect 1066 471365 338874 471931
rect 1066 470277 338874 470843
rect 1066 469189 338874 469755
rect 1066 468101 338874 468667
rect 1066 467013 338874 467579
rect 1066 465925 338874 466491
rect 1066 464837 338874 465403
rect 1066 463749 338874 464315
rect 1066 462661 338874 463227
rect 1066 461573 338874 462139
rect 1066 460485 338874 461051
rect 1066 459397 338874 459963
rect 1066 458309 338874 458875
rect 1066 457221 338874 457787
rect 1066 456133 338874 456699
rect 1066 455045 338874 455611
rect 1066 453957 338874 454523
rect 1066 452869 338874 453435
rect 1066 451781 338874 452347
rect 1066 450693 338874 451259
rect 1066 449605 338874 450171
rect 1066 448517 338874 449083
rect 1066 447429 338874 447995
rect 1066 446341 338874 446907
rect 1066 445253 338874 445819
rect 1066 444165 338874 444731
rect 1066 443077 338874 443643
rect 1066 441989 338874 442555
rect 1066 440901 338874 441467
rect 1066 439813 338874 440379
rect 1066 438725 338874 439291
rect 1066 437637 338874 438203
rect 1066 436549 338874 437115
rect 1066 435461 338874 436027
rect 1066 434373 338874 434939
rect 1066 433285 338874 433851
rect 1066 432197 338874 432763
rect 1066 431109 338874 431675
rect 1066 430021 338874 430587
rect 1066 428933 338874 429499
rect 1066 427845 338874 428411
rect 1066 426757 338874 427323
rect 1066 425669 338874 426235
rect 1066 424581 338874 425147
rect 1066 423493 338874 424059
rect 1066 422405 338874 422971
rect 1066 421317 338874 421883
rect 1066 420229 338874 420795
rect 1066 419141 338874 419707
rect 1066 418053 338874 418619
rect 1066 416965 338874 417531
rect 1066 415877 338874 416443
rect 1066 414789 338874 415355
rect 1066 413701 338874 414267
rect 1066 412613 338874 413179
rect 1066 411525 338874 412091
rect 1066 410437 338874 411003
rect 1066 409349 338874 409915
rect 1066 408261 338874 408827
rect 1066 407173 338874 407739
rect 1066 406085 338874 406651
rect 1066 404997 338874 405563
rect 1066 403909 338874 404475
rect 1066 402821 338874 403387
rect 1066 401733 338874 402299
rect 1066 400645 338874 401211
rect 1066 399557 338874 400123
rect 1066 398469 338874 399035
rect 1066 397381 338874 397947
rect 1066 396293 338874 396859
rect 1066 395205 338874 395771
rect 1066 394117 338874 394683
rect 1066 393029 338874 393595
rect 1066 391941 338874 392507
rect 1066 390853 338874 391419
rect 1066 389765 338874 390331
rect 1066 388677 338874 389243
rect 1066 387589 338874 388155
rect 1066 386501 338874 387067
rect 1066 385413 338874 385979
rect 1066 384325 338874 384891
rect 1066 383237 338874 383803
rect 1066 382149 338874 382715
rect 1066 381061 338874 381627
rect 1066 379973 338874 380539
rect 1066 378885 338874 379451
rect 1066 377797 338874 378363
rect 1066 376709 338874 377275
rect 1066 375621 338874 376187
rect 1066 374533 338874 375099
rect 1066 373445 338874 374011
rect 1066 372357 338874 372923
rect 1066 371269 338874 371835
rect 1066 370181 338874 370747
rect 1066 369093 338874 369659
rect 1066 368005 338874 368571
rect 1066 366917 338874 367483
rect 1066 365829 338874 366395
rect 1066 364741 338874 365307
rect 1066 363653 338874 364219
rect 1066 362565 338874 363131
rect 1066 361477 338874 362043
rect 1066 360389 338874 360955
rect 1066 359301 338874 359867
rect 1066 358213 338874 358779
rect 1066 357125 338874 357691
rect 1066 356037 338874 356603
rect 1066 354949 338874 355515
rect 1066 353861 338874 354427
rect 1066 352773 338874 353339
rect 1066 351685 338874 352251
rect 1066 350597 338874 351163
rect 1066 349509 338874 350075
rect 1066 348421 338874 348987
rect 1066 347333 338874 347899
rect 1066 346245 338874 346811
rect 1066 345157 338874 345723
rect 1066 344069 338874 344635
rect 1066 342981 338874 343547
rect 1066 341893 338874 342459
rect 1066 340805 338874 341371
rect 1066 339717 338874 340283
rect 1066 338629 338874 339195
rect 1066 337541 338874 338107
rect 1066 336453 338874 337019
rect 1066 335365 338874 335931
rect 1066 334277 338874 334843
rect 1066 333189 338874 333755
rect 1066 332101 338874 332667
rect 1066 331013 338874 331579
rect 1066 329925 338874 330491
rect 1066 328837 338874 329403
rect 1066 327749 338874 328315
rect 1066 326661 338874 327227
rect 1066 325573 338874 326139
rect 1066 324485 338874 325051
rect 1066 323397 338874 323963
rect 1066 322309 338874 322875
rect 1066 321221 338874 321787
rect 1066 320133 338874 320699
rect 1066 319045 338874 319611
rect 1066 317957 338874 318523
rect 1066 316869 338874 317435
rect 1066 315781 338874 316347
rect 1066 314693 338874 315259
rect 1066 313605 338874 314171
rect 1066 312517 338874 313083
rect 1066 311429 338874 311995
rect 1066 310341 338874 310907
rect 1066 309253 338874 309819
rect 1066 308165 338874 308731
rect 1066 307077 338874 307643
rect 1066 305989 338874 306555
rect 1066 304901 338874 305467
rect 1066 303813 338874 304379
rect 1066 302725 338874 303291
rect 1066 301637 338874 302203
rect 1066 300549 338874 301115
rect 1066 299461 338874 300027
rect 1066 298373 338874 298939
rect 1066 297285 338874 297851
rect 1066 296197 338874 296763
rect 1066 295109 338874 295675
rect 1066 294021 338874 294587
rect 1066 292933 338874 293499
rect 1066 291845 338874 292411
rect 1066 290757 338874 291323
rect 1066 289669 338874 290235
rect 1066 288581 338874 289147
rect 1066 287493 338874 288059
rect 1066 286405 338874 286971
rect 1066 285317 338874 285883
rect 1066 284229 338874 284795
rect 1066 283141 338874 283707
rect 1066 282053 338874 282619
rect 1066 280965 338874 281531
rect 1066 279877 338874 280443
rect 1066 278789 338874 279355
rect 1066 277701 338874 278267
rect 1066 276613 338874 277179
rect 1066 275525 338874 276091
rect 1066 274437 338874 275003
rect 1066 273349 338874 273915
rect 1066 272261 338874 272827
rect 1066 271173 338874 271739
rect 1066 270085 338874 270651
rect 1066 268997 338874 269563
rect 1066 267909 338874 268475
rect 1066 266821 338874 267387
rect 1066 265733 338874 266299
rect 1066 264645 338874 265211
rect 1066 263557 338874 264123
rect 1066 262469 338874 263035
rect 1066 261381 338874 261947
rect 1066 260293 338874 260859
rect 1066 259205 338874 259771
rect 1066 258117 338874 258683
rect 1066 257029 338874 257595
rect 1066 255941 338874 256507
rect 1066 254853 338874 255419
rect 1066 253765 338874 254331
rect 1066 252677 338874 253243
rect 1066 251589 338874 252155
rect 1066 250501 338874 251067
rect 1066 249413 338874 249979
rect 1066 248325 338874 248891
rect 1066 247237 338874 247803
rect 1066 246149 338874 246715
rect 1066 245061 338874 245627
rect 1066 243973 338874 244539
rect 1066 242885 338874 243451
rect 1066 241797 338874 242363
rect 1066 240709 338874 241275
rect 1066 239621 338874 240187
rect 1066 238533 338874 239099
rect 1066 237445 338874 238011
rect 1066 236357 338874 236923
rect 1066 235269 338874 235835
rect 1066 234181 338874 234747
rect 1066 233093 338874 233659
rect 1066 232005 338874 232571
rect 1066 230917 338874 231483
rect 1066 229829 338874 230395
rect 1066 228741 338874 229307
rect 1066 227653 338874 228219
rect 1066 226565 338874 227131
rect 1066 225477 338874 226043
rect 1066 224389 338874 224955
rect 1066 223301 338874 223867
rect 1066 222213 338874 222779
rect 1066 221125 338874 221691
rect 1066 220037 338874 220603
rect 1066 218949 338874 219515
rect 1066 217861 338874 218427
rect 1066 216773 338874 217339
rect 1066 215685 338874 216251
rect 1066 214597 338874 215163
rect 1066 213509 338874 214075
rect 1066 212421 338874 212987
rect 1066 211333 338874 211899
rect 1066 210245 338874 210811
rect 1066 209157 338874 209723
rect 1066 208069 338874 208635
rect 1066 206981 338874 207547
rect 1066 205893 338874 206459
rect 1066 204805 338874 205371
rect 1066 203717 338874 204283
rect 1066 202629 338874 203195
rect 1066 201541 338874 202107
rect 1066 200453 338874 201019
rect 1066 199365 338874 199931
rect 1066 198277 338874 198843
rect 1066 197189 338874 197755
rect 1066 196101 338874 196667
rect 1066 195013 338874 195579
rect 1066 193925 338874 194491
rect 1066 192837 338874 193403
rect 1066 191749 338874 192315
rect 1066 190661 338874 191227
rect 1066 189573 338874 190139
rect 1066 188485 338874 189051
rect 1066 187397 338874 187963
rect 1066 186309 338874 186875
rect 1066 185221 338874 185787
rect 1066 184133 338874 184699
rect 1066 183045 338874 183611
rect 1066 181957 338874 182523
rect 1066 180869 338874 181435
rect 1066 179781 338874 180347
rect 1066 178693 338874 179259
rect 1066 177605 338874 178171
rect 1066 176517 338874 177083
rect 1066 175429 338874 175995
rect 1066 174341 338874 174907
rect 1066 173253 338874 173819
rect 1066 172165 338874 172731
rect 1066 171077 338874 171643
rect 1066 169989 338874 170555
rect 1066 168901 338874 169467
rect 1066 167813 338874 168379
rect 1066 166725 338874 167291
rect 1066 165637 338874 166203
rect 1066 164549 338874 165115
rect 1066 163461 338874 164027
rect 1066 162373 338874 162939
rect 1066 161285 338874 161851
rect 1066 160197 338874 160763
rect 1066 159109 338874 159675
rect 1066 158021 338874 158587
rect 1066 156933 338874 157499
rect 1066 155845 338874 156411
rect 1066 154757 338874 155323
rect 1066 153669 338874 154235
rect 1066 152581 338874 153147
rect 1066 151493 338874 152059
rect 1066 150405 338874 150971
rect 1066 149317 338874 149883
rect 1066 148229 338874 148795
rect 1066 147141 338874 147707
rect 1066 146053 338874 146619
rect 1066 144965 338874 145531
rect 1066 143877 338874 144443
rect 1066 142789 338874 143355
rect 1066 141701 338874 142267
rect 1066 140613 338874 141179
rect 1066 139525 338874 140091
rect 1066 138437 338874 139003
rect 1066 137349 338874 137915
rect 1066 136261 338874 136827
rect 1066 135173 338874 135739
rect 1066 134085 338874 134651
rect 1066 132997 338874 133563
rect 1066 131909 338874 132475
rect 1066 130821 338874 131387
rect 1066 129733 338874 130299
rect 1066 128645 338874 129211
rect 1066 127557 338874 128123
rect 1066 126469 338874 127035
rect 1066 125381 338874 125947
rect 1066 124293 338874 124859
rect 1066 123205 338874 123771
rect 1066 122117 338874 122683
rect 1066 121029 338874 121595
rect 1066 119941 338874 120507
rect 1066 118853 338874 119419
rect 1066 117765 338874 118331
rect 1066 116677 338874 117243
rect 1066 115589 338874 116155
rect 1066 114501 338874 115067
rect 1066 113413 338874 113979
rect 1066 112325 338874 112891
rect 1066 111237 338874 111803
rect 1066 110149 338874 110715
rect 1066 109061 338874 109627
rect 1066 107973 338874 108539
rect 1066 106885 338874 107451
rect 1066 105797 338874 106363
rect 1066 104709 338874 105275
rect 1066 103621 338874 104187
rect 1066 102533 338874 103099
rect 1066 101445 338874 102011
rect 1066 100357 338874 100923
rect 1066 99269 338874 99835
rect 1066 98181 338874 98747
rect 1066 97093 338874 97659
rect 1066 96005 338874 96571
rect 1066 94917 338874 95483
rect 1066 93829 338874 94395
rect 1066 92741 338874 93307
rect 1066 91653 338874 92219
rect 1066 90565 338874 91131
rect 1066 89477 338874 90043
rect 1066 88389 338874 88955
rect 1066 87301 338874 87867
rect 1066 86213 338874 86779
rect 1066 85125 338874 85691
rect 1066 84037 338874 84603
rect 1066 82949 338874 83515
rect 1066 81861 338874 82427
rect 1066 80773 338874 81339
rect 1066 79685 338874 80251
rect 1066 78597 338874 79163
rect 1066 77509 338874 78075
rect 1066 76421 338874 76987
rect 1066 75333 338874 75899
rect 1066 74245 338874 74811
rect 1066 73157 338874 73723
rect 1066 72069 338874 72635
rect 1066 70981 338874 71547
rect 1066 69893 338874 70459
rect 1066 68805 338874 69371
rect 1066 67717 338874 68283
rect 1066 66629 338874 67195
rect 1066 65541 338874 66107
rect 1066 64453 338874 65019
rect 1066 63365 338874 63931
rect 1066 62277 338874 62843
rect 1066 61189 338874 61755
rect 1066 60101 338874 60667
rect 1066 59013 338874 59579
rect 1066 57925 338874 58491
rect 1066 56837 338874 57403
rect 1066 55749 338874 56315
rect 1066 54661 338874 55227
rect 1066 53573 338874 54139
rect 1066 52485 338874 53051
rect 1066 51397 338874 51963
rect 1066 50309 338874 50875
rect 1066 49221 338874 49787
rect 1066 48133 338874 48699
rect 1066 47045 338874 47611
rect 1066 45957 338874 46523
rect 1066 44869 338874 45435
rect 1066 43781 338874 44347
rect 1066 42693 338874 43259
rect 1066 41605 338874 42171
rect 1066 40517 338874 41083
rect 1066 39429 338874 39995
rect 1066 38341 338874 38907
rect 1066 37253 338874 37819
rect 1066 36165 338874 36731
rect 1066 35077 338874 35643
rect 1066 33989 338874 34555
rect 1066 32901 338874 33467
rect 1066 31813 338874 32379
rect 1066 30725 338874 31291
rect 1066 29637 338874 30203
rect 1066 28549 338874 29115
rect 1066 27461 338874 28027
rect 1066 26373 338874 26939
rect 1066 25285 338874 25851
rect 1066 24197 338874 24763
rect 1066 23109 338874 23675
rect 1066 22021 338874 22587
rect 1066 20933 338874 21499
rect 1066 19845 338874 20411
rect 1066 18757 338874 19323
rect 1066 17669 338874 18235
rect 1066 16581 338874 17147
rect 1066 15493 338874 16059
rect 1066 14405 338874 14971
rect 1066 13317 338874 13883
rect 1066 12229 338874 12795
rect 1066 11141 338874 11707
rect 1066 10053 338874 10619
rect 1066 8965 338874 9531
rect 1066 7877 338874 8443
rect 1066 6789 338874 7355
rect 1066 5701 338874 6267
rect 1066 4613 338874 5179
rect 1066 3525 338874 4091
rect 1066 2437 338874 3003
<< obsli1 >>
rect 1104 2159 338836 637585
<< obsm1 >>
rect 1104 2128 339374 637616
<< obsm2 >>
rect 1584 2139 339368 637605
<< metal3 >>
rect 339200 633904 340000 634024
rect 339200 622888 340000 623008
rect 339200 611872 340000 611992
rect 339200 600856 340000 600976
rect 339200 589840 340000 589960
rect 339200 578824 340000 578944
rect 339200 567808 340000 567928
rect 339200 556792 340000 556912
rect 339200 545776 340000 545896
rect 339200 534760 340000 534880
rect 339200 523744 340000 523864
rect 339200 512728 340000 512848
rect 339200 501712 340000 501832
rect 339200 490696 340000 490816
rect 339200 479680 340000 479800
rect 339200 468664 340000 468784
rect 339200 457648 340000 457768
rect 339200 446632 340000 446752
rect 339200 435616 340000 435736
rect 339200 424600 340000 424720
rect 339200 413584 340000 413704
rect 339200 402568 340000 402688
rect 339200 391552 340000 391672
rect 339200 380536 340000 380656
rect 339200 369520 340000 369640
rect 339200 358504 340000 358624
rect 339200 347488 340000 347608
rect 339200 336472 340000 336592
rect 339200 325456 340000 325576
rect 339200 314440 340000 314560
rect 339200 303424 340000 303544
rect 339200 292408 340000 292528
rect 339200 281392 340000 281512
rect 339200 270376 340000 270496
rect 339200 259360 340000 259480
rect 339200 248344 340000 248464
rect 339200 237328 340000 237448
rect 339200 226312 340000 226432
rect 339200 215296 340000 215416
rect 339200 204280 340000 204400
rect 339200 193264 340000 193384
rect 339200 182248 340000 182368
rect 339200 171232 340000 171352
rect 339200 160216 340000 160336
rect 339200 149200 340000 149320
rect 339200 138184 340000 138304
rect 339200 127168 340000 127288
rect 339200 116152 340000 116272
rect 339200 105136 340000 105256
rect 339200 94120 340000 94240
rect 339200 83104 340000 83224
rect 339200 72088 340000 72208
rect 339200 61072 340000 61192
rect 339200 50056 340000 50176
rect 339200 39040 340000 39160
rect 339200 28024 340000 28144
rect 339200 17008 340000 17128
rect 339200 5992 340000 6112
<< obsm3 >>
rect 4210 634104 339200 637601
rect 4210 633824 339120 634104
rect 4210 623088 339200 633824
rect 4210 622808 339120 623088
rect 4210 612072 339200 622808
rect 4210 611792 339120 612072
rect 4210 601056 339200 611792
rect 4210 600776 339120 601056
rect 4210 590040 339200 600776
rect 4210 589760 339120 590040
rect 4210 579024 339200 589760
rect 4210 578744 339120 579024
rect 4210 568008 339200 578744
rect 4210 567728 339120 568008
rect 4210 556992 339200 567728
rect 4210 556712 339120 556992
rect 4210 545976 339200 556712
rect 4210 545696 339120 545976
rect 4210 534960 339200 545696
rect 4210 534680 339120 534960
rect 4210 523944 339200 534680
rect 4210 523664 339120 523944
rect 4210 512928 339200 523664
rect 4210 512648 339120 512928
rect 4210 501912 339200 512648
rect 4210 501632 339120 501912
rect 4210 490896 339200 501632
rect 4210 490616 339120 490896
rect 4210 479880 339200 490616
rect 4210 479600 339120 479880
rect 4210 468864 339200 479600
rect 4210 468584 339120 468864
rect 4210 457848 339200 468584
rect 4210 457568 339120 457848
rect 4210 446832 339200 457568
rect 4210 446552 339120 446832
rect 4210 435816 339200 446552
rect 4210 435536 339120 435816
rect 4210 424800 339200 435536
rect 4210 424520 339120 424800
rect 4210 413784 339200 424520
rect 4210 413504 339120 413784
rect 4210 402768 339200 413504
rect 4210 402488 339120 402768
rect 4210 391752 339200 402488
rect 4210 391472 339120 391752
rect 4210 380736 339200 391472
rect 4210 380456 339120 380736
rect 4210 369720 339200 380456
rect 4210 369440 339120 369720
rect 4210 358704 339200 369440
rect 4210 358424 339120 358704
rect 4210 347688 339200 358424
rect 4210 347408 339120 347688
rect 4210 336672 339200 347408
rect 4210 336392 339120 336672
rect 4210 325656 339200 336392
rect 4210 325376 339120 325656
rect 4210 314640 339200 325376
rect 4210 314360 339120 314640
rect 4210 303624 339200 314360
rect 4210 303344 339120 303624
rect 4210 292608 339200 303344
rect 4210 292328 339120 292608
rect 4210 281592 339200 292328
rect 4210 281312 339120 281592
rect 4210 270576 339200 281312
rect 4210 270296 339120 270576
rect 4210 259560 339200 270296
rect 4210 259280 339120 259560
rect 4210 248544 339200 259280
rect 4210 248264 339120 248544
rect 4210 237528 339200 248264
rect 4210 237248 339120 237528
rect 4210 226512 339200 237248
rect 4210 226232 339120 226512
rect 4210 215496 339200 226232
rect 4210 215216 339120 215496
rect 4210 204480 339200 215216
rect 4210 204200 339120 204480
rect 4210 193464 339200 204200
rect 4210 193184 339120 193464
rect 4210 182448 339200 193184
rect 4210 182168 339120 182448
rect 4210 171432 339200 182168
rect 4210 171152 339120 171432
rect 4210 160416 339200 171152
rect 4210 160136 339120 160416
rect 4210 149400 339200 160136
rect 4210 149120 339120 149400
rect 4210 138384 339200 149120
rect 4210 138104 339120 138384
rect 4210 127368 339200 138104
rect 4210 127088 339120 127368
rect 4210 116352 339200 127088
rect 4210 116072 339120 116352
rect 4210 105336 339200 116072
rect 4210 105056 339120 105336
rect 4210 94320 339200 105056
rect 4210 94040 339120 94320
rect 4210 83304 339200 94040
rect 4210 83024 339120 83304
rect 4210 72288 339200 83024
rect 4210 72008 339120 72288
rect 4210 61272 339200 72008
rect 4210 60992 339120 61272
rect 4210 50256 339200 60992
rect 4210 49976 339120 50256
rect 4210 39240 339200 49976
rect 4210 38960 339120 39240
rect 4210 28224 339200 38960
rect 4210 27944 339120 28224
rect 4210 17208 339200 27944
rect 4210 16928 339120 17208
rect 4210 6192 339200 16928
rect 4210 5912 339120 6192
rect 4210 2143 339200 5912
<< metal4 >>
rect 4208 2128 4528 637616
rect 19568 2128 19888 637616
rect 34928 2128 35248 637616
rect 50288 2128 50608 637616
rect 65648 2128 65968 637616
rect 81008 2128 81328 637616
rect 96368 2128 96688 637616
rect 111728 2128 112048 637616
rect 127088 2128 127408 637616
rect 142448 2128 142768 637616
rect 157808 2128 158128 637616
rect 173168 2128 173488 637616
rect 188528 2128 188848 637616
rect 203888 2128 204208 637616
rect 219248 2128 219568 637616
rect 234608 2128 234928 637616
rect 249968 2128 250288 637616
rect 265328 2128 265648 637616
rect 280688 2128 281008 637616
rect 296048 2128 296368 637616
rect 311408 2128 311728 637616
rect 326768 2128 327088 637616
<< obsm4 >>
rect 12203 6427 19488 627333
rect 19968 6427 34848 627333
rect 35328 6427 50208 627333
rect 50688 6427 65568 627333
rect 66048 6427 80928 627333
rect 81408 6427 96288 627333
rect 96768 6427 111648 627333
rect 112128 6427 127008 627333
rect 127488 6427 142368 627333
rect 142848 6427 157728 627333
rect 158208 6427 173088 627333
rect 173568 6427 188448 627333
rect 188928 6427 203808 627333
rect 204288 6427 219168 627333
rect 219648 6427 234528 627333
rect 235008 6427 249888 627333
rect 250368 6427 265248 627333
rect 265728 6427 280608 627333
rect 281088 6427 295968 627333
rect 296448 6427 311328 627333
rect 311808 6427 326688 627333
rect 327168 6427 336845 627333
<< labels >>
rlabel metal3 s 339200 303424 340000 303544 6 clk
port 1 nsew signal input
rlabel metal3 s 339200 5992 340000 6112 6 io_in[0]
port 2 nsew signal input
rlabel metal3 s 339200 116152 340000 116272 6 io_in[10]
port 3 nsew signal input
rlabel metal3 s 339200 127168 340000 127288 6 io_in[11]
port 4 nsew signal input
rlabel metal3 s 339200 138184 340000 138304 6 io_in[12]
port 5 nsew signal input
rlabel metal3 s 339200 149200 340000 149320 6 io_in[13]
port 6 nsew signal input
rlabel metal3 s 339200 160216 340000 160336 6 io_in[14]
port 7 nsew signal input
rlabel metal3 s 339200 171232 340000 171352 6 io_in[15]
port 8 nsew signal input
rlabel metal3 s 339200 182248 340000 182368 6 io_in[16]
port 9 nsew signal input
rlabel metal3 s 339200 193264 340000 193384 6 io_in[17]
port 10 nsew signal input
rlabel metal3 s 339200 204280 340000 204400 6 io_in[18]
port 11 nsew signal input
rlabel metal3 s 339200 215296 340000 215416 6 io_in[19]
port 12 nsew signal input
rlabel metal3 s 339200 17008 340000 17128 6 io_in[1]
port 13 nsew signal input
rlabel metal3 s 339200 226312 340000 226432 6 io_in[20]
port 14 nsew signal input
rlabel metal3 s 339200 237328 340000 237448 6 io_in[21]
port 15 nsew signal input
rlabel metal3 s 339200 248344 340000 248464 6 io_in[22]
port 16 nsew signal input
rlabel metal3 s 339200 259360 340000 259480 6 io_in[23]
port 17 nsew signal input
rlabel metal3 s 339200 270376 340000 270496 6 io_in[24]
port 18 nsew signal input
rlabel metal3 s 339200 281392 340000 281512 6 io_in[25]
port 19 nsew signal input
rlabel metal3 s 339200 292408 340000 292528 6 io_in[26]
port 20 nsew signal input
rlabel metal3 s 339200 28024 340000 28144 6 io_in[2]
port 21 nsew signal input
rlabel metal3 s 339200 39040 340000 39160 6 io_in[3]
port 22 nsew signal input
rlabel metal3 s 339200 50056 340000 50176 6 io_in[4]
port 23 nsew signal input
rlabel metal3 s 339200 61072 340000 61192 6 io_in[5]
port 24 nsew signal input
rlabel metal3 s 339200 72088 340000 72208 6 io_in[6]
port 25 nsew signal input
rlabel metal3 s 339200 83104 340000 83224 6 io_in[7]
port 26 nsew signal input
rlabel metal3 s 339200 94120 340000 94240 6 io_in[8]
port 27 nsew signal input
rlabel metal3 s 339200 105136 340000 105256 6 io_in[9]
port 28 nsew signal input
rlabel metal3 s 339200 633904 340000 634024 6 io_oeb
port 29 nsew signal output
rlabel metal3 s 339200 325456 340000 325576 6 io_out[0]
port 30 nsew signal output
rlabel metal3 s 339200 435616 340000 435736 6 io_out[10]
port 31 nsew signal output
rlabel metal3 s 339200 446632 340000 446752 6 io_out[11]
port 32 nsew signal output
rlabel metal3 s 339200 457648 340000 457768 6 io_out[12]
port 33 nsew signal output
rlabel metal3 s 339200 468664 340000 468784 6 io_out[13]
port 34 nsew signal output
rlabel metal3 s 339200 479680 340000 479800 6 io_out[14]
port 35 nsew signal output
rlabel metal3 s 339200 490696 340000 490816 6 io_out[15]
port 36 nsew signal output
rlabel metal3 s 339200 501712 340000 501832 6 io_out[16]
port 37 nsew signal output
rlabel metal3 s 339200 512728 340000 512848 6 io_out[17]
port 38 nsew signal output
rlabel metal3 s 339200 523744 340000 523864 6 io_out[18]
port 39 nsew signal output
rlabel metal3 s 339200 534760 340000 534880 6 io_out[19]
port 40 nsew signal output
rlabel metal3 s 339200 336472 340000 336592 6 io_out[1]
port 41 nsew signal output
rlabel metal3 s 339200 545776 340000 545896 6 io_out[20]
port 42 nsew signal output
rlabel metal3 s 339200 556792 340000 556912 6 io_out[21]
port 43 nsew signal output
rlabel metal3 s 339200 567808 340000 567928 6 io_out[22]
port 44 nsew signal output
rlabel metal3 s 339200 578824 340000 578944 6 io_out[23]
port 45 nsew signal output
rlabel metal3 s 339200 589840 340000 589960 6 io_out[24]
port 46 nsew signal output
rlabel metal3 s 339200 600856 340000 600976 6 io_out[25]
port 47 nsew signal output
rlabel metal3 s 339200 611872 340000 611992 6 io_out[26]
port 48 nsew signal output
rlabel metal3 s 339200 622888 340000 623008 6 io_out[27]
port 49 nsew signal output
rlabel metal3 s 339200 347488 340000 347608 6 io_out[2]
port 50 nsew signal output
rlabel metal3 s 339200 358504 340000 358624 6 io_out[3]
port 51 nsew signal output
rlabel metal3 s 339200 369520 340000 369640 6 io_out[4]
port 52 nsew signal output
rlabel metal3 s 339200 380536 340000 380656 6 io_out[5]
port 53 nsew signal output
rlabel metal3 s 339200 391552 340000 391672 6 io_out[6]
port 54 nsew signal output
rlabel metal3 s 339200 402568 340000 402688 6 io_out[7]
port 55 nsew signal output
rlabel metal3 s 339200 413584 340000 413704 6 io_out[8]
port 56 nsew signal output
rlabel metal3 s 339200 424600 340000 424720 6 io_out[9]
port 57 nsew signal output
rlabel metal3 s 339200 314440 340000 314560 6 rst
port 58 nsew signal input
rlabel metal4 s 4208 2128 4528 637616 6 vccd1
port 59 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 637616 6 vccd1
port 59 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 637616 6 vccd1
port 59 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 637616 6 vccd1
port 59 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 637616 6 vccd1
port 59 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 637616 6 vccd1
port 59 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 637616 6 vccd1
port 59 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 637616 6 vccd1
port 59 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 637616 6 vccd1
port 59 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 637616 6 vccd1
port 59 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 637616 6 vccd1
port 59 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 637616 6 vssd1
port 60 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 637616 6 vssd1
port 60 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 637616 6 vssd1
port 60 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 637616 6 vssd1
port 60 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 637616 6 vssd1
port 60 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 637616 6 vssd1
port 60 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 637616 6 vssd1
port 60 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 637616 6 vssd1
port 60 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 637616 6 vssd1
port 60 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 637616 6 vssd1
port 60 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 637616 6 vssd1
port 60 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 340000 640000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 264297370
string GDS_FILE /media/lucah/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/AS512512512/runs/23_05_10_09_08/results/signoff/wrapped_as512512512.magic.gds
string GDS_START 1780936
<< end >>

