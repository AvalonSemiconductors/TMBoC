VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_6502
  CLASS BLOCK ;
  FOREIGN wrapped_6502 ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 200.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 196.000 174.710 200.000 ;
    END
  END clk
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 196.000 9.110 200.000 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 196.000 25.670 200.000 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 196.000 42.230 200.000 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 196.000 58.790 200.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 196.000 75.350 200.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 196.000 91.910 200.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 196.000 108.470 200.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 196.000 125.030 200.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 196.000 141.590 200.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 196.000 158.150 200.000 ;
    END
  END io_in[9]
  PIN io_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 191.120 200.000 191.720 ;
    END
  END io_oeb
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 7.520 200.000 8.120 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 75.520 200.000 76.120 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 82.320 200.000 82.920 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 89.120 200.000 89.720 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 95.920 200.000 96.520 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 102.720 200.000 103.320 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 109.520 200.000 110.120 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 116.320 200.000 116.920 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 123.120 200.000 123.720 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 129.920 200.000 130.520 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 136.720 200.000 137.320 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 14.320 200.000 14.920 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 143.520 200.000 144.120 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 150.320 200.000 150.920 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 157.120 200.000 157.720 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 163.920 200.000 164.520 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 170.720 200.000 171.320 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 177.520 200.000 178.120 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 184.320 200.000 184.920 ;
    END
  END io_out[26]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 21.120 200.000 21.720 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 27.920 200.000 28.520 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 34.720 200.000 35.320 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 41.520 200.000 42.120 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 48.320 200.000 48.920 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 55.120 200.000 55.720 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 61.920 200.000 62.520 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 68.720 200.000 69.320 ;
    END
  END io_out[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 196.000 191.270 200.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 187.920 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 186.265 194.310 187.870 ;
        RECT 5.330 180.825 194.310 183.655 ;
        RECT 5.330 175.385 194.310 178.215 ;
        RECT 5.330 169.945 194.310 172.775 ;
        RECT 5.330 164.505 194.310 167.335 ;
        RECT 5.330 159.065 194.310 161.895 ;
        RECT 5.330 153.625 194.310 156.455 ;
        RECT 5.330 148.185 194.310 151.015 ;
        RECT 5.330 142.745 194.310 145.575 ;
        RECT 5.330 137.305 194.310 140.135 ;
        RECT 5.330 131.865 194.310 134.695 ;
        RECT 5.330 126.425 194.310 129.255 ;
        RECT 5.330 120.985 194.310 123.815 ;
        RECT 5.330 115.545 194.310 118.375 ;
        RECT 5.330 110.105 194.310 112.935 ;
        RECT 5.330 104.665 194.310 107.495 ;
        RECT 5.330 99.225 194.310 102.055 ;
        RECT 5.330 93.785 194.310 96.615 ;
        RECT 5.330 88.345 194.310 91.175 ;
        RECT 5.330 82.905 194.310 85.735 ;
        RECT 5.330 77.465 194.310 80.295 ;
        RECT 5.330 72.025 194.310 74.855 ;
        RECT 5.330 66.585 194.310 69.415 ;
        RECT 5.330 61.145 194.310 63.975 ;
        RECT 5.330 55.705 194.310 58.535 ;
        RECT 5.330 50.265 194.310 53.095 ;
        RECT 5.330 44.825 194.310 47.655 ;
        RECT 5.330 39.385 194.310 42.215 ;
        RECT 5.330 33.945 194.310 36.775 ;
        RECT 5.330 28.505 194.310 31.335 ;
        RECT 5.330 23.065 194.310 25.895 ;
        RECT 5.330 17.625 194.310 20.455 ;
        RECT 5.330 12.185 194.310 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 194.120 187.765 ;
      LAYER met1 ;
        RECT 5.520 10.640 198.190 196.480 ;
      LAYER met2 ;
        RECT 8.370 195.720 8.550 197.045 ;
        RECT 9.390 195.720 25.110 197.045 ;
        RECT 25.950 195.720 41.670 197.045 ;
        RECT 42.510 195.720 58.230 197.045 ;
        RECT 59.070 195.720 74.790 197.045 ;
        RECT 75.630 195.720 91.350 197.045 ;
        RECT 92.190 195.720 107.910 197.045 ;
        RECT 108.750 195.720 124.470 197.045 ;
        RECT 125.310 195.720 141.030 197.045 ;
        RECT 141.870 195.720 157.590 197.045 ;
        RECT 158.430 195.720 174.150 197.045 ;
        RECT 174.990 195.720 190.710 197.045 ;
        RECT 191.550 195.720 198.170 197.045 ;
        RECT 8.370 7.635 198.170 195.720 ;
      LAYER met3 ;
        RECT 8.345 192.120 198.195 197.025 ;
        RECT 8.345 190.720 195.600 192.120 ;
        RECT 8.345 185.320 198.195 190.720 ;
        RECT 8.345 183.920 195.600 185.320 ;
        RECT 8.345 178.520 198.195 183.920 ;
        RECT 8.345 177.120 195.600 178.520 ;
        RECT 8.345 171.720 198.195 177.120 ;
        RECT 8.345 170.320 195.600 171.720 ;
        RECT 8.345 164.920 198.195 170.320 ;
        RECT 8.345 163.520 195.600 164.920 ;
        RECT 8.345 158.120 198.195 163.520 ;
        RECT 8.345 156.720 195.600 158.120 ;
        RECT 8.345 151.320 198.195 156.720 ;
        RECT 8.345 149.920 195.600 151.320 ;
        RECT 8.345 144.520 198.195 149.920 ;
        RECT 8.345 143.120 195.600 144.520 ;
        RECT 8.345 137.720 198.195 143.120 ;
        RECT 8.345 136.320 195.600 137.720 ;
        RECT 8.345 130.920 198.195 136.320 ;
        RECT 8.345 129.520 195.600 130.920 ;
        RECT 8.345 124.120 198.195 129.520 ;
        RECT 8.345 122.720 195.600 124.120 ;
        RECT 8.345 117.320 198.195 122.720 ;
        RECT 8.345 115.920 195.600 117.320 ;
        RECT 8.345 110.520 198.195 115.920 ;
        RECT 8.345 109.120 195.600 110.520 ;
        RECT 8.345 103.720 198.195 109.120 ;
        RECT 8.345 102.320 195.600 103.720 ;
        RECT 8.345 96.920 198.195 102.320 ;
        RECT 8.345 95.520 195.600 96.920 ;
        RECT 8.345 90.120 198.195 95.520 ;
        RECT 8.345 88.720 195.600 90.120 ;
        RECT 8.345 83.320 198.195 88.720 ;
        RECT 8.345 81.920 195.600 83.320 ;
        RECT 8.345 76.520 198.195 81.920 ;
        RECT 8.345 75.120 195.600 76.520 ;
        RECT 8.345 69.720 198.195 75.120 ;
        RECT 8.345 68.320 195.600 69.720 ;
        RECT 8.345 62.920 198.195 68.320 ;
        RECT 8.345 61.520 195.600 62.920 ;
        RECT 8.345 56.120 198.195 61.520 ;
        RECT 8.345 54.720 195.600 56.120 ;
        RECT 8.345 49.320 198.195 54.720 ;
        RECT 8.345 47.920 195.600 49.320 ;
        RECT 8.345 42.520 198.195 47.920 ;
        RECT 8.345 41.120 195.600 42.520 ;
        RECT 8.345 35.720 198.195 41.120 ;
        RECT 8.345 34.320 195.600 35.720 ;
        RECT 8.345 28.920 198.195 34.320 ;
        RECT 8.345 27.520 195.600 28.920 ;
        RECT 8.345 22.120 198.195 27.520 ;
        RECT 8.345 20.720 195.600 22.120 ;
        RECT 8.345 15.320 198.195 20.720 ;
        RECT 8.345 13.920 195.600 15.320 ;
        RECT 8.345 8.520 198.195 13.920 ;
        RECT 8.345 7.655 195.600 8.520 ;
      LAYER met4 ;
        RECT 24.215 188.320 185.545 197.025 ;
        RECT 24.215 12.415 97.440 188.320 ;
        RECT 99.840 12.415 174.240 188.320 ;
        RECT 176.640 12.415 185.545 188.320 ;
  END
END wrapped_6502
END LIBRARY

