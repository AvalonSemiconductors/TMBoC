magic
tech sky130B
magscale 1 2
timestamp 1675976272
<< obsli1 >>
rect 1104 2159 22816 21777
<< obsm1 >>
rect 1104 2128 22976 21808
<< obsm2 >>
rect 1584 2139 22970 21797
<< metal3 >>
rect 0 19668 800 19908
rect 0 11780 800 12020
rect 0 3892 800 4132
<< obsm3 >>
rect 800 19988 22974 21793
rect 880 19588 22974 19988
rect 800 12100 22974 19588
rect 880 11700 22974 12100
rect 800 4212 22974 11700
rect 880 3812 22974 4212
rect 800 2143 22974 3812
<< metal4 >>
rect 3658 2128 3978 21808
rect 6372 2128 6692 21808
rect 9086 2128 9406 21808
rect 11800 2128 12120 21808
rect 14514 2128 14834 21808
rect 17228 2128 17548 21808
rect 19942 2128 20262 21808
rect 22656 2128 22976 21808
<< obsm4 >>
rect 15147 3979 17148 10573
rect 17628 3979 19629 10573
<< labels >>
rlabel metal3 s 0 19668 800 19908 6 OP
port 1 nsew signal output
rlabel metal3 s 0 3892 800 4132 6 clk
port 2 nsew signal input
rlabel metal3 s 0 11780 800 12020 6 rst
port 3 nsew signal input
rlabel metal4 s 3658 2128 3978 21808 6 vccd1
port 4 nsew power bidirectional
rlabel metal4 s 9086 2128 9406 21808 6 vccd1
port 4 nsew power bidirectional
rlabel metal4 s 14514 2128 14834 21808 6 vccd1
port 4 nsew power bidirectional
rlabel metal4 s 19942 2128 20262 21808 6 vccd1
port 4 nsew power bidirectional
rlabel metal4 s 6372 2128 6692 21808 6 vssd1
port 5 nsew ground bidirectional
rlabel metal4 s 11800 2128 12120 21808 6 vssd1
port 5 nsew ground bidirectional
rlabel metal4 s 17228 2128 17548 21808 6 vssd1
port 5 nsew ground bidirectional
rlabel metal4 s 22656 2128 22976 21808 6 vssd1
port 5 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 24000 24000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1275808
string GDS_FILE /run/media/tholin/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/TunePlayer/runs/23_02_09_21_56/results/signoff/tune_player.magic.gds
string GDS_START 416620
<< end >>

