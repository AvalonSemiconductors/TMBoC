magic
tech sky130B
magscale 1 2
timestamp 1679913442
<< nwell >>
rect 1066 617157 358930 617478
rect 1066 616069 358930 616635
rect 1066 614981 358930 615547
rect 1066 613893 358930 614459
rect 1066 612805 358930 613371
rect 1066 611717 358930 612283
rect 1066 610629 358930 611195
rect 1066 609541 358930 610107
rect 1066 608453 358930 609019
rect 1066 607365 358930 607931
rect 1066 606277 358930 606843
rect 1066 605189 358930 605755
rect 1066 604101 358930 604667
rect 1066 603013 358930 603579
rect 1066 601925 358930 602491
rect 1066 600837 358930 601403
rect 1066 599749 358930 600315
rect 1066 598661 358930 599227
rect 1066 597573 358930 598139
rect 1066 596485 358930 597051
rect 1066 595397 358930 595963
rect 1066 594309 358930 594875
rect 1066 593221 358930 593787
rect 1066 592133 358930 592699
rect 1066 591045 358930 591611
rect 1066 589957 358930 590523
rect 1066 588869 358930 589435
rect 1066 587781 358930 588347
rect 1066 586693 358930 587259
rect 1066 585605 358930 586171
rect 1066 584517 358930 585083
rect 1066 583429 358930 583995
rect 1066 582341 358930 582907
rect 1066 581253 358930 581819
rect 1066 580165 358930 580731
rect 1066 579077 358930 579643
rect 1066 577989 358930 578555
rect 1066 576901 358930 577467
rect 1066 575813 358930 576379
rect 1066 574725 358930 575291
rect 1066 573637 358930 574203
rect 1066 572549 358930 573115
rect 1066 571461 358930 572027
rect 1066 570373 358930 570939
rect 1066 569285 358930 569851
rect 1066 568197 358930 568763
rect 1066 567109 358930 567675
rect 1066 566021 358930 566587
rect 1066 564933 358930 565499
rect 1066 563845 358930 564411
rect 1066 562757 358930 563323
rect 1066 561669 358930 562235
rect 1066 560581 358930 561147
rect 1066 559493 358930 560059
rect 1066 558405 358930 558971
rect 1066 557317 358930 557883
rect 1066 556229 358930 556795
rect 1066 555141 358930 555707
rect 1066 554053 358930 554619
rect 1066 552965 358930 553531
rect 1066 551877 358930 552443
rect 1066 550789 358930 551355
rect 1066 549701 358930 550267
rect 1066 548613 358930 549179
rect 1066 547525 358930 548091
rect 1066 546437 358930 547003
rect 1066 545349 358930 545915
rect 1066 544261 358930 544827
rect 1066 543173 358930 543739
rect 1066 542085 358930 542651
rect 1066 540997 358930 541563
rect 1066 539909 358930 540475
rect 1066 538821 358930 539387
rect 1066 537733 358930 538299
rect 1066 536645 358930 537211
rect 1066 535557 358930 536123
rect 1066 534469 358930 535035
rect 1066 533381 358930 533947
rect 1066 532293 358930 532859
rect 1066 531205 358930 531771
rect 1066 530117 358930 530683
rect 1066 529029 358930 529595
rect 1066 527941 358930 528507
rect 1066 526853 358930 527419
rect 1066 525765 358930 526331
rect 1066 524677 358930 525243
rect 1066 523589 358930 524155
rect 1066 522501 358930 523067
rect 1066 521413 358930 521979
rect 1066 520325 358930 520891
rect 1066 519237 358930 519803
rect 1066 518149 358930 518715
rect 1066 517061 358930 517627
rect 1066 515973 358930 516539
rect 1066 514885 358930 515451
rect 1066 513797 358930 514363
rect 1066 512709 358930 513275
rect 1066 511621 358930 512187
rect 1066 510533 358930 511099
rect 1066 509445 358930 510011
rect 1066 508357 358930 508923
rect 1066 507269 358930 507835
rect 1066 506181 358930 506747
rect 1066 505093 358930 505659
rect 1066 504005 358930 504571
rect 1066 502917 358930 503483
rect 1066 501829 358930 502395
rect 1066 500741 358930 501307
rect 1066 499653 358930 500219
rect 1066 498565 358930 499131
rect 1066 497477 358930 498043
rect 1066 496389 358930 496955
rect 1066 495301 358930 495867
rect 1066 494213 358930 494779
rect 1066 493125 358930 493691
rect 1066 492037 358930 492603
rect 1066 490949 358930 491515
rect 1066 489861 358930 490427
rect 1066 488773 358930 489339
rect 1066 487685 358930 488251
rect 1066 486597 358930 487163
rect 1066 485509 358930 486075
rect 1066 484421 358930 484987
rect 1066 483333 358930 483899
rect 1066 482245 358930 482811
rect 1066 481157 358930 481723
rect 1066 480069 358930 480635
rect 1066 478981 358930 479547
rect 1066 477893 358930 478459
rect 1066 476805 358930 477371
rect 1066 475717 358930 476283
rect 1066 474629 358930 475195
rect 1066 473541 358930 474107
rect 1066 472453 358930 473019
rect 1066 471365 358930 471931
rect 1066 470277 358930 470843
rect 1066 469189 358930 469755
rect 1066 468101 358930 468667
rect 1066 467013 358930 467579
rect 1066 465925 358930 466491
rect 1066 464837 358930 465403
rect 1066 463749 358930 464315
rect 1066 462661 358930 463227
rect 1066 461573 358930 462139
rect 1066 460485 358930 461051
rect 1066 459397 358930 459963
rect 1066 458309 358930 458875
rect 1066 457221 358930 457787
rect 1066 456133 358930 456699
rect 1066 455045 358930 455611
rect 1066 453957 358930 454523
rect 1066 452869 358930 453435
rect 1066 451781 358930 452347
rect 1066 450693 358930 451259
rect 1066 449605 358930 450171
rect 1066 448517 358930 449083
rect 1066 447429 358930 447995
rect 1066 446341 358930 446907
rect 1066 445253 358930 445819
rect 1066 444165 358930 444731
rect 1066 443077 358930 443643
rect 1066 441989 358930 442555
rect 1066 440901 358930 441467
rect 1066 439813 358930 440379
rect 1066 438725 358930 439291
rect 1066 437637 358930 438203
rect 1066 436549 358930 437115
rect 1066 435461 358930 436027
rect 1066 434373 358930 434939
rect 1066 433285 358930 433851
rect 1066 432197 358930 432763
rect 1066 431109 358930 431675
rect 1066 430021 358930 430587
rect 1066 428933 358930 429499
rect 1066 427845 358930 428411
rect 1066 426757 358930 427323
rect 1066 425669 358930 426235
rect 1066 424581 358930 425147
rect 1066 423493 358930 424059
rect 1066 422405 358930 422971
rect 1066 421317 358930 421883
rect 1066 420229 358930 420795
rect 1066 419141 358930 419707
rect 1066 418053 358930 418619
rect 1066 416965 358930 417531
rect 1066 415877 358930 416443
rect 1066 414789 358930 415355
rect 1066 413701 358930 414267
rect 1066 412613 358930 413179
rect 1066 411525 358930 412091
rect 1066 410437 358930 411003
rect 1066 409349 358930 409915
rect 1066 408261 358930 408827
rect 1066 407173 358930 407739
rect 1066 406085 358930 406651
rect 1066 404997 358930 405563
rect 1066 403909 358930 404475
rect 1066 402821 358930 403387
rect 1066 401733 358930 402299
rect 1066 400645 358930 401211
rect 1066 399557 358930 400123
rect 1066 398469 358930 399035
rect 1066 397381 358930 397947
rect 1066 396293 358930 396859
rect 1066 395205 358930 395771
rect 1066 394117 358930 394683
rect 1066 393029 358930 393595
rect 1066 391941 358930 392507
rect 1066 390853 358930 391419
rect 1066 389765 358930 390331
rect 1066 388677 358930 389243
rect 1066 387589 358930 388155
rect 1066 386501 358930 387067
rect 1066 385413 358930 385979
rect 1066 384325 358930 384891
rect 1066 383237 358930 383803
rect 1066 382149 358930 382715
rect 1066 381061 358930 381627
rect 1066 379973 358930 380539
rect 1066 378885 358930 379451
rect 1066 377797 358930 378363
rect 1066 376709 358930 377275
rect 1066 375621 358930 376187
rect 1066 374533 358930 375099
rect 1066 373445 358930 374011
rect 1066 372357 358930 372923
rect 1066 371269 358930 371835
rect 1066 370181 358930 370747
rect 1066 369093 358930 369659
rect 1066 368005 358930 368571
rect 1066 366917 358930 367483
rect 1066 365829 358930 366395
rect 1066 364741 358930 365307
rect 1066 363653 358930 364219
rect 1066 362565 358930 363131
rect 1066 361477 358930 362043
rect 1066 360389 358930 360955
rect 1066 359301 358930 359867
rect 1066 358213 358930 358779
rect 1066 357125 358930 357691
rect 1066 356037 358930 356603
rect 1066 354949 358930 355515
rect 1066 353861 358930 354427
rect 1066 352773 358930 353339
rect 1066 351685 358930 352251
rect 1066 350597 358930 351163
rect 1066 349509 358930 350075
rect 1066 348421 358930 348987
rect 1066 347333 358930 347899
rect 1066 346245 358930 346811
rect 1066 345157 358930 345723
rect 1066 344069 358930 344635
rect 1066 342981 358930 343547
rect 1066 341893 358930 342459
rect 1066 340805 358930 341371
rect 1066 339717 358930 340283
rect 1066 338629 358930 339195
rect 1066 337541 358930 338107
rect 1066 336453 358930 337019
rect 1066 335365 358930 335931
rect 1066 334277 358930 334843
rect 1066 333189 358930 333755
rect 1066 332101 358930 332667
rect 1066 331013 358930 331579
rect 1066 329925 358930 330491
rect 1066 328837 358930 329403
rect 1066 327749 358930 328315
rect 1066 326661 358930 327227
rect 1066 325573 358930 326139
rect 1066 324485 358930 325051
rect 1066 323397 358930 323963
rect 1066 322309 358930 322875
rect 1066 321221 358930 321787
rect 1066 320133 358930 320699
rect 1066 319045 358930 319611
rect 1066 317957 358930 318523
rect 1066 316869 358930 317435
rect 1066 315781 358930 316347
rect 1066 314693 358930 315259
rect 1066 313605 358930 314171
rect 1066 312517 358930 313083
rect 1066 311429 358930 311995
rect 1066 310341 358930 310907
rect 1066 309253 358930 309819
rect 1066 308165 358930 308731
rect 1066 307077 358930 307643
rect 1066 305989 358930 306555
rect 1066 304901 358930 305467
rect 1066 303813 358930 304379
rect 1066 302725 358930 303291
rect 1066 301637 358930 302203
rect 1066 300549 358930 301115
rect 1066 299461 358930 300027
rect 1066 298373 358930 298939
rect 1066 297285 358930 297851
rect 1066 296197 358930 296763
rect 1066 295109 358930 295675
rect 1066 294021 358930 294587
rect 1066 292933 358930 293499
rect 1066 291845 358930 292411
rect 1066 290757 358930 291323
rect 1066 289669 358930 290235
rect 1066 288581 358930 289147
rect 1066 287493 358930 288059
rect 1066 286405 358930 286971
rect 1066 285317 358930 285883
rect 1066 284229 358930 284795
rect 1066 283141 358930 283707
rect 1066 282053 358930 282619
rect 1066 280965 358930 281531
rect 1066 279877 358930 280443
rect 1066 278789 358930 279355
rect 1066 277701 358930 278267
rect 1066 276613 358930 277179
rect 1066 275525 358930 276091
rect 1066 274437 358930 275003
rect 1066 273349 358930 273915
rect 1066 272261 358930 272827
rect 1066 271173 358930 271739
rect 1066 270085 358930 270651
rect 1066 268997 358930 269563
rect 1066 267909 358930 268475
rect 1066 266821 358930 267387
rect 1066 265733 358930 266299
rect 1066 264645 358930 265211
rect 1066 263557 358930 264123
rect 1066 262469 358930 263035
rect 1066 261381 358930 261947
rect 1066 260293 358930 260859
rect 1066 259205 358930 259771
rect 1066 258117 358930 258683
rect 1066 257029 358930 257595
rect 1066 255941 358930 256507
rect 1066 254853 358930 255419
rect 1066 253765 358930 254331
rect 1066 252677 358930 253243
rect 1066 251589 358930 252155
rect 1066 250501 358930 251067
rect 1066 249413 358930 249979
rect 1066 248325 358930 248891
rect 1066 247237 358930 247803
rect 1066 246149 358930 246715
rect 1066 245061 358930 245627
rect 1066 243973 358930 244539
rect 1066 242885 358930 243451
rect 1066 241797 358930 242363
rect 1066 240709 358930 241275
rect 1066 239621 358930 240187
rect 1066 238533 358930 239099
rect 1066 237445 358930 238011
rect 1066 236357 358930 236923
rect 1066 235269 358930 235835
rect 1066 234181 358930 234747
rect 1066 233093 358930 233659
rect 1066 232005 358930 232571
rect 1066 230917 358930 231483
rect 1066 229829 358930 230395
rect 1066 228741 358930 229307
rect 1066 227653 358930 228219
rect 1066 226565 358930 227131
rect 1066 225477 358930 226043
rect 1066 224389 358930 224955
rect 1066 223301 358930 223867
rect 1066 222213 358930 222779
rect 1066 221125 358930 221691
rect 1066 220037 358930 220603
rect 1066 218949 358930 219515
rect 1066 217861 358930 218427
rect 1066 216773 358930 217339
rect 1066 215685 358930 216251
rect 1066 214597 358930 215163
rect 1066 213509 358930 214075
rect 1066 212421 358930 212987
rect 1066 211333 358930 211899
rect 1066 210245 358930 210811
rect 1066 209157 358930 209723
rect 1066 208069 358930 208635
rect 1066 206981 358930 207547
rect 1066 205893 358930 206459
rect 1066 204805 358930 205371
rect 1066 203717 358930 204283
rect 1066 202629 358930 203195
rect 1066 201541 358930 202107
rect 1066 200453 358930 201019
rect 1066 199365 358930 199931
rect 1066 198277 358930 198843
rect 1066 197189 358930 197755
rect 1066 196101 358930 196667
rect 1066 195013 358930 195579
rect 1066 193925 358930 194491
rect 1066 192837 358930 193403
rect 1066 191749 358930 192315
rect 1066 190661 358930 191227
rect 1066 189573 358930 190139
rect 1066 188485 358930 189051
rect 1066 187397 358930 187963
rect 1066 186309 358930 186875
rect 1066 185221 358930 185787
rect 1066 184133 358930 184699
rect 1066 183045 358930 183611
rect 1066 181957 358930 182523
rect 1066 180869 358930 181435
rect 1066 179781 358930 180347
rect 1066 178693 358930 179259
rect 1066 177605 358930 178171
rect 1066 176517 358930 177083
rect 1066 175429 358930 175995
rect 1066 174341 358930 174907
rect 1066 173253 358930 173819
rect 1066 172165 358930 172731
rect 1066 171077 358930 171643
rect 1066 169989 358930 170555
rect 1066 168901 358930 169467
rect 1066 167813 358930 168379
rect 1066 166725 358930 167291
rect 1066 165637 358930 166203
rect 1066 164549 358930 165115
rect 1066 163461 358930 164027
rect 1066 162373 358930 162939
rect 1066 161285 358930 161851
rect 1066 160197 358930 160763
rect 1066 159109 358930 159675
rect 1066 158021 358930 158587
rect 1066 156933 358930 157499
rect 1066 155845 358930 156411
rect 1066 154757 358930 155323
rect 1066 153669 358930 154235
rect 1066 152581 358930 153147
rect 1066 151493 358930 152059
rect 1066 150405 358930 150971
rect 1066 149317 358930 149883
rect 1066 148229 358930 148795
rect 1066 147141 358930 147707
rect 1066 146053 358930 146619
rect 1066 144965 358930 145531
rect 1066 143877 358930 144443
rect 1066 142789 358930 143355
rect 1066 141701 358930 142267
rect 1066 140613 358930 141179
rect 1066 139525 358930 140091
rect 1066 138437 358930 139003
rect 1066 137349 358930 137915
rect 1066 136261 358930 136827
rect 1066 135173 358930 135739
rect 1066 134085 358930 134651
rect 1066 132997 358930 133563
rect 1066 131909 358930 132475
rect 1066 130821 358930 131387
rect 1066 129733 358930 130299
rect 1066 128645 358930 129211
rect 1066 127557 358930 128123
rect 1066 126469 358930 127035
rect 1066 125381 358930 125947
rect 1066 124293 358930 124859
rect 1066 123205 358930 123771
rect 1066 122117 358930 122683
rect 1066 121029 358930 121595
rect 1066 119941 358930 120507
rect 1066 118853 358930 119419
rect 1066 117765 358930 118331
rect 1066 116677 358930 117243
rect 1066 115589 358930 116155
rect 1066 114501 358930 115067
rect 1066 113413 358930 113979
rect 1066 112325 358930 112891
rect 1066 111237 358930 111803
rect 1066 110149 358930 110715
rect 1066 109061 358930 109627
rect 1066 107973 358930 108539
rect 1066 106885 358930 107451
rect 1066 105797 358930 106363
rect 1066 104709 358930 105275
rect 1066 103621 358930 104187
rect 1066 102533 358930 103099
rect 1066 101445 358930 102011
rect 1066 100357 358930 100923
rect 1066 99269 358930 99835
rect 1066 98181 358930 98747
rect 1066 97093 358930 97659
rect 1066 96005 358930 96571
rect 1066 94917 358930 95483
rect 1066 93829 358930 94395
rect 1066 92741 358930 93307
rect 1066 91653 358930 92219
rect 1066 90565 358930 91131
rect 1066 89477 358930 90043
rect 1066 88389 358930 88955
rect 1066 87301 358930 87867
rect 1066 86213 358930 86779
rect 1066 85125 358930 85691
rect 1066 84037 358930 84603
rect 1066 82949 358930 83515
rect 1066 81861 358930 82427
rect 1066 80773 358930 81339
rect 1066 79685 358930 80251
rect 1066 78597 358930 79163
rect 1066 77509 358930 78075
rect 1066 76421 358930 76987
rect 1066 75333 358930 75899
rect 1066 74245 358930 74811
rect 1066 73157 358930 73723
rect 1066 72069 358930 72635
rect 1066 70981 358930 71547
rect 1066 69893 358930 70459
rect 1066 68805 358930 69371
rect 1066 67717 358930 68283
rect 1066 66629 358930 67195
rect 1066 65541 358930 66107
rect 1066 64453 358930 65019
rect 1066 63365 358930 63931
rect 1066 62277 358930 62843
rect 1066 61189 358930 61755
rect 1066 60101 358930 60667
rect 1066 59013 358930 59579
rect 1066 57925 358930 58491
rect 1066 56837 358930 57403
rect 1066 55749 358930 56315
rect 1066 54661 358930 55227
rect 1066 53573 358930 54139
rect 1066 52485 358930 53051
rect 1066 51397 358930 51963
rect 1066 50309 358930 50875
rect 1066 49221 358930 49787
rect 1066 48133 358930 48699
rect 1066 47045 358930 47611
rect 1066 45957 358930 46523
rect 1066 44869 358930 45435
rect 1066 43781 358930 44347
rect 1066 42693 358930 43259
rect 1066 41605 358930 42171
rect 1066 40517 358930 41083
rect 1066 39429 358930 39995
rect 1066 38341 358930 38907
rect 1066 37253 358930 37819
rect 1066 36165 358930 36731
rect 1066 35077 358930 35643
rect 1066 33989 358930 34555
rect 1066 32901 358930 33467
rect 1066 31813 358930 32379
rect 1066 30725 358930 31291
rect 1066 29637 358930 30203
rect 1066 28549 358930 29115
rect 1066 27461 358930 28027
rect 1066 26373 358930 26939
rect 1066 25285 358930 25851
rect 1066 24197 358930 24763
rect 1066 23109 358930 23675
rect 1066 22021 358930 22587
rect 1066 20933 358930 21499
rect 1066 19845 358930 20411
rect 1066 18757 358930 19323
rect 1066 17669 358930 18235
rect 1066 16581 358930 17147
rect 1066 15493 358930 16059
rect 1066 14405 358930 14971
rect 1066 13317 358930 13883
rect 1066 12229 358930 12795
rect 1066 11141 358930 11707
rect 1066 10053 358930 10619
rect 1066 8965 358930 9531
rect 1066 7877 358930 8443
rect 1066 6789 358930 7355
rect 1066 5701 358930 6267
rect 1066 4613 358930 5179
rect 1066 3525 358930 4091
rect 1066 2437 358930 3003
<< obsli1 >>
rect 1104 2159 358892 617457
<< obsm1 >>
rect 1104 2128 359430 617488
<< obsm2 >>
rect 4214 2139 359424 617477
<< metal3 >>
rect 359200 612280 360000 612400
rect 359200 601672 360000 601792
rect 359200 591064 360000 591184
rect 359200 580456 360000 580576
rect 359200 569848 360000 569968
rect 359200 559240 360000 559360
rect 359200 548632 360000 548752
rect 359200 538024 360000 538144
rect 359200 527416 360000 527536
rect 359200 516808 360000 516928
rect 359200 506200 360000 506320
rect 359200 495592 360000 495712
rect 359200 484984 360000 485104
rect 359200 474376 360000 474496
rect 359200 463768 360000 463888
rect 359200 453160 360000 453280
rect 359200 442552 360000 442672
rect 359200 431944 360000 432064
rect 359200 421336 360000 421456
rect 359200 410728 360000 410848
rect 359200 400120 360000 400240
rect 359200 389512 360000 389632
rect 359200 378904 360000 379024
rect 359200 368296 360000 368416
rect 359200 357688 360000 357808
rect 359200 347080 360000 347200
rect 359200 336472 360000 336592
rect 359200 325864 360000 325984
rect 359200 315256 360000 315376
rect 359200 304648 360000 304768
rect 359200 294040 360000 294160
rect 359200 283432 360000 283552
rect 359200 272824 360000 272944
rect 359200 262216 360000 262336
rect 359200 251608 360000 251728
rect 359200 241000 360000 241120
rect 359200 230392 360000 230512
rect 359200 219784 360000 219904
rect 359200 209176 360000 209296
rect 359200 198568 360000 198688
rect 359200 187960 360000 188080
rect 359200 177352 360000 177472
rect 359200 166744 360000 166864
rect 359200 156136 360000 156256
rect 359200 145528 360000 145648
rect 359200 134920 360000 135040
rect 359200 124312 360000 124432
rect 359200 113704 360000 113824
rect 359200 103096 360000 103216
rect 359200 92488 360000 92608
rect 359200 81880 360000 82000
rect 359200 71272 360000 71392
rect 359200 60664 360000 60784
rect 359200 50056 360000 50176
rect 359200 39448 360000 39568
rect 359200 28840 360000 28960
rect 359200 18232 360000 18352
rect 359200 7624 360000 7744
<< obsm3 >>
rect 4210 612480 359247 617473
rect 4210 612200 359120 612480
rect 4210 601872 359247 612200
rect 4210 601592 359120 601872
rect 4210 591264 359247 601592
rect 4210 590984 359120 591264
rect 4210 580656 359247 590984
rect 4210 580376 359120 580656
rect 4210 570048 359247 580376
rect 4210 569768 359120 570048
rect 4210 559440 359247 569768
rect 4210 559160 359120 559440
rect 4210 548832 359247 559160
rect 4210 548552 359120 548832
rect 4210 538224 359247 548552
rect 4210 537944 359120 538224
rect 4210 527616 359247 537944
rect 4210 527336 359120 527616
rect 4210 517008 359247 527336
rect 4210 516728 359120 517008
rect 4210 506400 359247 516728
rect 4210 506120 359120 506400
rect 4210 495792 359247 506120
rect 4210 495512 359120 495792
rect 4210 485184 359247 495512
rect 4210 484904 359120 485184
rect 4210 474576 359247 484904
rect 4210 474296 359120 474576
rect 4210 463968 359247 474296
rect 4210 463688 359120 463968
rect 4210 453360 359247 463688
rect 4210 453080 359120 453360
rect 4210 442752 359247 453080
rect 4210 442472 359120 442752
rect 4210 432144 359247 442472
rect 4210 431864 359120 432144
rect 4210 421536 359247 431864
rect 4210 421256 359120 421536
rect 4210 410928 359247 421256
rect 4210 410648 359120 410928
rect 4210 400320 359247 410648
rect 4210 400040 359120 400320
rect 4210 389712 359247 400040
rect 4210 389432 359120 389712
rect 4210 379104 359247 389432
rect 4210 378824 359120 379104
rect 4210 368496 359247 378824
rect 4210 368216 359120 368496
rect 4210 357888 359247 368216
rect 4210 357608 359120 357888
rect 4210 347280 359247 357608
rect 4210 347000 359120 347280
rect 4210 336672 359247 347000
rect 4210 336392 359120 336672
rect 4210 326064 359247 336392
rect 4210 325784 359120 326064
rect 4210 315456 359247 325784
rect 4210 315176 359120 315456
rect 4210 304848 359247 315176
rect 4210 304568 359120 304848
rect 4210 294240 359247 304568
rect 4210 293960 359120 294240
rect 4210 283632 359247 293960
rect 4210 283352 359120 283632
rect 4210 273024 359247 283352
rect 4210 272744 359120 273024
rect 4210 262416 359247 272744
rect 4210 262136 359120 262416
rect 4210 251808 359247 262136
rect 4210 251528 359120 251808
rect 4210 241200 359247 251528
rect 4210 240920 359120 241200
rect 4210 230592 359247 240920
rect 4210 230312 359120 230592
rect 4210 219984 359247 230312
rect 4210 219704 359120 219984
rect 4210 209376 359247 219704
rect 4210 209096 359120 209376
rect 4210 198768 359247 209096
rect 4210 198488 359120 198768
rect 4210 188160 359247 198488
rect 4210 187880 359120 188160
rect 4210 177552 359247 187880
rect 4210 177272 359120 177552
rect 4210 166944 359247 177272
rect 4210 166664 359120 166944
rect 4210 156336 359247 166664
rect 4210 156056 359120 156336
rect 4210 145728 359247 156056
rect 4210 145448 359120 145728
rect 4210 135120 359247 145448
rect 4210 134840 359120 135120
rect 4210 124512 359247 134840
rect 4210 124232 359120 124512
rect 4210 113904 359247 124232
rect 4210 113624 359120 113904
rect 4210 103296 359247 113624
rect 4210 103016 359120 103296
rect 4210 92688 359247 103016
rect 4210 92408 359120 92688
rect 4210 82080 359247 92408
rect 4210 81800 359120 82080
rect 4210 71472 359247 81800
rect 4210 71192 359120 71472
rect 4210 60864 359247 71192
rect 4210 60584 359120 60864
rect 4210 50256 359247 60584
rect 4210 49976 359120 50256
rect 4210 39648 359247 49976
rect 4210 39368 359120 39648
rect 4210 29040 359247 39368
rect 4210 28760 359120 29040
rect 4210 18432 359247 28760
rect 4210 18152 359120 18432
rect 4210 7824 359247 18152
rect 4210 7544 359120 7824
rect 4210 2143 359247 7544
<< metal4 >>
rect 4208 2128 4528 617488
rect 19568 2128 19888 617488
rect 34928 2128 35248 617488
rect 50288 2128 50608 617488
rect 65648 2128 65968 617488
rect 81008 2128 81328 617488
rect 96368 2128 96688 617488
rect 111728 2128 112048 617488
rect 127088 2128 127408 617488
rect 142448 2128 142768 617488
rect 157808 2128 158128 617488
rect 173168 2128 173488 617488
rect 188528 2128 188848 617488
rect 203888 2128 204208 617488
rect 219248 2128 219568 617488
rect 234608 2128 234928 617488
rect 249968 2128 250288 617488
rect 265328 2128 265648 617488
rect 280688 2128 281008 617488
rect 296048 2128 296368 617488
rect 311408 2128 311728 617488
rect 326768 2128 327088 617488
rect 342128 2128 342448 617488
rect 357488 2128 357808 617488
<< obsm4 >>
rect 50843 10915 65568 614957
rect 66048 10915 80928 614957
rect 81408 10915 96288 614957
rect 96768 10915 111648 614957
rect 112128 10915 127008 614957
rect 127488 10915 142368 614957
rect 142848 10915 157728 614957
rect 158208 10915 173088 614957
rect 173568 10915 188448 614957
rect 188928 10915 203808 614957
rect 204288 10915 219168 614957
rect 219648 10915 234528 614957
rect 235008 10915 249888 614957
rect 250368 10915 265248 614957
rect 265728 10915 280608 614957
rect 281088 10915 295968 614957
rect 296448 10915 311328 614957
rect 311808 10915 326688 614957
rect 327168 10915 342048 614957
rect 342528 10915 353037 614957
<< labels >>
rlabel metal3 s 359200 294040 360000 294160 6 clk
port 1 nsew signal input
rlabel metal3 s 359200 7624 360000 7744 6 io_in[0]
port 2 nsew signal input
rlabel metal3 s 359200 113704 360000 113824 6 io_in[10]
port 3 nsew signal input
rlabel metal3 s 359200 124312 360000 124432 6 io_in[11]
port 4 nsew signal input
rlabel metal3 s 359200 134920 360000 135040 6 io_in[12]
port 5 nsew signal input
rlabel metal3 s 359200 145528 360000 145648 6 io_in[13]
port 6 nsew signal input
rlabel metal3 s 359200 156136 360000 156256 6 io_in[14]
port 7 nsew signal input
rlabel metal3 s 359200 166744 360000 166864 6 io_in[15]
port 8 nsew signal input
rlabel metal3 s 359200 177352 360000 177472 6 io_in[16]
port 9 nsew signal input
rlabel metal3 s 359200 187960 360000 188080 6 io_in[17]
port 10 nsew signal input
rlabel metal3 s 359200 198568 360000 198688 6 io_in[18]
port 11 nsew signal input
rlabel metal3 s 359200 209176 360000 209296 6 io_in[19]
port 12 nsew signal input
rlabel metal3 s 359200 18232 360000 18352 6 io_in[1]
port 13 nsew signal input
rlabel metal3 s 359200 219784 360000 219904 6 io_in[20]
port 14 nsew signal input
rlabel metal3 s 359200 230392 360000 230512 6 io_in[21]
port 15 nsew signal input
rlabel metal3 s 359200 241000 360000 241120 6 io_in[22]
port 16 nsew signal input
rlabel metal3 s 359200 251608 360000 251728 6 io_in[23]
port 17 nsew signal input
rlabel metal3 s 359200 262216 360000 262336 6 io_in[24]
port 18 nsew signal input
rlabel metal3 s 359200 272824 360000 272944 6 io_in[25]
port 19 nsew signal input
rlabel metal3 s 359200 283432 360000 283552 6 io_in[26]
port 20 nsew signal input
rlabel metal3 s 359200 28840 360000 28960 6 io_in[2]
port 21 nsew signal input
rlabel metal3 s 359200 39448 360000 39568 6 io_in[3]
port 22 nsew signal input
rlabel metal3 s 359200 50056 360000 50176 6 io_in[4]
port 23 nsew signal input
rlabel metal3 s 359200 60664 360000 60784 6 io_in[5]
port 24 nsew signal input
rlabel metal3 s 359200 71272 360000 71392 6 io_in[6]
port 25 nsew signal input
rlabel metal3 s 359200 81880 360000 82000 6 io_in[7]
port 26 nsew signal input
rlabel metal3 s 359200 92488 360000 92608 6 io_in[8]
port 27 nsew signal input
rlabel metal3 s 359200 103096 360000 103216 6 io_in[9]
port 28 nsew signal input
rlabel metal3 s 359200 612280 360000 612400 6 io_oeb
port 29 nsew signal output
rlabel metal3 s 359200 315256 360000 315376 6 io_out[0]
port 30 nsew signal output
rlabel metal3 s 359200 421336 360000 421456 6 io_out[10]
port 31 nsew signal output
rlabel metal3 s 359200 431944 360000 432064 6 io_out[11]
port 32 nsew signal output
rlabel metal3 s 359200 442552 360000 442672 6 io_out[12]
port 33 nsew signal output
rlabel metal3 s 359200 453160 360000 453280 6 io_out[13]
port 34 nsew signal output
rlabel metal3 s 359200 463768 360000 463888 6 io_out[14]
port 35 nsew signal output
rlabel metal3 s 359200 474376 360000 474496 6 io_out[15]
port 36 nsew signal output
rlabel metal3 s 359200 484984 360000 485104 6 io_out[16]
port 37 nsew signal output
rlabel metal3 s 359200 495592 360000 495712 6 io_out[17]
port 38 nsew signal output
rlabel metal3 s 359200 506200 360000 506320 6 io_out[18]
port 39 nsew signal output
rlabel metal3 s 359200 516808 360000 516928 6 io_out[19]
port 40 nsew signal output
rlabel metal3 s 359200 325864 360000 325984 6 io_out[1]
port 41 nsew signal output
rlabel metal3 s 359200 527416 360000 527536 6 io_out[20]
port 42 nsew signal output
rlabel metal3 s 359200 538024 360000 538144 6 io_out[21]
port 43 nsew signal output
rlabel metal3 s 359200 548632 360000 548752 6 io_out[22]
port 44 nsew signal output
rlabel metal3 s 359200 559240 360000 559360 6 io_out[23]
port 45 nsew signal output
rlabel metal3 s 359200 569848 360000 569968 6 io_out[24]
port 46 nsew signal output
rlabel metal3 s 359200 580456 360000 580576 6 io_out[25]
port 47 nsew signal output
rlabel metal3 s 359200 591064 360000 591184 6 io_out[26]
port 48 nsew signal output
rlabel metal3 s 359200 601672 360000 601792 6 io_out[27]
port 49 nsew signal output
rlabel metal3 s 359200 336472 360000 336592 6 io_out[2]
port 50 nsew signal output
rlabel metal3 s 359200 347080 360000 347200 6 io_out[3]
port 51 nsew signal output
rlabel metal3 s 359200 357688 360000 357808 6 io_out[4]
port 52 nsew signal output
rlabel metal3 s 359200 368296 360000 368416 6 io_out[5]
port 53 nsew signal output
rlabel metal3 s 359200 378904 360000 379024 6 io_out[6]
port 54 nsew signal output
rlabel metal3 s 359200 389512 360000 389632 6 io_out[7]
port 55 nsew signal output
rlabel metal3 s 359200 400120 360000 400240 6 io_out[8]
port 56 nsew signal output
rlabel metal3 s 359200 410728 360000 410848 6 io_out[9]
port 57 nsew signal output
rlabel metal3 s 359200 304648 360000 304768 6 rst
port 58 nsew signal input
rlabel metal4 s 4208 2128 4528 617488 6 vccd1
port 59 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 617488 6 vccd1
port 59 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 617488 6 vccd1
port 59 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 617488 6 vccd1
port 59 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 617488 6 vccd1
port 59 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 617488 6 vccd1
port 59 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 617488 6 vccd1
port 59 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 617488 6 vccd1
port 59 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 617488 6 vccd1
port 59 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 617488 6 vccd1
port 59 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 617488 6 vccd1
port 59 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 617488 6 vccd1
port 59 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 617488 6 vssd1
port 60 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 617488 6 vssd1
port 60 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 617488 6 vssd1
port 60 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 617488 6 vssd1
port 60 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 617488 6 vssd1
port 60 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 617488 6 vssd1
port 60 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 617488 6 vssd1
port 60 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 617488 6 vssd1
port 60 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 617488 6 vssd1
port 60 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 617488 6 vssd1
port 60 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 617488 6 vssd1
port 60 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 617488 6 vssd1
port 60 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 360000 620000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 261593458
string GDS_FILE /run/media/tholin/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/AS512512512/runs/23_03_27_08_03/results/signoff/wrapped_as512512512.magic.gds
string GDS_START 1763644
<< end >>

