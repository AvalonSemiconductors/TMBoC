magic
tech sky130B
magscale 1 2
timestamp 1682095682
<< nwell >>
rect 1066 22021 23866 22342
rect 1066 20933 23866 21499
rect 1066 19845 23866 20411
rect 1066 18757 23866 19323
rect 1066 17669 23866 18235
rect 1066 16581 23866 17147
rect 1066 15493 23866 16059
rect 1066 14405 23866 14971
rect 1066 13317 23866 13883
rect 1066 12229 23866 12795
rect 1066 11141 23866 11707
rect 1066 10053 23866 10619
rect 1066 8965 23866 9531
rect 1066 7877 23866 8443
rect 1066 6789 23866 7355
rect 1066 5701 23866 6267
rect 1066 4613 23866 5179
rect 1066 3525 23866 4091
rect 1066 2437 23866 3003
<< obsli1 >>
rect 1104 2159 23828 22321
<< obsm1 >>
rect 1104 1164 23987 22352
<< metal2 >>
rect 2502 24200 2558 25000
rect 7470 24200 7526 25000
rect 12438 24200 12494 25000
rect 17406 24200 17462 25000
rect 22374 24200 22430 25000
rect 1490 0 1546 800
rect 2134 0 2190 800
rect 2778 0 2834 800
rect 3422 0 3478 800
rect 4066 0 4122 800
rect 4710 0 4766 800
rect 5354 0 5410 800
rect 5998 0 6054 800
rect 6642 0 6698 800
rect 7286 0 7342 800
rect 7930 0 7986 800
rect 8574 0 8630 800
rect 9218 0 9274 800
rect 9862 0 9918 800
rect 10506 0 10562 800
rect 11150 0 11206 800
rect 11794 0 11850 800
rect 12438 0 12494 800
rect 13082 0 13138 800
rect 13726 0 13782 800
rect 14370 0 14426 800
rect 15014 0 15070 800
rect 15658 0 15714 800
rect 16302 0 16358 800
rect 16946 0 17002 800
rect 17590 0 17646 800
rect 18234 0 18290 800
rect 18878 0 18934 800
rect 19522 0 19578 800
rect 20166 0 20222 800
rect 20810 0 20866 800
rect 21454 0 21510 800
rect 22098 0 22154 800
rect 22742 0 22798 800
rect 23386 0 23442 800
<< obsm2 >>
rect 1492 24144 2446 24200
rect 2614 24144 7414 24200
rect 7582 24144 12382 24200
rect 12550 24144 17350 24200
rect 17518 24144 22318 24200
rect 22486 24144 23981 24200
rect 1492 856 23981 24144
rect 1602 734 2078 856
rect 2246 734 2722 856
rect 2890 734 3366 856
rect 3534 734 4010 856
rect 4178 734 4654 856
rect 4822 734 5298 856
rect 5466 734 5942 856
rect 6110 734 6586 856
rect 6754 734 7230 856
rect 7398 734 7874 856
rect 8042 734 8518 856
rect 8686 734 9162 856
rect 9330 734 9806 856
rect 9974 734 10450 856
rect 10618 734 11094 856
rect 11262 734 11738 856
rect 11906 734 12382 856
rect 12550 734 13026 856
rect 13194 734 13670 856
rect 13838 734 14314 856
rect 14482 734 14958 856
rect 15126 734 15602 856
rect 15770 734 16246 856
rect 16414 734 16890 856
rect 17058 734 17534 856
rect 17702 734 18178 856
rect 18346 734 18822 856
rect 18990 734 19466 856
rect 19634 734 20110 856
rect 20278 734 20754 856
rect 20922 734 21398 856
rect 21566 734 22042 856
rect 22210 734 22686 856
rect 22854 734 23330 856
rect 23498 734 23981 856
<< obsm3 >>
rect 2313 2143 23985 22337
<< metal4 >>
rect 3784 2128 4104 22352
rect 6624 2128 6944 22352
rect 9465 2128 9785 22352
rect 12305 2128 12625 22352
rect 15146 2128 15466 22352
rect 17986 2128 18306 22352
rect 20827 2128 21147 22352
rect 23667 2128 23987 22352
<< obsm4 >>
rect 5395 4659 6544 20773
rect 7024 4659 9385 20773
rect 9865 4659 12225 20773
rect 12705 4659 15066 20773
rect 15546 4659 17906 20773
rect 18386 4659 20747 20773
rect 21227 4659 22389 20773
<< labels >>
rlabel metal2 s 2502 24200 2558 25000 6 clk
port 1 nsew signal input
rlabel metal2 s 12438 24200 12494 25000 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 17406 24200 17462 25000 6 io_in[1]
port 3 nsew signal input
rlabel metal2 s 22374 24200 22430 25000 6 io_in[2]
port 4 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 io_oeb[0]
port 5 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 io_oeb[10]
port 6 nsew signal output
rlabel metal2 s 13726 0 13782 800 6 io_oeb[11]
port 7 nsew signal output
rlabel metal2 s 14370 0 14426 800 6 io_oeb[12]
port 8 nsew signal output
rlabel metal2 s 15014 0 15070 800 6 io_oeb[13]
port 9 nsew signal output
rlabel metal2 s 15658 0 15714 800 6 io_oeb[14]
port 10 nsew signal output
rlabel metal2 s 16302 0 16358 800 6 io_oeb[15]
port 11 nsew signal output
rlabel metal2 s 16946 0 17002 800 6 io_oeb[16]
port 12 nsew signal output
rlabel metal2 s 17590 0 17646 800 6 io_oeb[17]
port 13 nsew signal output
rlabel metal2 s 18234 0 18290 800 6 io_oeb[18]
port 14 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 io_oeb[19]
port 15 nsew signal output
rlabel metal2 s 7286 0 7342 800 6 io_oeb[1]
port 16 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 io_oeb[20]
port 17 nsew signal output
rlabel metal2 s 20166 0 20222 800 6 io_oeb[21]
port 18 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 io_oeb[22]
port 19 nsew signal output
rlabel metal2 s 21454 0 21510 800 6 io_oeb[23]
port 20 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 io_oeb[24]
port 21 nsew signal output
rlabel metal2 s 22742 0 22798 800 6 io_oeb[25]
port 22 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 io_oeb[26]
port 23 nsew signal output
rlabel metal2 s 7930 0 7986 800 6 io_oeb[2]
port 24 nsew signal output
rlabel metal2 s 8574 0 8630 800 6 io_oeb[3]
port 25 nsew signal output
rlabel metal2 s 9218 0 9274 800 6 io_oeb[4]
port 26 nsew signal output
rlabel metal2 s 9862 0 9918 800 6 io_oeb[5]
port 27 nsew signal output
rlabel metal2 s 10506 0 10562 800 6 io_oeb[6]
port 28 nsew signal output
rlabel metal2 s 11150 0 11206 800 6 io_oeb[7]
port 29 nsew signal output
rlabel metal2 s 11794 0 11850 800 6 io_oeb[8]
port 30 nsew signal output
rlabel metal2 s 12438 0 12494 800 6 io_oeb[9]
port 31 nsew signal output
rlabel metal2 s 1490 0 1546 800 6 io_out[0]
port 32 nsew signal output
rlabel metal2 s 2134 0 2190 800 6 io_out[1]
port 33 nsew signal output
rlabel metal2 s 2778 0 2834 800 6 io_out[2]
port 34 nsew signal output
rlabel metal2 s 3422 0 3478 800 6 io_out[3]
port 35 nsew signal output
rlabel metal2 s 4066 0 4122 800 6 io_out[4]
port 36 nsew signal output
rlabel metal2 s 4710 0 4766 800 6 io_out[5]
port 37 nsew signal output
rlabel metal2 s 5354 0 5410 800 6 io_out[6]
port 38 nsew signal output
rlabel metal2 s 5998 0 6054 800 6 io_out[7]
port 39 nsew signal output
rlabel metal2 s 7470 24200 7526 25000 6 rst
port 40 nsew signal input
rlabel metal4 s 3784 2128 4104 22352 6 vccd1
port 41 nsew power bidirectional
rlabel metal4 s 9465 2128 9785 22352 6 vccd1
port 41 nsew power bidirectional
rlabel metal4 s 15146 2128 15466 22352 6 vccd1
port 41 nsew power bidirectional
rlabel metal4 s 20827 2128 21147 22352 6 vccd1
port 41 nsew power bidirectional
rlabel metal4 s 6624 2128 6944 22352 6 vssd1
port 42 nsew ground bidirectional
rlabel metal4 s 12305 2128 12625 22352 6 vssd1
port 42 nsew ground bidirectional
rlabel metal4 s 17986 2128 18306 22352 6 vssd1
port 42 nsew ground bidirectional
rlabel metal4 s 23667 2128 23987 22352 6 vssd1
port 42 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 25000 25000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2588334
string GDS_FILE /run/media/tholin/Data/Projects/MPW/TMBoC/openlane/LCD/runs/23_04_21_18_46/results/signoff/tt2_tholin_namebadge.magic.gds
string GDS_START 906428
<< end >>

