VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_as2650
  CLASS BLOCK ;
  FOREIGN wrapped_as2650 ;
  ORIGIN 0.000 0.000 ;
  SIZE 350.000 BY 350.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END clk
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 4.000 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 0.000 143.430 4.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 0.000 206.910 4.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 4.000 ;
    END
  END io_in[8]
  PIN io_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 339.360 4.000 339.960 ;
    END
  END io_oeb
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.280 4.000 131.880 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.520 4.000 144.120 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.760 4.000 156.360 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 4.000 168.600 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.480 4.000 193.080 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.720 4.000 205.320 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.960 4.000 217.560 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.200 4.000 229.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.680 4.000 254.280 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.920 4.000 266.520 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.160 4.000 278.760 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 290.400 4.000 291.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.880 4.000 315.480 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.120 4.000 327.720 ;
    END
  END io_out[26]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 4.000 82.920 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.560 4.000 95.160 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END io_out[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 0.000 333.870 4.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 337.520 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 337.520 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 344.080 337.365 ;
      LAYER met1 ;
        RECT 1.910 9.220 344.080 337.520 ;
      LAYER met2 ;
        RECT 1.470 4.280 340.300 339.845 ;
        RECT 1.470 4.000 15.910 4.280 ;
        RECT 16.750 4.000 47.650 4.280 ;
        RECT 48.490 4.000 79.390 4.280 ;
        RECT 80.230 4.000 111.130 4.280 ;
        RECT 111.970 4.000 142.870 4.280 ;
        RECT 143.710 4.000 174.610 4.280 ;
        RECT 175.450 4.000 206.350 4.280 ;
        RECT 207.190 4.000 238.090 4.280 ;
        RECT 238.930 4.000 269.830 4.280 ;
        RECT 270.670 4.000 301.570 4.280 ;
        RECT 302.410 4.000 333.310 4.280 ;
        RECT 334.150 4.000 340.300 4.280 ;
      LAYER met3 ;
        RECT 4.400 338.960 329.830 339.825 ;
        RECT 1.445 328.120 329.830 338.960 ;
        RECT 4.400 326.720 329.830 328.120 ;
        RECT 1.445 315.880 329.830 326.720 ;
        RECT 4.400 314.480 329.830 315.880 ;
        RECT 1.445 303.640 329.830 314.480 ;
        RECT 4.400 302.240 329.830 303.640 ;
        RECT 1.445 291.400 329.830 302.240 ;
        RECT 4.400 290.000 329.830 291.400 ;
        RECT 1.445 279.160 329.830 290.000 ;
        RECT 4.400 277.760 329.830 279.160 ;
        RECT 1.445 266.920 329.830 277.760 ;
        RECT 4.400 265.520 329.830 266.920 ;
        RECT 1.445 254.680 329.830 265.520 ;
        RECT 4.400 253.280 329.830 254.680 ;
        RECT 1.445 242.440 329.830 253.280 ;
        RECT 4.400 241.040 329.830 242.440 ;
        RECT 1.445 230.200 329.830 241.040 ;
        RECT 4.400 228.800 329.830 230.200 ;
        RECT 1.445 217.960 329.830 228.800 ;
        RECT 4.400 216.560 329.830 217.960 ;
        RECT 1.445 205.720 329.830 216.560 ;
        RECT 4.400 204.320 329.830 205.720 ;
        RECT 1.445 193.480 329.830 204.320 ;
        RECT 4.400 192.080 329.830 193.480 ;
        RECT 1.445 181.240 329.830 192.080 ;
        RECT 4.400 179.840 329.830 181.240 ;
        RECT 1.445 169.000 329.830 179.840 ;
        RECT 4.400 167.600 329.830 169.000 ;
        RECT 1.445 156.760 329.830 167.600 ;
        RECT 4.400 155.360 329.830 156.760 ;
        RECT 1.445 144.520 329.830 155.360 ;
        RECT 4.400 143.120 329.830 144.520 ;
        RECT 1.445 132.280 329.830 143.120 ;
        RECT 4.400 130.880 329.830 132.280 ;
        RECT 1.445 120.040 329.830 130.880 ;
        RECT 4.400 118.640 329.830 120.040 ;
        RECT 1.445 107.800 329.830 118.640 ;
        RECT 4.400 106.400 329.830 107.800 ;
        RECT 1.445 95.560 329.830 106.400 ;
        RECT 4.400 94.160 329.830 95.560 ;
        RECT 1.445 83.320 329.830 94.160 ;
        RECT 4.400 81.920 329.830 83.320 ;
        RECT 1.445 71.080 329.830 81.920 ;
        RECT 4.400 69.680 329.830 71.080 ;
        RECT 1.445 58.840 329.830 69.680 ;
        RECT 4.400 57.440 329.830 58.840 ;
        RECT 1.445 46.600 329.830 57.440 ;
        RECT 4.400 45.200 329.830 46.600 ;
        RECT 1.445 34.360 329.830 45.200 ;
        RECT 4.400 32.960 329.830 34.360 ;
        RECT 1.445 22.120 329.830 32.960 ;
        RECT 4.400 20.720 329.830 22.120 ;
        RECT 1.445 9.880 329.830 20.720 ;
        RECT 4.400 9.015 329.830 9.880 ;
      LAYER met4 ;
        RECT 3.975 11.735 20.640 333.705 ;
        RECT 23.040 11.735 97.440 333.705 ;
        RECT 99.840 11.735 174.240 333.705 ;
        RECT 176.640 11.735 251.040 333.705 ;
        RECT 253.440 11.735 281.225 333.705 ;
  END
END wrapped_as2650
END LIBRARY

