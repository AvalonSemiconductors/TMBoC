magic
tech sky130B
magscale 1 2
timestamp 1687097953
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 429838 700748 429844 700800
rect 429896 700788 429902 700800
rect 445110 700788 445116 700800
rect 429896 700760 445116 700788
rect 429896 700748 429902 700760
rect 445110 700748 445116 700760
rect 445168 700748 445174 700800
rect 364978 700680 364984 700732
rect 365036 700720 365042 700732
rect 445018 700720 445024 700732
rect 365036 700692 445024 700720
rect 365036 700680 365042 700692
rect 445018 700680 445024 700692
rect 445076 700680 445082 700732
rect 332502 700612 332508 700664
rect 332560 700652 332566 700664
rect 446490 700652 446496 700664
rect 332560 700624 446496 700652
rect 332560 700612 332566 700624
rect 446490 700612 446496 700624
rect 446548 700612 446554 700664
rect 300118 700544 300124 700596
rect 300176 700584 300182 700596
rect 449158 700584 449164 700596
rect 300176 700556 449164 700584
rect 300176 700544 300182 700556
rect 449158 700544 449164 700556
rect 449216 700544 449222 700596
rect 283834 700476 283840 700528
rect 283892 700516 283898 700528
rect 446398 700516 446404 700528
rect 283892 700488 446404 700516
rect 283892 700476 283898 700488
rect 446398 700476 446404 700488
rect 446456 700476 446462 700528
rect 154114 700408 154120 700460
rect 154172 700448 154178 700460
rect 416038 700448 416044 700460
rect 154172 700420 416044 700448
rect 154172 700408 154178 700420
rect 416038 700408 416044 700420
rect 416096 700408 416102 700460
rect 444282 700408 444288 700460
rect 444340 700448 444346 700460
rect 494790 700448 494796 700460
rect 444340 700420 494796 700448
rect 444340 700408 444346 700420
rect 494790 700408 494796 700420
rect 494848 700408 494854 700460
rect 105446 700340 105452 700392
rect 105504 700380 105510 700392
rect 445202 700380 445208 700392
rect 105504 700352 445208 700380
rect 105504 700340 105510 700352
rect 445202 700340 445208 700352
rect 445260 700340 445266 700392
rect 445662 700340 445668 700392
rect 445720 700380 445726 700392
rect 478506 700380 478512 700392
rect 445720 700352 478512 700380
rect 445720 700340 445726 700352
rect 478506 700340 478512 700352
rect 478564 700340 478570 700392
rect 40494 700272 40500 700324
rect 40552 700312 40558 700324
rect 449250 700312 449256 700324
rect 40552 700284 449256 700312
rect 40552 700272 40558 700284
rect 449250 700272 449256 700284
rect 449308 700272 449314 700324
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 347774 685312 347780 685364
rect 347832 685352 347838 685364
rect 446674 685352 446680 685364
rect 347832 685324 446680 685352
rect 347832 685312 347838 685324
rect 446674 685312 446680 685324
rect 446732 685312 446738 685364
rect 218054 685244 218060 685296
rect 218112 685284 218118 685296
rect 446582 685284 446588 685296
rect 218112 685256 446588 685284
rect 218112 685244 218118 685256
rect 446582 685244 446588 685256
rect 446640 685244 446646 685296
rect 88334 685176 88340 685228
rect 88392 685216 88398 685228
rect 416222 685216 416228 685228
rect 88392 685188 416228 685216
rect 88392 685176 88398 685188
rect 416222 685176 416228 685188
rect 416280 685176 416286 685228
rect 71774 685108 71780 685160
rect 71832 685148 71838 685160
rect 419350 685148 419356 685160
rect 71832 685120 419356 685148
rect 71832 685108 71838 685120
rect 419350 685108 419356 685120
rect 419408 685108 419414 685160
rect 19978 684768 19984 684820
rect 20036 684808 20042 684820
rect 419442 684808 419448 684820
rect 20036 684780 419448 684808
rect 20036 684768 20042 684780
rect 419442 684768 419448 684780
rect 419500 684768 419506 684820
rect 3970 684700 3976 684752
rect 4028 684740 4034 684752
rect 418798 684740 418804 684752
rect 4028 684712 418804 684740
rect 4028 684700 4034 684712
rect 418798 684700 418804 684712
rect 418856 684700 418862 684752
rect 3602 684632 3608 684684
rect 3660 684672 3666 684684
rect 418982 684672 418988 684684
rect 3660 684644 418988 684672
rect 3660 684632 3666 684644
rect 418982 684632 418988 684644
rect 419040 684632 419046 684684
rect 3418 684564 3424 684616
rect 3476 684604 3482 684616
rect 419074 684604 419080 684616
rect 3476 684576 419080 684604
rect 3476 684564 3482 684576
rect 419074 684564 419080 684576
rect 419132 684564 419138 684616
rect 3326 684496 3332 684548
rect 3384 684536 3390 684548
rect 418890 684536 418896 684548
rect 3384 684508 418896 684536
rect 3384 684496 3390 684508
rect 418890 684496 418896 684508
rect 418948 684496 418954 684548
rect 266354 683748 266360 683800
rect 266412 683788 266418 683800
rect 446858 683788 446864 683800
rect 266412 683760 446864 683788
rect 266412 683748 266418 683760
rect 446858 683748 446864 683760
rect 446916 683748 446922 683800
rect 20806 683544 20812 683596
rect 20864 683584 20870 683596
rect 359458 683584 359464 683596
rect 20864 683556 359464 683584
rect 20864 683544 20870 683556
rect 359458 683544 359464 683556
rect 359516 683544 359522 683596
rect 21358 683476 21364 683528
rect 21416 683516 21422 683528
rect 416130 683516 416136 683528
rect 21416 683488 416136 683516
rect 21416 683476 21422 683488
rect 416130 683476 416136 683488
rect 416188 683476 416194 683528
rect 3878 683408 3884 683460
rect 3936 683448 3942 683460
rect 419166 683448 419172 683460
rect 3936 683420 419172 683448
rect 3936 683408 3942 683420
rect 419166 683408 419172 683420
rect 419224 683408 419230 683460
rect 3510 683340 3516 683392
rect 3568 683380 3574 683392
rect 419258 683380 419264 683392
rect 3568 683352 419264 683380
rect 3568 683340 3574 683352
rect 419258 683340 419264 683352
rect 419316 683340 419322 683392
rect 4062 683272 4068 683324
rect 4120 683312 4126 683324
rect 420178 683312 420184 683324
rect 4120 683284 420184 683312
rect 4120 683272 4126 683284
rect 420178 683272 420184 683284
rect 420236 683272 420242 683324
rect 3786 683204 3792 683256
rect 3844 683244 3850 683256
rect 445386 683244 445392 683256
rect 3844 683216 445392 683244
rect 3844 683204 3850 683216
rect 445386 683204 445392 683216
rect 445444 683204 445450 683256
rect 3234 683136 3240 683188
rect 3292 683176 3298 683188
rect 445478 683176 445484 683188
rect 3292 683148 445484 683176
rect 3292 683136 3298 683148
rect 445478 683136 445484 683148
rect 445536 683136 445542 683188
rect 3142 682660 3148 682712
rect 3200 682700 3206 682712
rect 420546 682700 420552 682712
rect 3200 682672 420552 682700
rect 3200 682660 3206 682672
rect 420546 682660 420552 682672
rect 420604 682660 420610 682712
rect 20070 681708 20076 681760
rect 20128 681748 20134 681760
rect 20806 681748 20812 681760
rect 20128 681720 20812 681748
rect 20128 681708 20134 681720
rect 20806 681708 20812 681720
rect 20864 681708 20870 681760
rect 3510 679192 3516 679244
rect 3568 679192 3574 679244
rect 3528 679040 3556 679192
rect 3510 678988 3516 679040
rect 3568 678988 3574 679040
rect 361758 678988 361764 679040
rect 361816 679028 361822 679040
rect 365070 679028 365076 679040
rect 361816 679000 365076 679028
rect 361816 678988 361822 679000
rect 365070 678988 365076 679000
rect 365128 678988 365134 679040
rect 3694 678512 3700 678564
rect 3752 678552 3758 678564
rect 3752 678524 3924 678552
rect 3752 678512 3758 678524
rect 3896 678224 3924 678524
rect 3878 678172 3884 678224
rect 3936 678172 3942 678224
rect 17678 670692 17684 670744
rect 17736 670732 17742 670744
rect 20070 670732 20076 670744
rect 17736 670704 20076 670732
rect 17736 670692 17742 670704
rect 20070 670692 20076 670704
rect 20128 670692 20134 670744
rect 450630 669944 450636 669996
rect 450688 669984 450694 669996
rect 462314 669984 462320 669996
rect 450688 669956 462320 669984
rect 450688 669944 450694 669956
rect 462314 669944 462320 669956
rect 462372 669944 462378 669996
rect 361758 667904 361764 667956
rect 361816 667944 361822 667956
rect 381538 667944 381544 667956
rect 361816 667916 381544 667944
rect 361816 667904 361822 667916
rect 381538 667904 381544 667916
rect 381596 667904 381602 667956
rect 13814 667360 13820 667412
rect 13872 667400 13878 667412
rect 17678 667400 17684 667412
rect 13872 667372 17684 667400
rect 13872 667360 13878 667372
rect 17678 667360 17684 667372
rect 17736 667360 17742 667412
rect 13814 665224 13820 665236
rect 12452 665196 13820 665224
rect 11790 665116 11796 665168
rect 11848 665156 11854 665168
rect 12452 665156 12480 665196
rect 13814 665184 13820 665196
rect 13872 665184 13878 665236
rect 11848 665128 12480 665156
rect 11848 665116 11854 665128
rect 11790 659716 11796 659728
rect 8312 659688 11796 659716
rect 7558 659608 7564 659660
rect 7616 659648 7622 659660
rect 8312 659648 8340 659688
rect 11790 659676 11796 659688
rect 11848 659676 11854 659728
rect 7616 659620 8340 659648
rect 7616 659608 7622 659620
rect 3142 658180 3148 658232
rect 3200 658220 3206 658232
rect 19978 658220 19984 658232
rect 3200 658192 19984 658220
rect 3200 658180 3206 658192
rect 19978 658180 19984 658192
rect 20036 658180 20042 658232
rect 361758 656888 361764 656940
rect 361816 656928 361822 656940
rect 406378 656928 406384 656940
rect 361816 656900 406384 656928
rect 361816 656888 361822 656900
rect 406378 656888 406384 656900
rect 406436 656888 406442 656940
rect 6178 655528 6184 655580
rect 6236 655568 6242 655580
rect 7558 655568 7564 655580
rect 6236 655540 7564 655568
rect 6236 655528 6242 655540
rect 7558 655528 7564 655540
rect 7616 655528 7622 655580
rect 4798 652740 4804 652792
rect 4856 652780 4862 652792
rect 6178 652780 6184 652792
rect 4856 652752 6184 652780
rect 4856 652740 4862 652752
rect 6178 652740 6184 652752
rect 6236 652740 6242 652792
rect 361758 645872 361764 645924
rect 361816 645912 361822 645924
rect 378778 645912 378784 645924
rect 361816 645884 378784 645912
rect 361816 645872 361822 645884
rect 378778 645872 378784 645884
rect 378836 645872 378842 645924
rect 569218 643084 569224 643136
rect 569276 643124 569282 643136
rect 579614 643124 579620 643136
rect 569276 643096 579620 643124
rect 569276 643084 569282 643096
rect 579614 643084 579620 643096
rect 579672 643084 579678 643136
rect 361574 634788 361580 634840
rect 361632 634828 361638 634840
rect 407758 634828 407764 634840
rect 361632 634800 407764 634828
rect 361632 634788 361638 634800
rect 407758 634788 407764 634800
rect 407816 634788 407822 634840
rect 3694 631320 3700 631372
rect 3752 631360 3758 631372
rect 20898 631360 20904 631372
rect 3752 631332 20904 631360
rect 3752 631320 3758 631332
rect 20898 631320 20904 631332
rect 20956 631320 20962 631372
rect 567838 630640 567844 630692
rect 567896 630680 567902 630692
rect 580166 630680 580172 630692
rect 567896 630652 580172 630680
rect 567896 630640 567902 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 361574 623772 361580 623824
rect 361632 623812 361638 623824
rect 376018 623812 376024 623824
rect 361632 623784 376024 623812
rect 361632 623772 361638 623784
rect 376018 623772 376024 623784
rect 376076 623772 376082 623824
rect 571978 616836 571984 616888
rect 572036 616876 572042 616888
rect 580166 616876 580172 616888
rect 572036 616848 580172 616876
rect 572036 616836 572042 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 359458 616768 359464 616820
rect 359516 616808 359522 616820
rect 360930 616808 360936 616820
rect 359516 616780 360936 616808
rect 359516 616768 359522 616780
rect 360930 616768 360936 616780
rect 360988 616768 360994 616820
rect 361574 612756 361580 612808
rect 361632 612796 361638 612808
rect 410518 612796 410524 612808
rect 361632 612768 410524 612796
rect 361632 612756 361638 612768
rect 410518 612756 410524 612768
rect 410576 612756 410582 612808
rect 360930 611192 360936 611244
rect 360988 611232 360994 611244
rect 362218 611232 362224 611244
rect 360988 611204 362224 611232
rect 360988 611192 360994 611204
rect 362218 611192 362224 611204
rect 362276 611192 362282 611244
rect 458726 603712 458732 603764
rect 458784 603752 458790 603764
rect 459002 603752 459008 603764
rect 458784 603724 459008 603752
rect 458784 603712 458790 603724
rect 459002 603712 459008 603724
rect 459060 603712 459066 603764
rect 361758 601672 361764 601724
rect 361816 601712 361822 601724
rect 374638 601712 374644 601724
rect 361816 601684 374644 601712
rect 361816 601672 361822 601684
rect 374638 601672 374644 601684
rect 374696 601672 374702 601724
rect 362218 600244 362224 600296
rect 362276 600284 362282 600296
rect 362954 600284 362960 600296
rect 362276 600256 362960 600284
rect 362276 600244 362282 600256
rect 362954 600244 362960 600256
rect 363012 600244 363018 600296
rect 457622 600244 457628 600296
rect 457680 600284 457686 600296
rect 461578 600284 461584 600296
rect 457680 600256 461584 600284
rect 457680 600244 457686 600256
rect 461578 600244 461584 600256
rect 461636 600244 461642 600296
rect 459002 599836 459008 599888
rect 459060 599876 459066 599888
rect 463694 599876 463700 599888
rect 459060 599848 463700 599876
rect 459060 599836 459066 599848
rect 463694 599836 463700 599848
rect 463752 599836 463758 599888
rect 458818 599700 458824 599752
rect 458876 599740 458882 599752
rect 465074 599740 465080 599752
rect 458876 599712 465080 599740
rect 458876 599700 458882 599712
rect 465074 599700 465080 599712
rect 465132 599700 465138 599752
rect 457530 599632 457536 599684
rect 457588 599672 457594 599684
rect 469858 599672 469864 599684
rect 457588 599644 469864 599672
rect 457588 599632 457594 599644
rect 469858 599632 469864 599644
rect 469916 599632 469922 599684
rect 457438 599564 457444 599616
rect 457496 599604 457502 599616
rect 469950 599604 469956 599616
rect 457496 599576 469956 599604
rect 457496 599564 457502 599576
rect 469950 599564 469956 599576
rect 470008 599564 470014 599616
rect 459922 598408 459928 598460
rect 459980 598448 459986 598460
rect 463786 598448 463792 598460
rect 459980 598420 463792 598448
rect 459980 598408 459986 598420
rect 463786 598408 463792 598420
rect 463844 598408 463850 598460
rect 458634 598340 458640 598392
rect 458692 598380 458698 598392
rect 465166 598380 465172 598392
rect 458692 598352 465172 598380
rect 458692 598340 458698 598352
rect 465166 598340 465172 598352
rect 465224 598340 465230 598392
rect 488626 598340 488632 598392
rect 488684 598380 488690 598392
rect 494238 598380 494244 598392
rect 488684 598352 494244 598380
rect 488684 598340 488690 598352
rect 494238 598340 494244 598352
rect 494296 598340 494302 598392
rect 449894 598272 449900 598324
rect 449952 598312 449958 598324
rect 526714 598312 526720 598324
rect 449952 598284 526720 598312
rect 449952 598272 449958 598284
rect 526714 598272 526720 598284
rect 526772 598272 526778 598324
rect 457898 598204 457904 598256
rect 457956 598244 457962 598256
rect 468478 598244 468484 598256
rect 457956 598216 468484 598244
rect 457956 598204 457962 598216
rect 468478 598204 468484 598216
rect 468536 598204 468542 598256
rect 482278 598204 482284 598256
rect 482336 598244 482342 598256
rect 494054 598244 494060 598256
rect 482336 598216 494060 598244
rect 482336 598204 482342 598216
rect 494054 598204 494060 598216
rect 494112 598204 494118 598256
rect 493318 598136 493324 598188
rect 493376 598176 493382 598188
rect 494974 598176 494980 598188
rect 493376 598148 494980 598176
rect 493376 598136 493382 598148
rect 494974 598136 494980 598148
rect 495032 598136 495038 598188
rect 519538 598136 519544 598188
rect 519596 598176 519602 598188
rect 520366 598176 520372 598188
rect 519596 598148 520372 598176
rect 519596 598136 519602 598148
rect 520366 598136 520372 598148
rect 520424 598136 520430 598188
rect 473262 598068 473268 598120
rect 473320 598108 473326 598120
rect 475930 598108 475936 598120
rect 473320 598080 475936 598108
rect 473320 598068 473326 598080
rect 475930 598068 475936 598080
rect 475988 598068 475994 598120
rect 457346 596844 457352 596896
rect 457404 596884 457410 596896
rect 465718 596884 465724 596896
rect 457404 596856 465724 596884
rect 457404 596844 457410 596856
rect 465718 596844 465724 596856
rect 465776 596844 465782 596896
rect 362954 596776 362960 596828
rect 363012 596816 363018 596828
rect 368382 596816 368388 596828
rect 363012 596788 368388 596816
rect 363012 596776 363018 596788
rect 368382 596776 368388 596788
rect 368440 596776 368446 596828
rect 449802 596776 449808 596828
rect 449860 596816 449866 596828
rect 469582 596816 469588 596828
rect 449860 596788 469588 596816
rect 449860 596776 449866 596788
rect 469582 596776 469588 596788
rect 469640 596776 469646 596828
rect 361758 590656 361764 590708
rect 361816 590696 361822 590708
rect 371970 590696 371976 590708
rect 361816 590668 371976 590696
rect 361816 590656 361822 590668
rect 371970 590656 371976 590668
rect 372028 590656 372034 590708
rect 567930 590656 567936 590708
rect 567988 590696 567994 590708
rect 580166 590696 580172 590708
rect 567988 590668 580172 590696
rect 567988 590656 567994 590668
rect 580166 590656 580172 590668
rect 580224 590656 580230 590708
rect 368474 589296 368480 589348
rect 368532 589336 368538 589348
rect 368532 589308 371280 589336
rect 368532 589296 368538 589308
rect 371252 589268 371280 589308
rect 372798 589268 372804 589280
rect 371252 589240 372804 589268
rect 372798 589228 372804 589240
rect 372856 589228 372862 589280
rect 372798 584400 372804 584452
rect 372856 584440 372862 584452
rect 379514 584440 379520 584452
rect 372856 584412 379520 584440
rect 372856 584400 372862 584412
rect 379514 584400 379520 584412
rect 379572 584400 379578 584452
rect 379514 582632 379520 582684
rect 379572 582672 379578 582684
rect 381630 582672 381636 582684
rect 379572 582644 381636 582672
rect 379572 582632 379578 582644
rect 381630 582632 381636 582644
rect 381688 582632 381694 582684
rect 361758 579640 361764 579692
rect 361816 579680 361822 579692
rect 370498 579680 370504 579692
rect 361816 579652 370504 579680
rect 361816 579640 361822 579652
rect 370498 579640 370504 579652
rect 370556 579640 370562 579692
rect 361758 568556 361764 568608
rect 361816 568596 361822 568608
rect 367738 568596 367744 568608
rect 361816 568568 367744 568596
rect 361816 568556 361822 568568
rect 367738 568556 367744 568568
rect 367796 568556 367802 568608
rect 459646 564340 459652 564392
rect 459704 564380 459710 564392
rect 462314 564380 462320 564392
rect 459704 564352 462320 564380
rect 459704 564340 459710 564352
rect 462314 564340 462320 564352
rect 462372 564340 462378 564392
rect 577498 563048 577504 563100
rect 577556 563088 577562 563100
rect 579614 563088 579620 563100
rect 577556 563060 579620 563088
rect 577556 563048 577562 563060
rect 579614 563048 579620 563060
rect 579672 563048 579678 563100
rect 381630 559308 381636 559360
rect 381688 559348 381694 559360
rect 383746 559348 383752 559360
rect 381688 559320 383752 559348
rect 381688 559308 381694 559320
rect 383746 559308 383752 559320
rect 383804 559308 383810 559360
rect 361574 557744 361580 557796
rect 361632 557784 361638 557796
rect 363598 557784 363604 557796
rect 361632 557756 363604 557784
rect 361632 557744 361638 557756
rect 363598 557744 363604 557756
rect 363656 557744 363662 557796
rect 383746 554140 383752 554192
rect 383804 554180 383810 554192
rect 385678 554180 385684 554192
rect 383804 554152 385684 554180
rect 383804 554140 383810 554152
rect 385678 554140 385684 554152
rect 385736 554140 385742 554192
rect 385678 550536 385684 550588
rect 385736 550576 385742 550588
rect 387426 550576 387432 550588
rect 385736 550548 387432 550576
rect 385736 550536 385742 550548
rect 387426 550536 387432 550548
rect 387484 550536 387490 550588
rect 361574 546592 361580 546644
rect 361632 546632 361638 546644
rect 363690 546632 363696 546644
rect 361632 546604 363696 546632
rect 361632 546592 361638 546604
rect 363690 546592 363696 546604
rect 363748 546592 363754 546644
rect 387426 546456 387432 546508
rect 387484 546496 387490 546508
rect 388438 546496 388444 546508
rect 387484 546468 388444 546496
rect 387484 546456 387490 546468
rect 388438 546456 388444 546468
rect 388496 546456 388502 546508
rect 457714 543056 457720 543108
rect 457772 543096 457778 543108
rect 464338 543096 464344 543108
rect 457772 543068 464344 543096
rect 457772 543056 457778 543068
rect 464338 543056 464344 543068
rect 464396 543056 464402 543108
rect 459830 542988 459836 543040
rect 459888 543028 459894 543040
rect 466454 543028 466460 543040
rect 459888 543000 466460 543028
rect 459888 542988 459894 543000
rect 466454 542988 466460 543000
rect 466512 542988 466518 543040
rect 361574 535712 361580 535764
rect 361632 535752 361638 535764
rect 363782 535752 363788 535764
rect 361632 535724 363788 535752
rect 361632 535712 361638 535724
rect 363782 535712 363788 535724
rect 363840 535712 363846 535764
rect 388438 535440 388444 535492
rect 388496 535480 388502 535492
rect 389818 535480 389824 535492
rect 388496 535452 389824 535480
rect 388496 535440 388502 535452
rect 389818 535440 389824 535452
rect 389876 535440 389882 535492
rect 448330 526396 448336 526448
rect 448388 526436 448394 526448
rect 500954 526436 500960 526448
rect 448388 526408 500960 526436
rect 448388 526396 448394 526408
rect 500954 526396 500960 526408
rect 501012 526396 501018 526448
rect 389818 524492 389824 524544
rect 389876 524532 389882 524544
rect 391198 524532 391204 524544
rect 389876 524504 391204 524532
rect 389876 524492 389882 524504
rect 391198 524492 391204 524504
rect 391256 524492 391262 524544
rect 361758 524424 361764 524476
rect 361816 524464 361822 524476
rect 411898 524464 411904 524476
rect 361816 524436 411904 524464
rect 361816 524424 361822 524436
rect 411898 524424 411904 524436
rect 411956 524424 411962 524476
rect 515398 524424 515404 524476
rect 515456 524464 515462 524476
rect 580166 524464 580172 524476
rect 515456 524436 580172 524464
rect 515456 524424 515462 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 448238 522248 448244 522300
rect 448296 522288 448302 522300
rect 493318 522288 493324 522300
rect 448296 522260 493324 522288
rect 448296 522248 448302 522260
rect 493318 522248 493324 522260
rect 493376 522248 493382 522300
rect 448422 520888 448428 520940
rect 448480 520928 448486 520940
rect 506474 520928 506480 520940
rect 448480 520900 506480 520928
rect 448480 520888 448486 520900
rect 506474 520888 506480 520900
rect 506532 520888 506538 520940
rect 462958 520412 462964 520464
rect 463016 520452 463022 520464
rect 488626 520452 488632 520464
rect 463016 520424 488632 520452
rect 463016 520412 463022 520424
rect 488626 520412 488632 520424
rect 488684 520412 488690 520464
rect 472894 520344 472900 520396
rect 472952 520384 472958 520396
rect 473262 520384 473268 520396
rect 472952 520356 473268 520384
rect 472952 520344 472958 520356
rect 473262 520344 473268 520356
rect 473320 520384 473326 520396
rect 494238 520384 494244 520396
rect 473320 520356 494244 520384
rect 473320 520344 473326 520356
rect 494238 520344 494244 520356
rect 494296 520344 494302 520396
rect 458082 520004 458088 520056
rect 458140 520044 458146 520056
rect 463050 520044 463056 520056
rect 458140 520016 463056 520044
rect 458140 520004 458146 520016
rect 463050 520004 463056 520016
rect 463108 520004 463114 520056
rect 457254 519596 457260 519648
rect 457312 519636 457318 519648
rect 467926 519636 467932 519648
rect 457312 519608 467932 519636
rect 457312 519596 457318 519608
rect 467926 519596 467932 519608
rect 467984 519596 467990 519648
rect 448054 519528 448060 519580
rect 448112 519568 448118 519580
rect 472894 519568 472900 519580
rect 448112 519540 472900 519568
rect 448112 519528 448118 519540
rect 472894 519528 472900 519540
rect 472952 519528 472958 519580
rect 459738 518712 459744 518764
rect 459796 518752 459802 518764
rect 462498 518752 462504 518764
rect 459796 518724 462504 518752
rect 459796 518712 459802 518724
rect 462498 518712 462504 518724
rect 462556 518712 462562 518764
rect 457806 518372 457812 518424
rect 457864 518412 457870 518424
rect 466546 518412 466552 518424
rect 457864 518384 466552 518412
rect 457864 518372 457870 518384
rect 466546 518372 466552 518384
rect 466604 518372 466610 518424
rect 459554 518304 459560 518356
rect 459612 518344 459618 518356
rect 470686 518344 470692 518356
rect 459612 518316 470692 518344
rect 459612 518304 459618 518316
rect 470686 518304 470692 518316
rect 470744 518304 470750 518356
rect 459094 518236 459100 518288
rect 459152 518276 459158 518288
rect 470870 518276 470876 518288
rect 459152 518248 470876 518276
rect 459152 518236 459158 518248
rect 470870 518236 470876 518248
rect 470928 518236 470934 518288
rect 447962 518168 447968 518220
rect 448020 518208 448026 518220
rect 462406 518208 462412 518220
rect 448020 518180 462412 518208
rect 448020 518168 448026 518180
rect 462406 518168 462412 518180
rect 462464 518168 462470 518220
rect 457990 517964 457996 518016
rect 458048 518004 458054 518016
rect 461670 518004 461676 518016
rect 458048 517976 461676 518004
rect 458048 517964 458054 517976
rect 461670 517964 461676 517976
rect 461728 517964 461734 518016
rect 391198 517488 391204 517540
rect 391256 517528 391262 517540
rect 391256 517500 393314 517528
rect 391256 517488 391262 517500
rect 393286 517460 393314 517500
rect 480162 517488 480168 517540
rect 480220 517528 480226 517540
rect 482646 517528 482652 517540
rect 480220 517500 482652 517528
rect 480220 517488 480226 517500
rect 482646 517488 482652 517500
rect 482704 517488 482710 517540
rect 394602 517460 394608 517472
rect 393286 517432 394608 517460
rect 394602 517420 394608 517432
rect 394660 517420 394666 517472
rect 448422 516128 448428 516180
rect 448480 516168 448486 516180
rect 491846 516168 491852 516180
rect 448480 516140 491852 516168
rect 448480 516128 448486 516140
rect 491846 516128 491852 516140
rect 491904 516128 491910 516180
rect 494054 515380 494060 515432
rect 494112 515420 494118 515432
rect 538214 515420 538220 515432
rect 494112 515392 538220 515420
rect 494112 515380 494118 515392
rect 538214 515380 538220 515392
rect 538272 515380 538278 515432
rect 3970 514768 3976 514820
rect 4028 514808 4034 514820
rect 4798 514808 4804 514820
rect 4028 514780 4804 514808
rect 4028 514768 4034 514780
rect 4798 514768 4804 514780
rect 4856 514768 4862 514820
rect 361758 513340 361764 513392
rect 361816 513380 361822 513392
rect 414658 513380 414664 513392
rect 361816 513352 414664 513380
rect 361816 513340 361822 513352
rect 414658 513340 414664 513352
rect 414716 513340 414722 513392
rect 494054 511980 494060 512032
rect 494112 512020 494118 512032
rect 535454 512020 535460 512032
rect 494112 511992 535460 512020
rect 494112 511980 494118 511992
rect 535454 511980 535460 511992
rect 535512 511980 535518 512032
rect 394694 510620 394700 510672
rect 394752 510660 394758 510672
rect 394752 510632 398880 510660
rect 394752 510620 394758 510632
rect 398852 510592 398880 510632
rect 402238 510592 402244 510604
rect 398852 510564 402244 510592
rect 402238 510552 402244 510564
rect 402296 510552 402302 510604
rect 494238 508512 494244 508564
rect 494296 508552 494302 508564
rect 532694 508552 532700 508564
rect 494296 508524 532700 508552
rect 494296 508512 494302 508524
rect 532694 508512 532700 508524
rect 532752 508512 532758 508564
rect 494974 505112 494980 505164
rect 495032 505152 495038 505164
rect 529934 505152 529940 505164
rect 495032 505124 529940 505152
rect 495032 505112 495038 505124
rect 529934 505112 529940 505124
rect 529992 505112 529998 505164
rect 361758 502324 361764 502376
rect 361816 502364 361822 502376
rect 416314 502364 416320 502376
rect 361816 502336 416320 502364
rect 361816 502324 361822 502336
rect 416314 502324 416320 502336
rect 416372 502324 416378 502376
rect 448514 500216 448520 500268
rect 448572 500256 448578 500268
rect 545114 500256 545120 500268
rect 448572 500228 545120 500256
rect 448572 500216 448578 500228
rect 545114 500216 545120 500228
rect 545172 500216 545178 500268
rect 450078 499808 450084 499860
rect 450136 499848 450142 499860
rect 450722 499848 450728 499860
rect 450136 499820 450728 499848
rect 450136 499808 450142 499820
rect 450722 499808 450728 499820
rect 450780 499808 450786 499860
rect 447318 499536 447324 499588
rect 447376 499576 447382 499588
rect 449710 499576 449716 499588
rect 447376 499548 449716 499576
rect 447376 499536 447382 499548
rect 449710 499536 449716 499548
rect 449768 499536 449774 499588
rect 447870 499468 447876 499520
rect 447928 499508 447934 499520
rect 494054 499508 494060 499520
rect 447928 499480 494060 499508
rect 447928 499468 447934 499480
rect 494054 499468 494060 499480
rect 494112 499468 494118 499520
rect 447962 499400 447968 499452
rect 448020 499440 448026 499452
rect 494146 499440 494152 499452
rect 448020 499412 494152 499440
rect 448020 499400 448026 499412
rect 494146 499400 494152 499412
rect 494204 499400 494210 499452
rect 448238 498856 448244 498908
rect 448296 498896 448302 498908
rect 542446 498896 542452 498908
rect 448296 498868 542452 498896
rect 448296 498856 448302 498868
rect 542446 498856 542452 498868
rect 542504 498856 542510 498908
rect 449710 498788 449716 498840
rect 449768 498828 449774 498840
rect 547874 498828 547880 498840
rect 449768 498800 547880 498828
rect 449768 498788 449774 498800
rect 547874 498788 547880 498800
rect 547932 498788 547938 498840
rect 452010 497564 452016 497616
rect 452068 497604 452074 497616
rect 481634 497604 481640 497616
rect 452068 497576 481640 497604
rect 452068 497564 452074 497576
rect 481634 497564 481640 497576
rect 481692 497564 481698 497616
rect 449802 497496 449808 497548
rect 449860 497536 449866 497548
rect 486234 497536 486240 497548
rect 449860 497508 486240 497536
rect 449860 497496 449866 497508
rect 486234 497496 486240 497508
rect 486292 497496 486298 497548
rect 451918 497428 451924 497480
rect 451976 497468 451982 497480
rect 488626 497468 488632 497480
rect 451976 497440 488632 497468
rect 451976 497428 451982 497440
rect 488626 497428 488632 497440
rect 488684 497428 488690 497480
rect 454034 497088 454040 497140
rect 454092 497128 454098 497140
rect 459554 497128 459560 497140
rect 454092 497100 459560 497128
rect 454092 497088 454098 497100
rect 459554 497088 459560 497100
rect 459612 497088 459618 497140
rect 454126 497020 454132 497072
rect 454184 497060 454190 497072
rect 458082 497060 458088 497072
rect 454184 497032 458088 497060
rect 454184 497020 454190 497032
rect 458082 497020 458088 497032
rect 458140 497020 458146 497072
rect 455414 496952 455420 497004
rect 455472 496992 455478 497004
rect 461026 496992 461032 497004
rect 455472 496964 461032 496992
rect 455472 496952 455478 496964
rect 461026 496952 461032 496964
rect 461084 496952 461090 497004
rect 452838 496884 452844 496936
rect 452896 496924 452902 496936
rect 455138 496924 455144 496936
rect 452896 496896 455144 496924
rect 452896 496884 452902 496896
rect 455138 496884 455144 496896
rect 455196 496884 455202 496936
rect 451366 496816 451372 496868
rect 451424 496856 451430 496868
rect 453666 496856 453672 496868
rect 451424 496828 453672 496856
rect 451424 496816 451430 496828
rect 453666 496816 453672 496828
rect 453724 496816 453730 496868
rect 454678 496816 454684 496868
rect 454736 496856 454742 496868
rect 456610 496856 456616 496868
rect 454736 496828 456616 496856
rect 454736 496816 454742 496828
rect 456610 496816 456616 496828
rect 456668 496816 456674 496868
rect 569310 484372 569316 484424
rect 569368 484412 569374 484424
rect 580166 484412 580172 484424
rect 569368 484384 580172 484412
rect 569368 484372 569374 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 361758 480224 361764 480276
rect 361816 480264 361822 480276
rect 418706 480264 418712 480276
rect 361816 480236 418712 480264
rect 361816 480224 361822 480236
rect 418706 480224 418712 480236
rect 418764 480224 418770 480276
rect 511258 470568 511264 470620
rect 511316 470608 511322 470620
rect 579982 470608 579988 470620
rect 511316 470580 579988 470608
rect 511316 470568 511322 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 402238 469276 402244 469328
rect 402296 469316 402302 469328
rect 404998 469316 405004 469328
rect 402296 469288 405004 469316
rect 402296 469276 402302 469288
rect 404998 469276 405004 469288
rect 405056 469276 405062 469328
rect 361758 469208 361764 469260
rect 361816 469248 361822 469260
rect 417418 469248 417424 469260
rect 361816 469220 417424 469248
rect 361816 469208 361822 469220
rect 417418 469208 417424 469220
rect 417476 469208 417482 469260
rect 494698 462476 494704 462528
rect 494756 462516 494762 462528
rect 527634 462516 527640 462528
rect 494756 462488 527640 462516
rect 494756 462476 494762 462488
rect 527634 462476 527640 462488
rect 527692 462476 527698 462528
rect 436094 462408 436100 462460
rect 436152 462448 436158 462460
rect 554130 462448 554136 462460
rect 436152 462420 554136 462448
rect 436152 462408 436158 462420
rect 554130 462408 554136 462420
rect 554188 462408 554194 462460
rect 433242 462340 433248 462392
rect 433300 462380 433306 462392
rect 551186 462380 551192 462392
rect 433300 462352 551192 462380
rect 433300 462340 433306 462352
rect 551186 462340 551192 462352
rect 551244 462340 551250 462392
rect 515490 461660 515496 461712
rect 515548 461700 515554 461712
rect 542354 461700 542360 461712
rect 515548 461672 542360 461700
rect 515548 461660 515554 461672
rect 542354 461660 542360 461672
rect 542412 461660 542418 461712
rect 480162 461592 480168 461644
rect 480220 461632 480226 461644
rect 521746 461632 521752 461644
rect 480220 461604 521752 461632
rect 480220 461592 480226 461604
rect 521746 461592 521752 461604
rect 521804 461592 521810 461644
rect 449986 460912 449992 460964
rect 450044 460952 450050 460964
rect 524414 460952 524420 460964
rect 450044 460924 524420 460952
rect 450044 460912 450050 460924
rect 524414 460912 524420 460924
rect 524472 460912 524478 460964
rect 361758 458192 361764 458244
rect 361816 458232 361822 458244
rect 382918 458232 382924 458244
rect 361816 458204 382924 458232
rect 361816 458192 361822 458204
rect 382918 458192 382924 458204
rect 382976 458192 382982 458244
rect 449434 457444 449440 457496
rect 449492 457484 449498 457496
rect 487154 457484 487160 457496
rect 449492 457456 487160 457484
rect 449492 457444 449498 457456
rect 487154 457444 487160 457456
rect 487212 457444 487218 457496
rect 473722 456764 473728 456816
rect 473780 456804 473786 456816
rect 480162 456804 480168 456816
rect 473780 456776 480168 456804
rect 473780 456764 473786 456776
rect 480162 456764 480168 456776
rect 480220 456764 480226 456816
rect 449526 456016 449532 456068
rect 449584 456056 449590 456068
rect 484394 456056 484400 456068
rect 449584 456028 484400 456056
rect 449584 456016 449590 456028
rect 484394 456016 484400 456028
rect 484452 456016 484458 456068
rect 488258 456016 488264 456068
rect 488316 456056 488322 456068
rect 494698 456056 494704 456068
rect 488316 456028 494704 456056
rect 488316 456016 488322 456028
rect 494698 456016 494704 456028
rect 494756 456016 494762 456068
rect 450170 455472 450176 455524
rect 450228 455512 450234 455524
rect 480990 455512 480996 455524
rect 450228 455484 480996 455512
rect 450228 455472 450234 455484
rect 480990 455472 480996 455484
rect 481048 455472 481054 455524
rect 422294 455404 422300 455456
rect 422352 455444 422358 455456
rect 473722 455444 473728 455456
rect 422352 455416 473728 455444
rect 422352 455404 422358 455416
rect 473722 455404 473728 455416
rect 473780 455404 473786 455456
rect 404998 455336 405004 455388
rect 405056 455376 405062 455388
rect 406470 455376 406476 455388
rect 405056 455348 406476 455376
rect 405056 455336 405062 455348
rect 406470 455336 406476 455348
rect 406528 455336 406534 455388
rect 450262 454792 450268 454844
rect 450320 454832 450326 454844
rect 480254 454832 480260 454844
rect 450320 454804 480260 454832
rect 450320 454792 450326 454804
rect 480254 454792 480260 454804
rect 480312 454792 480318 454844
rect 449710 454724 449716 454776
rect 449768 454764 449774 454776
rect 481910 454764 481916 454776
rect 449768 454736 481916 454764
rect 449768 454724 449774 454736
rect 481910 454724 481916 454736
rect 481968 454724 481974 454776
rect 449618 454656 449624 454708
rect 449676 454696 449682 454708
rect 483106 454696 483112 454708
rect 449676 454668 483112 454696
rect 449676 454656 449682 454668
rect 483106 454656 483112 454668
rect 483164 454656 483170 454708
rect 406470 450916 406476 450968
rect 406528 450956 406534 450968
rect 408494 450956 408500 450968
rect 406528 450928 408500 450956
rect 406528 450916 406534 450928
rect 408494 450916 408500 450928
rect 408552 450916 408558 450968
rect 427446 447108 427452 447160
rect 427504 447148 427510 447160
rect 446950 447148 446956 447160
rect 427504 447120 446956 447148
rect 427504 447108 427510 447120
rect 446950 447108 446956 447120
rect 447008 447108 447014 447160
rect 432414 445748 432420 445800
rect 432472 445788 432478 445800
rect 433242 445788 433248 445800
rect 432472 445760 433248 445788
rect 432472 445748 432478 445760
rect 433242 445748 433248 445760
rect 433300 445788 433306 445800
rect 444098 445788 444104 445800
rect 433300 445760 444104 445788
rect 433300 445748 433306 445760
rect 444098 445748 444104 445760
rect 444156 445748 444162 445800
rect 436094 445680 436100 445732
rect 436152 445720 436158 445732
rect 437382 445720 437388 445732
rect 436152 445692 437388 445720
rect 436152 445680 436158 445692
rect 437382 445680 437388 445692
rect 437440 445680 437446 445732
rect 437290 444524 437296 444576
rect 437348 444564 437354 444576
rect 445846 444564 445852 444576
rect 437348 444536 445852 444564
rect 437348 444524 437354 444536
rect 445846 444524 445852 444536
rect 445904 444524 445910 444576
rect 442626 444456 442632 444508
rect 442684 444496 442690 444508
rect 445754 444496 445760 444508
rect 442684 444468 445760 444496
rect 442684 444456 442690 444468
rect 445754 444456 445760 444468
rect 445812 444456 445818 444508
rect 422754 444388 422760 444440
rect 422812 444428 422818 444440
rect 445570 444428 445576 444440
rect 422812 444400 445576 444428
rect 422812 444388 422818 444400
rect 445570 444388 445576 444400
rect 445628 444388 445634 444440
rect 408494 441600 408500 441652
rect 408552 441640 408558 441652
rect 408552 441612 411300 441640
rect 408552 441600 408558 441612
rect 411272 441572 411300 441612
rect 413738 441572 413744 441584
rect 411272 441544 413744 441572
rect 413738 441532 413744 441544
rect 413796 441532 413802 441584
rect 413738 437520 413744 437572
rect 413796 437560 413802 437572
rect 414750 437560 414756 437572
rect 413796 437532 414756 437560
rect 413796 437520 413802 437532
rect 414750 437520 414756 437532
rect 414808 437520 414814 437572
rect 361758 436092 361764 436144
rect 361816 436132 361822 436144
rect 418614 436132 418620 436144
rect 361816 436104 418620 436132
rect 361816 436092 361822 436104
rect 418614 436092 418620 436104
rect 418672 436092 418678 436144
rect 414750 431332 414756 431384
rect 414808 431372 414814 431384
rect 416682 431372 416688 431384
rect 414808 431344 416688 431372
rect 414808 431332 414814 431344
rect 416682 431332 416688 431344
rect 416740 431332 416746 431384
rect 569402 430584 569408 430636
rect 569460 430624 569466 430636
rect 580166 430624 580172 430636
rect 569460 430596 580172 430624
rect 569460 430584 569466 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 456886 429836 456892 429888
rect 456944 429876 456950 429888
rect 474274 429876 474280 429888
rect 456944 429848 474280 429876
rect 456944 429836 456950 429848
rect 474274 429836 474280 429848
rect 474332 429836 474338 429888
rect 478138 429156 478144 429208
rect 478196 429196 478202 429208
rect 479610 429196 479616 429208
rect 478196 429168 479616 429196
rect 478196 429156 478202 429168
rect 479610 429156 479616 429168
rect 479668 429156 479674 429208
rect 482278 429156 482284 429208
rect 482336 429196 482342 429208
rect 484946 429196 484952 429208
rect 482336 429168 484952 429196
rect 482336 429156 482342 429168
rect 484946 429156 484952 429168
rect 485004 429156 485010 429208
rect 486418 429156 486424 429208
rect 486476 429196 486482 429208
rect 487614 429196 487620 429208
rect 486476 429168 487620 429196
rect 486476 429156 486482 429168
rect 487614 429156 487620 429168
rect 487672 429156 487678 429208
rect 416682 429020 416688 429072
rect 416740 429060 416746 429072
rect 420362 429060 420368 429072
rect 416740 429032 420368 429060
rect 416740 429020 416746 429032
rect 420362 429020 420368 429032
rect 420420 429020 420426 429072
rect 457438 428408 457444 428460
rect 457496 428448 457502 428460
rect 471606 428448 471612 428460
rect 457496 428420 471612 428448
rect 457496 428408 457502 428420
rect 471606 428408 471612 428420
rect 471664 428408 471670 428460
rect 529198 423580 529204 423632
rect 529256 423620 529262 423632
rect 530210 423620 530216 423632
rect 529256 423592 530216 423620
rect 529256 423580 529262 423592
rect 530210 423580 530216 423592
rect 530268 423580 530274 423632
rect 530578 423580 530584 423632
rect 530636 423620 530642 423632
rect 532786 423620 532792 423632
rect 530636 423592 532792 423620
rect 530636 423580 530642 423592
rect 532786 423580 532792 423592
rect 532844 423580 532850 423632
rect 502978 423512 502984 423564
rect 503036 423552 503042 423564
rect 523770 423552 523776 423564
rect 503036 423524 523776 423552
rect 503036 423512 503042 423524
rect 523770 423512 523776 423524
rect 523828 423512 523834 423564
rect 522298 423444 522304 423496
rect 522356 423484 522362 423496
rect 549530 423484 549536 423496
rect 522356 423456 549536 423484
rect 522356 423444 522362 423456
rect 549530 423444 549536 423456
rect 549588 423444 549594 423496
rect 483014 423376 483020 423428
rect 483072 423416 483078 423428
rect 522482 423416 522488 423428
rect 483072 423388 522488 423416
rect 483072 423376 483078 423388
rect 522482 423376 522488 423388
rect 522540 423376 522546 423428
rect 523678 423376 523684 423428
rect 523736 423416 523742 423428
rect 552106 423416 552112 423428
rect 523736 423388 552112 423416
rect 523736 423376 523742 423388
rect 552106 423376 552112 423388
rect 552164 423376 552170 423428
rect 485774 423308 485780 423360
rect 485832 423348 485838 423360
rect 526346 423348 526352 423360
rect 485832 423320 526352 423348
rect 485832 423308 485838 423320
rect 526346 423308 526352 423320
rect 526404 423308 526410 423360
rect 526438 423308 526444 423360
rect 526496 423348 526502 423360
rect 554682 423348 554688 423360
rect 526496 423320 554688 423348
rect 526496 423308 526502 423320
rect 554682 423308 554688 423320
rect 554740 423308 554746 423360
rect 487154 423240 487160 423292
rect 487212 423280 487218 423292
rect 528922 423280 528928 423292
rect 487212 423252 528928 423280
rect 487212 423240 487218 423252
rect 528922 423240 528928 423252
rect 528980 423240 528986 423292
rect 488534 423172 488540 423224
rect 488592 423212 488598 423224
rect 531498 423212 531504 423224
rect 488592 423184 531504 423212
rect 488592 423172 488598 423184
rect 531498 423172 531504 423184
rect 531556 423172 531562 423224
rect 496814 423104 496820 423156
rect 496872 423144 496878 423156
rect 545666 423144 545672 423156
rect 496872 423116 545672 423144
rect 496872 423104 496878 423116
rect 545666 423104 545672 423116
rect 545724 423104 545730 423156
rect 498194 423036 498200 423088
rect 498252 423076 498258 423088
rect 548242 423076 548248 423088
rect 498252 423048 548248 423076
rect 498252 423036 498258 423048
rect 548242 423036 548248 423048
rect 548300 423036 548306 423088
rect 499574 422968 499580 423020
rect 499632 423008 499638 423020
rect 550818 423008 550824 423020
rect 499632 422980 550824 423008
rect 499632 422968 499638 422980
rect 550818 422968 550824 422980
rect 550876 422968 550882 423020
rect 501046 422900 501052 422952
rect 501104 422940 501110 422952
rect 553394 422940 553400 422952
rect 501104 422912 553400 422940
rect 501104 422900 501110 422912
rect 553394 422900 553400 422912
rect 553452 422900 553458 422952
rect 483106 421540 483112 421592
rect 483164 421580 483170 421592
rect 521194 421580 521200 421592
rect 483164 421552 521200 421580
rect 483164 421540 483170 421552
rect 521194 421540 521200 421552
rect 521252 421540 521258 421592
rect 494054 420180 494060 420232
rect 494112 420220 494118 420232
rect 541802 420220 541808 420232
rect 494112 420192 541808 420220
rect 494112 420180 494118 420192
rect 541802 420180 541808 420192
rect 541860 420180 541866 420232
rect 362402 418752 362408 418804
rect 362460 418792 362466 418804
rect 440878 418792 440884 418804
rect 362460 418764 440884 418792
rect 362460 418752 362466 418764
rect 440878 418752 440884 418764
rect 440936 418752 440942 418804
rect 420362 418140 420368 418192
rect 420420 418180 420426 418192
rect 420420 418152 422294 418180
rect 420420 418140 420426 418152
rect 422266 418112 422294 418152
rect 426434 418112 426440 418124
rect 422266 418084 426440 418112
rect 426434 418072 426440 418084
rect 426492 418072 426498 418124
rect 425974 417732 425980 417784
rect 426032 417772 426038 417784
rect 507854 417772 507860 417784
rect 426032 417744 507860 417772
rect 426032 417732 426038 417744
rect 507854 417732 507860 417744
rect 507912 417732 507918 417784
rect 421466 417664 421472 417716
rect 421524 417704 421530 417716
rect 503714 417704 503720 417716
rect 421524 417676 503720 417704
rect 421524 417664 421530 417676
rect 503714 417664 503720 417676
rect 503772 417664 503778 417716
rect 424686 417596 424692 417648
rect 424744 417636 424750 417648
rect 506474 417636 506480 417648
rect 424744 417608 506480 417636
rect 424744 417596 424750 417608
rect 506474 417596 506480 417608
rect 506532 417596 506538 417648
rect 424042 417528 424048 417580
rect 424100 417568 424106 417580
rect 506566 417568 506572 417580
rect 424100 417540 506572 417568
rect 424100 417528 424106 417540
rect 506566 417528 506572 417540
rect 506624 417528 506630 417580
rect 425330 417460 425336 417512
rect 425388 417500 425394 417512
rect 507946 417500 507952 417512
rect 425388 417472 507952 417500
rect 425388 417460 425394 417472
rect 507946 417460 507952 417472
rect 508004 417460 508010 417512
rect 422110 417392 422116 417444
rect 422168 417432 422174 417444
rect 503990 417432 503996 417444
rect 422168 417404 503996 417432
rect 422168 417392 422174 417404
rect 503990 417392 503996 417404
rect 504048 417392 504054 417444
rect 362310 416032 362316 416084
rect 362368 416072 362374 416084
rect 436738 416072 436744 416084
rect 362368 416044 436744 416072
rect 362368 416032 362374 416044
rect 436738 416032 436744 416044
rect 436796 416032 436802 416084
rect 426434 415624 426440 415676
rect 426492 415664 426498 415676
rect 429838 415664 429844 415676
rect 426492 415636 429844 415664
rect 426492 415624 426498 415636
rect 429838 415624 429844 415636
rect 429896 415624 429902 415676
rect 361574 413992 361580 414044
rect 361632 414032 361638 414044
rect 439498 414032 439504 414044
rect 361632 414004 439504 414032
rect 361632 413992 361638 414004
rect 439498 413992 439504 414004
rect 439556 413992 439562 414044
rect 429838 410184 429844 410236
rect 429896 410224 429902 410236
rect 431218 410224 431224 410236
rect 429896 410196 431224 410224
rect 429896 410184 429902 410196
rect 431218 410184 431224 410196
rect 431276 410184 431282 410236
rect 361574 402976 361580 403028
rect 361632 403016 361638 403028
rect 442258 403016 442264 403028
rect 361632 402988 442264 403016
rect 361632 402976 361638 402988
rect 442258 402976 442264 402988
rect 442316 402976 442322 403028
rect 502610 402228 502616 402280
rect 502668 402268 502674 402280
rect 557534 402268 557540 402280
rect 502668 402240 557540 402268
rect 502668 402228 502674 402240
rect 557534 402228 557540 402240
rect 557592 402228 557598 402280
rect 497458 400868 497464 400920
rect 497516 400908 497522 400920
rect 546494 400908 546500 400920
rect 497516 400880 546500 400908
rect 497516 400868 497522 400880
rect 546494 400868 546500 400880
rect 546552 400868 546558 400920
rect 494146 399440 494152 399492
rect 494204 399480 494210 399492
rect 539594 399480 539600 399492
rect 494204 399452 539600 399480
rect 494204 399440 494210 399452
rect 539594 399440 539600 399452
rect 539652 399440 539658 399492
rect 431218 398760 431224 398812
rect 431276 398800 431282 398812
rect 432598 398800 432604 398812
rect 431276 398772 432604 398800
rect 431276 398760 431282 398772
rect 432598 398760 432604 398772
rect 432656 398760 432662 398812
rect 492674 398080 492680 398132
rect 492732 398120 492738 398132
rect 538214 398120 538220 398132
rect 492732 398092 538220 398120
rect 492732 398080 492738 398092
rect 538214 398080 538220 398092
rect 538272 398080 538278 398132
rect 492766 396720 492772 396772
rect 492824 396760 492830 396772
rect 536834 396760 536840 396772
rect 492824 396732 536840 396760
rect 492824 396720 492830 396732
rect 536834 396720 536840 396732
rect 536892 396720 536898 396772
rect 461394 395292 461400 395344
rect 461452 395332 461458 395344
rect 490006 395332 490012 395344
rect 461452 395304 490012 395332
rect 461452 395292 461458 395304
rect 490006 395292 490012 395304
rect 490064 395292 490070 395344
rect 491570 395292 491576 395344
rect 491628 395332 491634 395344
rect 535454 395332 535460 395344
rect 491628 395304 535460 395332
rect 491628 395292 491634 395304
rect 535454 395292 535460 395304
rect 535512 395292 535518 395344
rect 458450 393932 458456 393984
rect 458508 393972 458514 393984
rect 478138 393972 478144 393984
rect 458508 393944 478144 393972
rect 458508 393932 458514 393944
rect 478138 393932 478144 393944
rect 478196 393932 478202 393984
rect 491386 393932 491392 393984
rect 491444 393972 491450 393984
rect 534166 393972 534172 393984
rect 491444 393944 534172 393972
rect 491444 393932 491450 393944
rect 534166 393932 534172 393944
rect 534224 393932 534230 393984
rect 458174 392640 458180 392692
rect 458232 392680 458238 392692
rect 476114 392680 476120 392692
rect 458232 392652 476120 392680
rect 458232 392640 458238 392652
rect 476114 392640 476120 392652
rect 476172 392640 476178 392692
rect 461118 392572 461124 392624
rect 461176 392612 461182 392624
rect 486418 392612 486424 392624
rect 461176 392584 486424 392612
rect 461176 392572 461182 392584
rect 486418 392572 486424 392584
rect 486476 392572 486482 392624
rect 490558 392572 490564 392624
rect 490616 392612 490622 392624
rect 534074 392612 534080 392624
rect 490616 392584 534080 392612
rect 490616 392572 490622 392584
rect 534074 392572 534080 392584
rect 534132 392572 534138 392624
rect 440970 392068 440976 392080
rect 431926 392040 440976 392068
rect 361574 391960 361580 392012
rect 361632 392000 361638 392012
rect 431926 392000 431954 392040
rect 440970 392028 440976 392040
rect 441028 392028 441034 392080
rect 361632 391972 431954 392000
rect 361632 391960 361638 391972
rect 432598 391960 432604 392012
rect 432656 392000 432662 392012
rect 433978 392000 433984 392012
rect 432656 391972 433984 392000
rect 432656 391960 432662 391972
rect 433978 391960 433984 391972
rect 434036 391960 434042 392012
rect 460382 391348 460388 391400
rect 460440 391388 460446 391400
rect 482278 391388 482284 391400
rect 460440 391360 482284 391388
rect 460440 391348 460446 391360
rect 482278 391348 482284 391360
rect 482336 391348 482342 391400
rect 450446 391280 450452 391332
rect 450504 391320 450510 391332
rect 491294 391320 491300 391332
rect 450504 391292 491300 391320
rect 450504 391280 450510 391292
rect 491294 391280 491300 391292
rect 491352 391280 491358 391332
rect 496446 391280 496452 391332
rect 496504 391320 496510 391332
rect 543734 391320 543740 391332
rect 496504 391292 543740 391320
rect 496504 391280 496510 391292
rect 543734 391280 543740 391292
rect 543792 391280 543798 391332
rect 422386 391212 422392 391264
rect 422444 391252 422450 391264
rect 506014 391252 506020 391264
rect 422444 391224 506020 391252
rect 422444 391212 422450 391224
rect 506014 391212 506020 391224
rect 506072 391212 506078 391264
rect 461670 389852 461676 389904
rect 461728 389892 461734 389904
rect 481634 389892 481640 389904
rect 461728 389864 481640 389892
rect 461728 389852 461734 389864
rect 481634 389852 481640 389864
rect 481692 389852 481698 389904
rect 495710 389852 495716 389904
rect 495768 389892 495774 389904
rect 542354 389892 542360 389904
rect 495768 389864 542360 389892
rect 495768 389852 495774 389864
rect 542354 389852 542360 389864
rect 542412 389852 542418 389904
rect 422294 389784 422300 389836
rect 422352 389824 422358 389836
rect 505278 389824 505284 389836
rect 422352 389796 505284 389824
rect 422352 389784 422358 389796
rect 505278 389784 505284 389796
rect 505336 389784 505342 389836
rect 450078 389240 450084 389292
rect 450136 389280 450142 389292
rect 450722 389280 450728 389292
rect 450136 389252 450728 389280
rect 450136 389240 450142 389252
rect 450722 389240 450728 389252
rect 450780 389240 450786 389292
rect 454034 389240 454040 389292
rect 454092 389280 454098 389292
rect 454862 389280 454868 389292
rect 454092 389252 454868 389280
rect 454092 389240 454098 389252
rect 454862 389240 454868 389252
rect 454920 389240 454926 389292
rect 465074 389240 465080 389292
rect 465132 389280 465138 389292
rect 465902 389280 465908 389292
rect 465132 389252 465908 389280
rect 465132 389240 465138 389252
rect 465902 389240 465908 389252
rect 465960 389240 465966 389292
rect 483014 389240 483020 389292
rect 483072 389280 483078 389292
rect 483566 389280 483572 389292
rect 483072 389252 483572 389280
rect 483072 389240 483078 389252
rect 483566 389240 483572 389252
rect 483624 389240 483630 389292
rect 492674 389240 492680 389292
rect 492732 389280 492738 389292
rect 493134 389280 493140 389292
rect 492732 389252 493140 389280
rect 492732 389240 492738 389252
rect 493134 389240 493140 389252
rect 493192 389240 493198 389292
rect 494054 389240 494060 389292
rect 494112 389280 494118 389292
rect 494606 389280 494612 389292
rect 494112 389252 494612 389280
rect 494112 389240 494118 389252
rect 494606 389240 494612 389252
rect 494664 389240 494670 389292
rect 506474 389240 506480 389292
rect 506532 389280 506538 389292
rect 507118 389280 507124 389292
rect 506532 389252 507124 389280
rect 506532 389240 506538 389252
rect 507118 389240 507124 389252
rect 507176 389240 507182 389292
rect 507854 389240 507860 389292
rect 507912 389280 507918 389292
rect 508590 389280 508596 389292
rect 507912 389252 508596 389280
rect 507912 389240 507918 389252
rect 508590 389240 508596 389252
rect 508648 389240 508654 389292
rect 453758 389104 453764 389156
rect 453816 389144 453822 389156
rect 454678 389144 454684 389156
rect 453816 389116 454684 389144
rect 453816 389104 453822 389116
rect 454678 389104 454684 389116
rect 454736 389104 454742 389156
rect 469950 388900 469956 388952
rect 470008 388940 470014 388952
rect 477310 388940 477316 388952
rect 470008 388912 477316 388940
rect 470008 388900 470014 388912
rect 477310 388900 477316 388912
rect 477368 388900 477374 388952
rect 484670 388900 484676 388952
rect 484728 388940 484734 388952
rect 502978 388940 502984 388952
rect 484728 388912 502984 388940
rect 484728 388900 484734 388912
rect 502978 388900 502984 388912
rect 503036 388900 503042 388952
rect 468478 388832 468484 388884
rect 468536 388872 468542 388884
rect 475838 388872 475844 388884
rect 468536 388844 475844 388872
rect 468536 388832 468542 388844
rect 475838 388832 475844 388844
rect 475896 388832 475902 388884
rect 500862 388832 500868 388884
rect 500920 388872 500926 388884
rect 523678 388872 523684 388884
rect 500920 388844 523684 388872
rect 500920 388832 500926 388844
rect 523678 388832 523684 388844
rect 523736 388832 523742 388884
rect 468570 388764 468576 388816
rect 468628 388804 468634 388816
rect 481726 388804 481732 388816
rect 468628 388776 481732 388804
rect 468628 388764 468634 388776
rect 481726 388764 481732 388776
rect 481784 388764 481790 388816
rect 499390 388764 499396 388816
rect 499448 388804 499454 388816
rect 522298 388804 522304 388816
rect 499448 388776 522304 388804
rect 499448 388764 499454 388776
rect 522298 388764 522304 388776
rect 522356 388764 522362 388816
rect 469858 388696 469864 388748
rect 469916 388736 469922 388748
rect 478046 388736 478052 388748
rect 469916 388708 478052 388736
rect 469916 388696 469922 388708
rect 478046 388696 478052 388708
rect 478104 388696 478110 388748
rect 502334 388696 502340 388748
rect 502392 388736 502398 388748
rect 526438 388736 526444 388748
rect 502392 388708 526444 388736
rect 502392 388696 502398 388708
rect 526438 388696 526444 388708
rect 526496 388696 526502 388748
rect 467098 388628 467104 388680
rect 467156 388668 467162 388680
rect 482462 388668 482468 388680
rect 467156 388640 482468 388668
rect 467156 388628 467162 388640
rect 482462 388628 482468 388640
rect 482520 388628 482526 388680
rect 485406 388628 485412 388680
rect 485464 388668 485470 388680
rect 524414 388668 524420 388680
rect 485464 388640 524420 388668
rect 485464 388628 485470 388640
rect 524414 388628 524420 388640
rect 524472 388628 524478 388680
rect 463050 388560 463056 388612
rect 463108 388600 463114 388612
rect 480990 388600 480996 388612
rect 463108 388572 480996 388600
rect 463108 388560 463114 388572
rect 480990 388560 480996 388572
rect 481048 388560 481054 388612
rect 486878 388560 486884 388612
rect 486936 388600 486942 388612
rect 527174 388600 527180 388612
rect 486936 388572 527180 388600
rect 486936 388560 486942 388572
rect 527174 388560 527180 388572
rect 527232 388560 527238 388612
rect 461578 388492 461584 388544
rect 461636 388532 461642 388544
rect 478782 388532 478788 388544
rect 461636 388504 478788 388532
rect 461636 388492 461642 388504
rect 478782 388492 478788 388504
rect 478840 388492 478846 388544
rect 489822 388492 489828 388544
rect 489880 388532 489886 388544
rect 530578 388532 530584 388544
rect 489880 388504 530584 388532
rect 489880 388492 489886 388504
rect 530578 388492 530584 388504
rect 530636 388492 530642 388544
rect 456702 388424 456708 388476
rect 456760 388464 456766 388476
rect 457438 388464 457444 388476
rect 456760 388436 457444 388464
rect 456760 388424 456766 388436
rect 457438 388424 457444 388436
rect 457496 388424 457502 388476
rect 461762 388424 461768 388476
rect 461820 388464 461826 388476
rect 480254 388464 480260 388476
rect 461820 388436 480260 388464
rect 461820 388424 461826 388436
rect 480254 388424 480260 388436
rect 480312 388424 480318 388476
rect 488350 388424 488356 388476
rect 488408 388464 488414 388476
rect 529198 388464 529204 388476
rect 488408 388436 529204 388464
rect 488408 388424 488414 388436
rect 529198 388424 529204 388436
rect 529256 388424 529262 388476
rect 464338 388016 464344 388068
rect 464396 388056 464402 388068
rect 469214 388056 469220 388068
rect 464396 388028 469220 388056
rect 464396 388016 464402 388028
rect 469214 388016 469220 388028
rect 469272 388016 469278 388068
rect 465718 387948 465724 388000
rect 465776 387988 465782 388000
rect 469950 387988 469956 388000
rect 465776 387960 469956 387988
rect 465776 387948 465782 387960
rect 469950 387948 469956 387960
rect 470008 387948 470014 388000
rect 459646 387812 459652 387864
rect 459704 387852 459710 387864
rect 461670 387852 461676 387864
rect 459704 387824 461676 387852
rect 459704 387812 459710 387824
rect 461670 387812 461676 387824
rect 461728 387812 461734 387864
rect 447686 387404 447692 387456
rect 447744 387444 447750 387456
rect 452010 387444 452016 387456
rect 447744 387416 452016 387444
rect 447744 387404 447750 387416
rect 452010 387404 452016 387416
rect 452068 387404 452074 387456
rect 447778 387200 447784 387252
rect 447836 387240 447842 387252
rect 462958 387240 462964 387252
rect 447836 387212 462964 387240
rect 447836 387200 447842 387212
rect 462958 387200 462964 387212
rect 463016 387200 463022 387252
rect 448974 387132 448980 387184
rect 449032 387172 449038 387184
rect 491110 387172 491116 387184
rect 449032 387144 491116 387172
rect 449032 387132 449038 387144
rect 491110 387132 491116 387144
rect 491168 387132 491174 387184
rect 449066 387064 449072 387116
rect 449124 387104 449130 387116
rect 513374 387104 513380 387116
rect 449124 387076 513380 387104
rect 449124 387064 449130 387076
rect 513374 387064 513380 387076
rect 513432 387064 513438 387116
rect 445570 386588 445576 386640
rect 445628 386628 445634 386640
rect 553946 386628 553952 386640
rect 445628 386600 553952 386628
rect 445628 386588 445634 386600
rect 553946 386588 553952 386600
rect 554004 386588 554010 386640
rect 371878 386520 371884 386572
rect 371936 386560 371942 386572
rect 512270 386560 512276 386572
rect 371936 386532 512276 386560
rect 371936 386520 371942 386532
rect 512270 386520 512276 386532
rect 512328 386520 512334 386572
rect 364978 386452 364984 386504
rect 365036 386492 365042 386504
rect 512178 386492 512184 386504
rect 365036 386464 512184 386492
rect 365036 386452 365042 386464
rect 512178 386452 512184 386464
rect 512236 386452 512242 386504
rect 360838 386384 360844 386436
rect 360896 386424 360902 386436
rect 512086 386424 512092 386436
rect 360896 386396 512092 386424
rect 360896 386384 360902 386396
rect 512086 386384 512092 386396
rect 512144 386384 512150 386436
rect 448422 385976 448428 386028
rect 448480 386016 448486 386028
rect 451918 386016 451924 386028
rect 448480 385988 451924 386016
rect 448480 385976 448486 385988
rect 451918 385976 451924 385988
rect 451976 385976 451982 386028
rect 450354 385092 450360 385144
rect 450412 385132 450418 385144
rect 563422 385132 563428 385144
rect 450412 385104 563428 385132
rect 450412 385092 450418 385104
rect 563422 385092 563428 385104
rect 563480 385092 563486 385144
rect 366358 385024 366364 385076
rect 366416 385064 366422 385076
rect 511994 385064 512000 385076
rect 366416 385036 512000 385064
rect 366416 385024 366422 385036
rect 511994 385024 512000 385036
rect 512052 385024 512058 385076
rect 365070 384956 365076 385008
rect 365128 384996 365134 385008
rect 447134 384996 447140 385008
rect 365128 384968 447140 384996
rect 365128 384956 365134 384968
rect 447134 384956 447140 384968
rect 447192 384956 447198 385008
rect 512730 383732 512736 383784
rect 512788 383772 512794 383784
rect 530578 383772 530584 383784
rect 512788 383744 530584 383772
rect 512788 383732 512794 383744
rect 530578 383732 530584 383744
rect 530636 383732 530642 383784
rect 513282 383664 513288 383716
rect 513340 383704 513346 383716
rect 547138 383704 547144 383716
rect 513340 383676 547144 383704
rect 513340 383664 513346 383676
rect 547138 383664 547144 383676
rect 547196 383664 547202 383716
rect 381538 383596 381544 383648
rect 381596 383636 381602 383648
rect 447134 383636 447140 383648
rect 381596 383608 447140 383636
rect 381596 383596 381602 383608
rect 447134 383596 447140 383608
rect 447192 383596 447198 383648
rect 406378 383528 406384 383580
rect 406436 383568 406442 383580
rect 447226 383568 447232 383580
rect 406436 383540 447232 383568
rect 406436 383528 406442 383540
rect 447226 383528 447232 383540
rect 447284 383528 447290 383580
rect 511994 383528 512000 383580
rect 512052 383568 512058 383580
rect 512546 383568 512552 383580
rect 512052 383540 512552 383568
rect 512052 383528 512058 383540
rect 512546 383528 512552 383540
rect 512604 383528 512610 383580
rect 512822 382984 512828 383036
rect 512880 383024 512886 383036
rect 518158 383024 518164 383036
rect 512880 382996 518164 383024
rect 512880 382984 512886 382996
rect 518158 382984 518164 382996
rect 518216 382984 518222 383036
rect 512454 382440 512460 382492
rect 512512 382480 512518 382492
rect 515582 382480 515588 382492
rect 512512 382452 515588 382480
rect 512512 382440 512518 382452
rect 515582 382440 515588 382452
rect 515640 382440 515646 382492
rect 513006 382372 513012 382424
rect 513064 382412 513070 382424
rect 519630 382412 519636 382424
rect 513064 382384 519636 382412
rect 513064 382372 513070 382384
rect 519630 382372 519636 382384
rect 519688 382372 519694 382424
rect 378778 382168 378784 382220
rect 378836 382208 378842 382220
rect 447134 382208 447140 382220
rect 378836 382180 447140 382208
rect 378836 382168 378842 382180
rect 447134 382168 447140 382180
rect 447192 382168 447198 382220
rect 407758 382100 407764 382152
rect 407816 382140 407822 382152
rect 447226 382140 447232 382152
rect 407816 382112 447232 382140
rect 407816 382100 407822 382112
rect 447226 382100 447232 382112
rect 447284 382100 447290 382152
rect 361574 380876 361580 380928
rect 361632 380916 361638 380928
rect 442350 380916 442356 380928
rect 361632 380888 442356 380916
rect 361632 380876 361638 380888
rect 442350 380876 442356 380888
rect 442408 380876 442414 380928
rect 513282 380876 513288 380928
rect 513340 380916 513346 380928
rect 549898 380916 549904 380928
rect 513340 380888 549904 380916
rect 513340 380876 513346 380888
rect 549898 380876 549904 380888
rect 549956 380876 549962 380928
rect 376018 380808 376024 380860
rect 376076 380848 376082 380860
rect 447134 380848 447140 380860
rect 376076 380820 447140 380848
rect 376076 380808 376082 380820
rect 447134 380808 447140 380820
rect 447192 380808 447198 380860
rect 410518 380740 410524 380792
rect 410576 380780 410582 380792
rect 447226 380780 447232 380792
rect 410576 380752 447232 380780
rect 410576 380740 410582 380752
rect 447226 380740 447232 380752
rect 447284 380740 447290 380792
rect 512086 379856 512092 379908
rect 512144 379896 512150 379908
rect 514110 379896 514116 379908
rect 512144 379868 514116 379896
rect 512144 379856 512150 379868
rect 514110 379856 514116 379868
rect 514168 379856 514174 379908
rect 513282 379516 513288 379568
rect 513340 379556 513346 379568
rect 544378 379556 544384 379568
rect 513340 379528 544384 379556
rect 513340 379516 513346 379528
rect 544378 379516 544384 379528
rect 544436 379516 544442 379568
rect 371970 379448 371976 379500
rect 372028 379488 372034 379500
rect 447226 379488 447232 379500
rect 372028 379460 447232 379488
rect 372028 379448 372034 379460
rect 447226 379448 447232 379460
rect 447284 379448 447290 379500
rect 374638 379380 374644 379432
rect 374696 379420 374702 379432
rect 447134 379420 447140 379432
rect 374696 379392 447140 379420
rect 374696 379380 374702 379392
rect 447134 379380 447140 379392
rect 447192 379380 447198 379432
rect 512178 378292 512184 378344
rect 512236 378332 512242 378344
rect 522298 378332 522304 378344
rect 512236 378304 522304 378332
rect 512236 378292 512242 378304
rect 522298 378292 522304 378304
rect 522356 378292 522362 378344
rect 513282 378224 513288 378276
rect 513340 378264 513346 378276
rect 548518 378264 548524 378276
rect 513340 378236 548524 378264
rect 513340 378224 513346 378236
rect 548518 378224 548524 378236
rect 548576 378224 548582 378276
rect 514018 378156 514024 378208
rect 514076 378196 514082 378208
rect 579798 378196 579804 378208
rect 514076 378168 579804 378196
rect 514076 378156 514082 378168
rect 579798 378156 579804 378168
rect 579856 378156 579862 378208
rect 367738 378088 367744 378140
rect 367796 378128 367802 378140
rect 447226 378128 447232 378140
rect 367796 378100 447232 378128
rect 367796 378088 367802 378100
rect 447226 378088 447232 378100
rect 447284 378088 447290 378140
rect 370498 378020 370504 378072
rect 370556 378060 370562 378072
rect 447134 378060 447140 378072
rect 370556 378032 447140 378060
rect 370556 378020 370562 378032
rect 447134 378020 447140 378032
rect 447192 378020 447198 378072
rect 512822 377408 512828 377460
rect 512880 377448 512886 377460
rect 549990 377448 549996 377460
rect 512880 377420 549996 377448
rect 512880 377408 512886 377420
rect 549990 377408 549996 377420
rect 550048 377408 550054 377460
rect 513282 376796 513288 376848
rect 513340 376836 513346 376848
rect 517514 376836 517520 376848
rect 513340 376808 517520 376836
rect 513340 376796 513346 376808
rect 517514 376796 517520 376808
rect 517572 376796 517578 376848
rect 363690 376660 363696 376712
rect 363748 376700 363754 376712
rect 447226 376700 447232 376712
rect 363748 376672 447232 376700
rect 363748 376660 363754 376672
rect 447226 376660 447232 376672
rect 447284 376660 447290 376712
rect 363598 376592 363604 376644
rect 363656 376632 363662 376644
rect 447134 376632 447140 376644
rect 363656 376604 447140 376632
rect 363656 376592 363662 376604
rect 447134 376592 447140 376604
rect 447192 376592 447198 376644
rect 512362 375980 512368 376032
rect 512420 376020 512426 376032
rect 547230 376020 547236 376032
rect 512420 375992 547236 376020
rect 512420 375980 512426 375992
rect 547230 375980 547236 375992
rect 547288 375980 547294 376032
rect 512454 375504 512460 375556
rect 512512 375544 512518 375556
rect 520274 375544 520280 375556
rect 512512 375516 520280 375544
rect 512512 375504 512518 375516
rect 520274 375504 520280 375516
rect 520332 375504 520338 375556
rect 512730 375368 512736 375420
rect 512788 375408 512794 375420
rect 516134 375408 516140 375420
rect 512788 375380 516140 375408
rect 512788 375368 512794 375380
rect 516134 375368 516140 375380
rect 516192 375368 516198 375420
rect 363782 375300 363788 375352
rect 363840 375340 363846 375352
rect 447134 375340 447140 375352
rect 363840 375312 447140 375340
rect 363840 375300 363846 375312
rect 447134 375300 447140 375312
rect 447192 375300 447198 375352
rect 411898 375232 411904 375284
rect 411956 375272 411962 375284
rect 447226 375272 447232 375284
rect 411956 375244 447232 375272
rect 411956 375232 411962 375244
rect 447226 375232 447232 375244
rect 447284 375232 447290 375284
rect 513282 374008 513288 374060
rect 513340 374048 513346 374060
rect 518894 374048 518900 374060
rect 513340 374020 518900 374048
rect 513340 374008 513346 374020
rect 518894 374008 518900 374020
rect 518952 374008 518958 374060
rect 414658 373940 414664 373992
rect 414716 373980 414722 373992
rect 447134 373980 447140 373992
rect 414716 373952 447140 373980
rect 414716 373940 414722 373952
rect 447134 373940 447140 373952
rect 447192 373940 447198 373992
rect 416314 373872 416320 373924
rect 416372 373912 416378 373924
rect 447226 373912 447232 373924
rect 416372 373884 447232 373912
rect 416372 373872 416378 373884
rect 447226 373872 447232 373884
rect 447284 373872 447290 373924
rect 512638 373328 512644 373380
rect 512696 373368 512702 373380
rect 517698 373368 517704 373380
rect 512696 373340 517704 373368
rect 512696 373328 512702 373340
rect 517698 373328 517704 373340
rect 517756 373328 517762 373380
rect 513282 372648 513288 372700
rect 513340 372688 513346 372700
rect 518986 372688 518992 372700
rect 513340 372660 518992 372688
rect 513340 372648 513346 372660
rect 518986 372648 518992 372660
rect 519044 372648 519050 372700
rect 512638 372580 512644 372632
rect 512696 372620 512702 372632
rect 523034 372620 523040 372632
rect 512696 372592 523040 372620
rect 512696 372580 512702 372592
rect 523034 372580 523040 372592
rect 523092 372580 523098 372632
rect 362218 372512 362224 372564
rect 362276 372552 362282 372564
rect 447134 372552 447140 372564
rect 362276 372524 447140 372552
rect 362276 372512 362282 372524
rect 447134 372512 447140 372524
rect 447192 372512 447198 372564
rect 418706 372444 418712 372496
rect 418764 372484 418770 372496
rect 447226 372484 447232 372496
rect 418764 372456 447232 372484
rect 418764 372444 418770 372456
rect 447226 372444 447232 372456
rect 447284 372444 447290 372496
rect 433978 371492 433984 371544
rect 434036 371532 434042 371544
rect 435358 371532 435364 371544
rect 434036 371504 435364 371532
rect 434036 371492 434042 371504
rect 435358 371492 435364 371504
rect 435416 371492 435422 371544
rect 512086 371356 512092 371408
rect 512144 371396 512150 371408
rect 514846 371396 514852 371408
rect 512144 371368 514852 371396
rect 512144 371356 512150 371368
rect 514846 371356 514852 371368
rect 514904 371356 514910 371408
rect 382918 371152 382924 371204
rect 382976 371192 382982 371204
rect 447226 371192 447232 371204
rect 382976 371164 447232 371192
rect 382976 371152 382982 371164
rect 447226 371152 447232 371164
rect 447284 371152 447290 371204
rect 417418 371084 417424 371136
rect 417476 371124 417482 371136
rect 447134 371124 447140 371136
rect 417476 371096 447140 371124
rect 417476 371084 417482 371096
rect 447134 371084 447140 371096
rect 447192 371084 447198 371136
rect 512086 370948 512092 371000
rect 512144 370988 512150 371000
rect 514754 370988 514760 371000
rect 512144 370960 514760 370988
rect 512144 370948 512150 370960
rect 514754 370948 514760 370960
rect 514812 370948 514818 371000
rect 361574 369860 361580 369912
rect 361632 369900 361638 369912
rect 429194 369900 429200 369912
rect 361632 369872 429200 369900
rect 361632 369860 361638 369872
rect 429194 369860 429200 369872
rect 429252 369860 429258 369912
rect 418614 369792 418620 369844
rect 418672 369832 418678 369844
rect 447226 369832 447232 369844
rect 418672 369804 447232 369832
rect 418672 369792 418678 369804
rect 447226 369792 447232 369804
rect 447284 369792 447290 369844
rect 436738 369724 436744 369776
rect 436796 369764 436802 369776
rect 447134 369764 447140 369776
rect 436796 369736 447140 369764
rect 436796 369724 436802 369736
rect 447134 369724 447140 369736
rect 447192 369724 447198 369776
rect 512270 368840 512276 368892
rect 512328 368880 512334 368892
rect 514938 368880 514944 368892
rect 512328 368852 514944 368880
rect 512328 368840 512334 368852
rect 514938 368840 514944 368852
rect 514996 368840 515002 368892
rect 512730 368500 512736 368552
rect 512788 368540 512794 368552
rect 516226 368540 516232 368552
rect 512788 368512 516232 368540
rect 512788 368500 512794 368512
rect 516226 368500 516232 368512
rect 516284 368500 516290 368552
rect 439498 368432 439504 368484
rect 439556 368472 439562 368484
rect 447226 368472 447232 368484
rect 439556 368444 447232 368472
rect 439556 368432 439562 368444
rect 447226 368432 447232 368444
rect 447284 368432 447290 368484
rect 440878 368364 440884 368416
rect 440936 368404 440942 368416
rect 447134 368404 447140 368416
rect 440936 368376 447140 368404
rect 440936 368364 440942 368376
rect 447134 368364 447140 368376
rect 447192 368364 447198 368416
rect 513282 367344 513288 367396
rect 513340 367384 513346 367396
rect 520366 367384 520372 367396
rect 513340 367356 520372 367384
rect 513340 367344 513346 367356
rect 520366 367344 520372 367356
rect 520424 367344 520430 367396
rect 511994 367140 512000 367192
rect 512052 367180 512058 367192
rect 514202 367180 514208 367192
rect 512052 367152 514208 367180
rect 512052 367140 512058 367152
rect 514202 367140 514208 367152
rect 514260 367140 514266 367192
rect 440970 367004 440976 367056
rect 441028 367044 441034 367056
rect 447134 367044 447140 367056
rect 441028 367016 447140 367044
rect 441028 367004 441034 367016
rect 447134 367004 447140 367016
rect 447192 367004 447198 367056
rect 442258 366936 442264 366988
rect 442316 366976 442322 366988
rect 447226 366976 447232 366988
rect 442316 366948 447232 366976
rect 442316 366936 442322 366948
rect 447226 366936 447232 366948
rect 447284 366936 447290 366988
rect 513282 365848 513288 365900
rect 513340 365888 513346 365900
rect 517790 365888 517796 365900
rect 513340 365860 517796 365888
rect 513340 365848 513346 365860
rect 517790 365848 517796 365860
rect 517848 365848 517854 365900
rect 513006 365712 513012 365764
rect 513064 365752 513070 365764
rect 516778 365752 516784 365764
rect 513064 365724 516784 365752
rect 513064 365712 513070 365724
rect 516778 365712 516784 365724
rect 516836 365712 516842 365764
rect 429194 365644 429200 365696
rect 429252 365684 429258 365696
rect 447134 365684 447140 365696
rect 429252 365656 447140 365684
rect 429252 365644 429258 365656
rect 447134 365644 447140 365656
rect 447192 365644 447198 365696
rect 442350 365576 442356 365628
rect 442408 365616 442414 365628
rect 447226 365616 447232 365628
rect 442408 365588 447232 365616
rect 442408 365576 442414 365588
rect 447226 365576 447232 365588
rect 447284 365576 447290 365628
rect 569494 364352 569500 364404
rect 569552 364392 569558 364404
rect 580166 364392 580172 364404
rect 569552 364364 580172 364392
rect 569552 364352 569558 364364
rect 580166 364352 580172 364364
rect 580224 364352 580230 364404
rect 511994 363332 512000 363384
rect 512052 363372 512058 363384
rect 513742 363372 513748 363384
rect 512052 363344 513748 363372
rect 512052 363332 512058 363344
rect 513742 363332 513748 363344
rect 513800 363332 513806 363384
rect 513282 363264 513288 363316
rect 513340 363304 513346 363316
rect 517606 363304 517612 363316
rect 513340 363276 517612 363304
rect 513340 363264 513346 363276
rect 517606 363264 517612 363276
rect 517664 363264 517670 363316
rect 436922 362992 436928 363044
rect 436980 363032 436986 363044
rect 447134 363032 447140 363044
rect 436980 363004 447140 363032
rect 436980 362992 436986 363004
rect 447134 362992 447140 363004
rect 447192 362992 447198 363044
rect 432598 362924 432604 362976
rect 432656 362964 432662 362976
rect 447226 362964 447232 362976
rect 432656 362936 447232 362964
rect 432656 362924 432662 362936
rect 447226 362924 447232 362936
rect 447284 362924 447290 362976
rect 442258 361632 442264 361684
rect 442316 361672 442322 361684
rect 447226 361672 447232 361684
rect 442316 361644 447232 361672
rect 442316 361632 442322 361644
rect 447226 361632 447232 361644
rect 447284 361632 447290 361684
rect 439682 361564 439688 361616
rect 439740 361604 439746 361616
rect 447134 361604 447140 361616
rect 439740 361576 447140 361604
rect 439740 361564 439746 361576
rect 447134 361564 447140 361576
rect 447192 361564 447198 361616
rect 511994 361224 512000 361276
rect 512052 361264 512058 361276
rect 513650 361264 513656 361276
rect 512052 361236 513656 361264
rect 512052 361224 512058 361236
rect 513650 361224 513656 361236
rect 513708 361224 513714 361276
rect 435542 360272 435548 360324
rect 435600 360312 435606 360324
rect 435600 360284 438348 360312
rect 435600 360272 435606 360284
rect 435358 360204 435364 360256
rect 435416 360244 435422 360256
rect 438118 360244 438124 360256
rect 435416 360216 438124 360244
rect 435416 360204 435422 360216
rect 438118 360204 438124 360216
rect 438176 360204 438182 360256
rect 438320 360244 438348 360284
rect 441062 360272 441068 360324
rect 441120 360312 441126 360324
rect 447134 360312 447140 360324
rect 441120 360284 447140 360312
rect 441120 360272 441126 360284
rect 447134 360272 447140 360284
rect 447192 360272 447198 360324
rect 447226 360244 447232 360256
rect 438320 360216 447232 360244
rect 447226 360204 447232 360216
rect 447284 360204 447290 360256
rect 513282 360204 513288 360256
rect 513340 360244 513346 360256
rect 520458 360244 520464 360256
rect 513340 360216 520464 360244
rect 513340 360204 513346 360216
rect 520458 360204 520464 360216
rect 520516 360204 520522 360256
rect 548518 360136 548524 360188
rect 548576 360176 548582 360188
rect 552014 360176 552020 360188
rect 548576 360148 552020 360176
rect 548576 360136 548582 360148
rect 552014 360136 552020 360148
rect 552072 360136 552078 360188
rect 549898 359116 549904 359168
rect 549956 359156 549962 359168
rect 558178 359156 558184 359168
rect 549956 359128 558184 359156
rect 549956 359116 549962 359128
rect 558178 359116 558184 359128
rect 558236 359116 558242 359168
rect 544378 359048 544384 359100
rect 544436 359088 544442 359100
rect 553762 359088 553768 359100
rect 544436 359060 553768 359088
rect 544436 359048 544442 359060
rect 553762 359048 553768 359060
rect 553820 359048 553826 359100
rect 547138 358980 547144 359032
rect 547196 359020 547202 359032
rect 565538 359020 565544 359032
rect 547196 358992 565544 359020
rect 547196 358980 547202 358992
rect 565538 358980 565544 358992
rect 565596 358980 565602 359032
rect 522298 358912 522304 358964
rect 522356 358952 522362 358964
rect 550818 358952 550824 358964
rect 522356 358924 550824 358952
rect 522356 358912 522362 358924
rect 550818 358912 550824 358924
rect 550876 358912 550882 358964
rect 442350 358844 442356 358896
rect 442408 358884 442414 358896
rect 447226 358884 447232 358896
rect 442408 358856 447232 358884
rect 442408 358844 442414 358856
rect 447226 358844 447232 358856
rect 447284 358844 447290 358896
rect 512638 358844 512644 358896
rect 512696 358884 512702 358896
rect 516410 358884 516416 358896
rect 512696 358856 516416 358884
rect 512696 358844 512702 358856
rect 516410 358844 516416 358856
rect 516468 358844 516474 358896
rect 530578 358844 530584 358896
rect 530636 358884 530642 358896
rect 567010 358884 567016 358896
rect 530636 358856 567016 358884
rect 530636 358844 530642 358856
rect 567010 358844 567016 358856
rect 567068 358844 567074 358896
rect 436830 358776 436836 358828
rect 436888 358816 436894 358828
rect 447134 358816 447140 358828
rect 436888 358788 447140 358816
rect 436888 358776 436894 358788
rect 447134 358776 447140 358788
rect 447192 358776 447198 358828
rect 514110 358776 514116 358828
rect 514168 358816 514174 358828
rect 555234 358816 555240 358828
rect 514168 358788 555240 358816
rect 514168 358776 514174 358788
rect 555234 358776 555240 358788
rect 555292 358776 555298 358828
rect 549990 358708 549996 358760
rect 550048 358748 550054 358760
rect 556706 358748 556712 358760
rect 550048 358720 556712 358748
rect 550048 358708 550054 358720
rect 556706 358708 556712 358720
rect 556764 358708 556770 358760
rect 518158 358640 518164 358692
rect 518216 358680 518222 358692
rect 562594 358680 562600 358692
rect 518216 358652 562600 358680
rect 518216 358640 518222 358652
rect 562594 358640 562600 358652
rect 562652 358640 562658 358692
rect 519630 358572 519636 358624
rect 519688 358612 519694 358624
rect 564066 358612 564072 358624
rect 519688 358584 564072 358612
rect 519688 358572 519694 358584
rect 564066 358572 564072 358584
rect 564124 358572 564130 358624
rect 547230 358504 547236 358556
rect 547288 358544 547294 358556
rect 559650 358544 559656 358556
rect 547288 358516 559656 358544
rect 547288 358504 547294 358516
rect 559650 358504 559656 358516
rect 559708 358504 559714 358556
rect 515582 358436 515588 358488
rect 515640 358476 515646 358488
rect 561122 358476 561128 358488
rect 515640 358448 561128 358476
rect 515640 358436 515646 358448
rect 561122 358436 561128 358448
rect 561180 358436 561186 358488
rect 513190 357688 513196 357740
rect 513248 357728 513254 357740
rect 517882 357728 517888 357740
rect 513248 357700 517888 357728
rect 513248 357688 513254 357700
rect 517882 357688 517888 357700
rect 517940 357688 517946 357740
rect 513282 356328 513288 356380
rect 513340 356368 513346 356380
rect 519078 356368 519084 356380
rect 513340 356340 519084 356368
rect 513340 356328 513346 356340
rect 519078 356328 519084 356340
rect 519136 356328 519142 356380
rect 512270 355376 512276 355428
rect 512328 355416 512334 355428
rect 515122 355416 515128 355428
rect 512328 355388 515128 355416
rect 512328 355376 512334 355388
rect 515122 355376 515128 355388
rect 515180 355376 515186 355428
rect 513282 354968 513288 355020
rect 513340 355008 513346 355020
rect 520550 355008 520556 355020
rect 513340 354980 520556 355008
rect 513340 354968 513346 354980
rect 520550 354968 520556 354980
rect 520608 354968 520614 355020
rect 513282 354696 513288 354748
rect 513340 354736 513346 354748
rect 517974 354736 517980 354748
rect 513340 354708 517980 354736
rect 513340 354696 513346 354708
rect 517974 354696 517980 354708
rect 518032 354696 518038 354748
rect 512822 353472 512828 353524
rect 512880 353512 512886 353524
rect 516318 353512 516324 353524
rect 512880 353484 516324 353512
rect 512880 353472 512886 353484
rect 516318 353472 516324 353484
rect 516376 353472 516382 353524
rect 512454 353336 512460 353388
rect 512512 353376 512518 353388
rect 515214 353376 515220 353388
rect 512512 353348 515220 353376
rect 512512 353336 512518 353348
rect 515214 353336 515220 353348
rect 515272 353336 515278 353388
rect 513006 352656 513012 352708
rect 513064 352696 513070 352708
rect 516594 352696 516600 352708
rect 513064 352668 516600 352696
rect 513064 352656 513070 352668
rect 516594 352656 516600 352668
rect 516652 352656 516658 352708
rect 512454 351976 512460 352028
rect 512512 352016 512518 352028
rect 515030 352016 515036 352028
rect 512512 351988 515036 352016
rect 512512 351976 512518 351988
rect 515030 351976 515036 351988
rect 515088 351976 515094 352028
rect 394694 351908 394700 351960
rect 394752 351948 394758 351960
rect 447134 351948 447140 351960
rect 394752 351920 447140 351948
rect 394752 351908 394758 351920
rect 447134 351908 447140 351920
rect 447192 351908 447198 351960
rect 513282 350888 513288 350940
rect 513340 350928 513346 350940
rect 518066 350928 518072 350940
rect 513340 350900 518072 350928
rect 513340 350888 513346 350900
rect 518066 350888 518072 350900
rect 518124 350888 518130 350940
rect 512454 350752 512460 350804
rect 512512 350792 512518 350804
rect 513926 350792 513932 350804
rect 512512 350764 513932 350792
rect 512512 350752 512518 350764
rect 513926 350752 513932 350764
rect 513984 350752 513990 350804
rect 405734 350548 405740 350600
rect 405792 350588 405798 350600
rect 447134 350588 447140 350600
rect 405792 350560 447140 350588
rect 405792 350548 405798 350560
rect 447134 350548 447140 350560
rect 447192 350548 447198 350600
rect 512822 349800 512828 349852
rect 512880 349840 512886 349852
rect 516502 349840 516508 349852
rect 512880 349812 516508 349840
rect 512880 349800 512886 349812
rect 516502 349800 516508 349812
rect 516560 349800 516566 349852
rect 512454 349256 512460 349308
rect 512512 349296 512518 349308
rect 513834 349296 513840 349308
rect 512512 349268 513840 349296
rect 512512 349256 512518 349268
rect 513834 349256 513840 349268
rect 513892 349256 513898 349308
rect 512546 349188 512552 349240
rect 512604 349228 512610 349240
rect 515306 349228 515312 349240
rect 512604 349200 515312 349228
rect 512604 349188 512610 349200
rect 515306 349188 515312 349200
rect 515364 349188 515370 349240
rect 446950 349052 446956 349104
rect 447008 349092 447014 349104
rect 447778 349092 447784 349104
rect 447008 349064 447784 349092
rect 447008 349052 447014 349064
rect 447778 349052 447784 349064
rect 447836 349052 447842 349104
rect 412634 348372 412640 348424
rect 412692 348412 412698 348424
rect 435634 348412 435640 348424
rect 412692 348384 435640 348412
rect 412692 348372 412698 348384
rect 435634 348372 435640 348384
rect 435692 348372 435698 348424
rect 513282 347896 513288 347948
rect 513340 347936 513346 347948
rect 519170 347936 519176 347948
rect 513340 347908 519176 347936
rect 513340 347896 513346 347908
rect 519170 347896 519176 347908
rect 519228 347896 519234 347948
rect 361758 347760 361764 347812
rect 361816 347800 361822 347812
rect 389818 347800 389824 347812
rect 361816 347772 389824 347800
rect 361816 347760 361822 347772
rect 389818 347760 389824 347772
rect 389876 347760 389882 347812
rect 513098 347760 513104 347812
rect 513156 347800 513162 347812
rect 516686 347800 516692 347812
rect 513156 347772 516692 347800
rect 513156 347760 513162 347772
rect 516686 347760 516692 347772
rect 516744 347760 516750 347812
rect 362310 347692 362316 347744
rect 362368 347732 362374 347744
rect 447134 347732 447140 347744
rect 362368 347704 447140 347732
rect 362368 347692 362374 347704
rect 447134 347692 447140 347704
rect 447192 347692 447198 347744
rect 513282 345176 513288 345228
rect 513340 345216 513346 345228
rect 520642 345216 520648 345228
rect 513340 345188 520648 345216
rect 513340 345176 513346 345188
rect 520642 345176 520648 345188
rect 520700 345176 520706 345228
rect 432690 344292 432696 344344
rect 432748 344332 432754 344344
rect 442258 344332 442264 344344
rect 432748 344304 442264 344332
rect 432748 344292 432754 344304
rect 442258 344292 442264 344304
rect 442316 344292 442322 344344
rect 513282 344224 513288 344276
rect 513340 344264 513346 344276
rect 518158 344264 518164 344276
rect 513340 344236 518164 344264
rect 513340 344224 513346 344236
rect 518158 344224 518164 344236
rect 518216 344224 518222 344276
rect 513282 343816 513288 343868
rect 513340 343856 513346 343868
rect 520734 343856 520740 343868
rect 513340 343828 520740 343856
rect 513340 343816 513346 343828
rect 520734 343816 520740 343828
rect 520792 343816 520798 343868
rect 445570 343068 445576 343120
rect 445628 343108 445634 343120
rect 449710 343108 449716 343120
rect 445628 343080 449716 343108
rect 445628 343068 445634 343080
rect 449710 343068 449716 343080
rect 449768 343068 449774 343120
rect 401594 342864 401600 342916
rect 401652 342904 401658 342916
rect 445570 342904 445576 342916
rect 401652 342876 445576 342904
rect 401652 342864 401658 342876
rect 445570 342864 445576 342876
rect 445628 342864 445634 342916
rect 512454 342524 512460 342576
rect 512512 342564 512518 342576
rect 515582 342564 515588 342576
rect 512512 342536 515588 342564
rect 512512 342524 512518 342536
rect 515582 342524 515588 342536
rect 515640 342524 515646 342576
rect 513282 342252 513288 342304
rect 513340 342292 513346 342304
rect 521654 342292 521660 342304
rect 513340 342264 521660 342292
rect 513340 342252 513346 342264
rect 521654 342252 521660 342264
rect 521712 342252 521718 342304
rect 513282 341232 513288 341284
rect 513340 341272 513346 341284
rect 519262 341272 519268 341284
rect 513340 341244 519268 341272
rect 513340 341232 513346 341244
rect 519262 341232 519268 341244
rect 519320 341232 519326 341284
rect 513098 341096 513104 341148
rect 513156 341136 513162 341148
rect 516870 341136 516876 341148
rect 513156 341108 516876 341136
rect 513156 341096 513162 341108
rect 516870 341096 516876 341108
rect 516928 341096 516934 341148
rect 442902 340960 442908 341012
rect 442960 341000 442966 341012
rect 447226 341000 447232 341012
rect 442960 340972 447232 341000
rect 442960 340960 442966 340972
rect 447226 340960 447232 340972
rect 447284 340960 447290 341012
rect 361758 340892 361764 340944
rect 361816 340932 361822 340944
rect 447134 340932 447140 340944
rect 361816 340904 447140 340932
rect 361816 340892 361822 340904
rect 447134 340892 447140 340904
rect 447192 340892 447198 340944
rect 513282 339600 513288 339652
rect 513340 339640 513346 339652
rect 520826 339640 520832 339652
rect 513340 339612 520832 339640
rect 513340 339600 513346 339612
rect 520826 339600 520832 339612
rect 520884 339600 520890 339652
rect 443730 339532 443736 339584
rect 443788 339572 443794 339584
rect 447226 339572 447232 339584
rect 443788 339544 447232 339572
rect 443788 339532 443794 339544
rect 447226 339532 447232 339544
rect 447284 339532 447290 339584
rect 399478 339464 399484 339516
rect 399536 339504 399542 339516
rect 447134 339504 447140 339516
rect 399536 339476 447140 339504
rect 399536 339464 399542 339476
rect 447134 339464 447140 339476
rect 447192 339464 447198 339516
rect 513282 339464 513288 339516
rect 513340 339504 513346 339516
rect 518250 339504 518256 339516
rect 513340 339476 518256 339504
rect 513340 339464 513346 339476
rect 518250 339464 518256 339476
rect 518308 339464 518314 339516
rect 513282 338240 513288 338292
rect 513340 338280 513346 338292
rect 519722 338280 519728 338292
rect 513340 338252 519728 338280
rect 513340 338240 513346 338252
rect 519722 338240 519728 338252
rect 519780 338240 519786 338292
rect 431218 338172 431224 338224
rect 431276 338212 431282 338224
rect 447134 338212 447140 338224
rect 431276 338184 447140 338212
rect 431276 338172 431282 338184
rect 447134 338172 447140 338184
rect 447192 338172 447198 338224
rect 385954 338104 385960 338156
rect 386012 338144 386018 338156
rect 447226 338144 447232 338156
rect 386012 338116 447232 338144
rect 386012 338104 386018 338116
rect 447226 338104 447232 338116
rect 447284 338104 447290 338156
rect 513006 338104 513012 338156
rect 513064 338144 513070 338156
rect 521746 338144 521752 338156
rect 513064 338116 521752 338144
rect 513064 338104 513070 338116
rect 521746 338104 521752 338116
rect 521804 338104 521810 338156
rect 513006 337152 513012 337204
rect 513064 337192 513070 337204
rect 516962 337192 516968 337204
rect 513064 337164 516968 337192
rect 513064 337152 513070 337164
rect 516962 337152 516968 337164
rect 517020 337152 517026 337204
rect 416774 336880 416780 336932
rect 416832 336920 416838 336932
rect 429930 336920 429936 336932
rect 416832 336892 429936 336920
rect 416832 336880 416838 336892
rect 429930 336880 429936 336892
rect 429988 336880 429994 336932
rect 513282 336880 513288 336932
rect 513340 336920 513346 336932
rect 520918 336920 520924 336932
rect 513340 336892 520924 336920
rect 513340 336880 513346 336892
rect 520918 336880 520924 336892
rect 520976 336880 520982 336932
rect 424134 336812 424140 336864
rect 424192 336852 424198 336864
rect 431402 336852 431408 336864
rect 424192 336824 431408 336852
rect 424192 336812 424198 336824
rect 431402 336812 431408 336824
rect 431460 336812 431466 336864
rect 440970 336812 440976 336864
rect 441028 336852 441034 336864
rect 447134 336852 447140 336864
rect 441028 336824 447140 336852
rect 441028 336812 441034 336824
rect 447134 336812 447140 336824
rect 447192 336812 447198 336864
rect 420454 336744 420460 336796
rect 420512 336784 420518 336796
rect 435726 336784 435732 336796
rect 420512 336756 435732 336784
rect 420512 336744 420518 336756
rect 435726 336744 435732 336756
rect 435784 336744 435790 336796
rect 439590 336744 439596 336796
rect 439648 336784 439654 336796
rect 447226 336784 447232 336796
rect 439648 336756 447232 336784
rect 439648 336744 439654 336756
rect 447226 336744 447232 336756
rect 447284 336744 447290 336796
rect 513098 336744 513104 336796
rect 513156 336784 513162 336796
rect 523126 336784 523132 336796
rect 513156 336756 523132 336784
rect 513156 336744 513162 336756
rect 523126 336744 523132 336756
rect 523184 336744 523190 336796
rect 416222 336336 416228 336388
rect 416280 336376 416286 336388
rect 438210 336376 438216 336388
rect 416280 336348 438216 336376
rect 416280 336336 416286 336348
rect 438210 336336 438216 336348
rect 438268 336336 438274 336388
rect 419442 336268 419448 336320
rect 419500 336308 419506 336320
rect 443822 336308 443828 336320
rect 419500 336280 443828 336308
rect 419500 336268 419506 336280
rect 443822 336268 443828 336280
rect 443880 336268 443886 336320
rect 416038 336200 416044 336252
rect 416096 336240 416102 336252
rect 441154 336240 441160 336252
rect 416096 336212 441160 336240
rect 416096 336200 416102 336212
rect 441154 336200 441160 336212
rect 441212 336200 441218 336252
rect 419350 336132 419356 336184
rect 419408 336172 419414 336184
rect 446950 336172 446956 336184
rect 419408 336144 446956 336172
rect 419408 336132 419414 336144
rect 446950 336132 446956 336144
rect 447008 336132 447014 336184
rect 397454 336064 397460 336116
rect 397512 336104 397518 336116
rect 449066 336104 449072 336116
rect 397512 336076 449072 336104
rect 397512 336064 397518 336076
rect 449066 336064 449072 336076
rect 449124 336064 449130 336116
rect 513282 336064 513288 336116
rect 513340 336104 513346 336116
rect 518342 336104 518348 336116
rect 513340 336076 518348 336104
rect 513340 336064 513346 336076
rect 518342 336064 518348 336076
rect 518400 336064 518406 336116
rect 362218 335996 362224 336048
rect 362276 336036 362282 336048
rect 442902 336036 442908 336048
rect 362276 336008 442908 336036
rect 362276 335996 362282 336008
rect 442902 335996 442908 336008
rect 442960 335996 442966 336048
rect 442258 335452 442264 335504
rect 442316 335492 442322 335504
rect 447318 335492 447324 335504
rect 442316 335464 447324 335492
rect 442316 335452 442322 335464
rect 447318 335452 447324 335464
rect 447376 335452 447382 335504
rect 409414 335384 409420 335436
rect 409472 335424 409478 335436
rect 431310 335424 431316 335436
rect 409472 335396 431316 335424
rect 409472 335384 409478 335396
rect 431310 335384 431316 335396
rect 431368 335384 431374 335436
rect 435450 335384 435456 335436
rect 435508 335424 435514 335436
rect 447226 335424 447232 335436
rect 435508 335396 447232 335424
rect 435508 335384 435514 335396
rect 447226 335384 447232 335396
rect 447284 335384 447290 335436
rect 413094 335316 413100 335368
rect 413152 335356 413158 335368
rect 439774 335356 439780 335368
rect 413152 335328 439780 335356
rect 413152 335316 413158 335328
rect 439774 335316 439780 335328
rect 439832 335316 439838 335368
rect 513282 335316 513288 335368
rect 513340 335356 513346 335368
rect 521838 335356 521844 335368
rect 513340 335328 521844 335356
rect 513340 335316 513346 335328
rect 521838 335316 521844 335328
rect 521896 335316 521902 335368
rect 420178 335044 420184 335096
rect 420236 335084 420242 335096
rect 442534 335084 442540 335096
rect 420236 335056 442540 335084
rect 420236 335044 420242 335056
rect 442534 335044 442540 335056
rect 442592 335044 442598 335096
rect 418798 334976 418804 335028
rect 418856 335016 418862 335028
rect 443914 335016 443920 335028
rect 418856 334988 443920 335016
rect 418856 334976 418862 334988
rect 443914 334976 443920 334988
rect 443972 334976 443978 335028
rect 416130 334908 416136 334960
rect 416188 334948 416194 334960
rect 444006 334948 444012 334960
rect 416188 334920 444012 334948
rect 416188 334908 416194 334920
rect 444006 334908 444012 334920
rect 444064 334908 444070 334960
rect 418890 334840 418896 334892
rect 418948 334880 418954 334892
rect 447042 334880 447048 334892
rect 418948 334852 447048 334880
rect 418948 334840 418954 334852
rect 447042 334840 447048 334852
rect 447100 334840 447106 334892
rect 419258 334772 419264 334824
rect 419316 334812 419322 334824
rect 448974 334812 448980 334824
rect 419316 334784 448980 334812
rect 419316 334772 419322 334784
rect 448974 334772 448980 334784
rect 449032 334772 449038 334824
rect 419074 334704 419080 334756
rect 419132 334744 419138 334756
rect 449526 334744 449532 334756
rect 419132 334716 449532 334744
rect 419132 334704 419138 334716
rect 449526 334704 449532 334716
rect 449584 334704 449590 334756
rect 418982 334636 418988 334688
rect 419040 334676 419046 334688
rect 449434 334676 449440 334688
rect 419040 334648 449440 334676
rect 419040 334636 419046 334648
rect 449434 334636 449440 334648
rect 449492 334636 449498 334688
rect 419166 334568 419172 334620
rect 419224 334608 419230 334620
rect 450722 334608 450728 334620
rect 419224 334580 450728 334608
rect 419224 334568 419230 334580
rect 450722 334568 450728 334580
rect 450780 334568 450786 334620
rect 512454 334500 512460 334552
rect 512512 334540 512518 334552
rect 514110 334540 514116 334552
rect 512512 334512 514116 334540
rect 512512 334500 512518 334512
rect 514110 334500 514116 334512
rect 514168 334500 514174 334552
rect 428090 334364 428096 334416
rect 428148 334404 428154 334416
rect 428148 334376 431954 334404
rect 428148 334364 428154 334376
rect 431926 334132 431954 334376
rect 438118 334228 438124 334280
rect 438176 334268 438182 334280
rect 440234 334268 440240 334280
rect 438176 334240 440240 334268
rect 438176 334228 438182 334240
rect 440234 334228 440240 334240
rect 440292 334228 440298 334280
rect 512822 334160 512828 334212
rect 512880 334200 512886 334212
rect 519446 334200 519452 334212
rect 512880 334172 519452 334200
rect 512880 334160 512886 334172
rect 519446 334160 519452 334172
rect 519504 334160 519510 334212
rect 448238 334132 448244 334144
rect 431926 334104 448244 334132
rect 448238 334092 448244 334104
rect 448296 334092 448302 334144
rect 443638 334024 443644 334076
rect 443696 334064 443702 334076
rect 447318 334064 447324 334076
rect 443696 334036 447324 334064
rect 443696 334024 443702 334036
rect 447318 334024 447324 334036
rect 447376 334024 447382 334076
rect 364058 333956 364064 334008
rect 364116 333996 364122 334008
rect 447226 333996 447232 334008
rect 364116 333968 447232 333996
rect 364116 333956 364122 333968
rect 447226 333956 447232 333968
rect 447284 333956 447290 334008
rect 509234 333956 509240 334008
rect 509292 333996 509298 334008
rect 509694 333996 509700 334008
rect 509292 333968 509700 333996
rect 509292 333956 509298 333968
rect 509694 333956 509700 333968
rect 509752 333956 509758 334008
rect 511350 333208 511356 333260
rect 511408 333248 511414 333260
rect 580258 333248 580264 333260
rect 511408 333220 580264 333248
rect 511408 333208 511414 333220
rect 580258 333208 580264 333220
rect 580316 333208 580322 333260
rect 439498 332664 439504 332716
rect 439556 332704 439562 332716
rect 447318 332704 447324 332716
rect 439556 332676 447324 332704
rect 439556 332664 439562 332676
rect 447318 332664 447324 332676
rect 447376 332664 447382 332716
rect 513282 332664 513288 332716
rect 513340 332704 513346 332716
rect 519630 332704 519636 332716
rect 513340 332676 519636 332704
rect 513340 332664 513346 332676
rect 519630 332664 519636 332676
rect 519688 332664 519694 332716
rect 429838 332596 429844 332648
rect 429896 332636 429902 332648
rect 447226 332636 447232 332648
rect 429896 332608 447232 332636
rect 429896 332596 429902 332608
rect 447226 332596 447232 332608
rect 447284 332596 447290 332648
rect 440234 332528 440240 332580
rect 440292 332568 440298 332580
rect 442626 332568 442632 332580
rect 440292 332540 442632 332568
rect 440292 332528 440298 332540
rect 442626 332528 442632 332540
rect 442684 332528 442690 332580
rect 512822 331440 512828 331492
rect 512880 331480 512886 331492
rect 519354 331480 519360 331492
rect 512880 331452 519360 331480
rect 512880 331440 512886 331452
rect 519354 331440 519360 331452
rect 519412 331440 519418 331492
rect 432874 331304 432880 331356
rect 432932 331344 432938 331356
rect 439682 331344 439688 331356
rect 432932 331316 439688 331344
rect 432932 331304 432938 331316
rect 439682 331304 439688 331316
rect 439740 331304 439746 331356
rect 440878 331304 440884 331356
rect 440936 331344 440942 331356
rect 447226 331344 447232 331356
rect 440936 331316 447232 331344
rect 440936 331304 440942 331316
rect 447226 331304 447232 331316
rect 447284 331304 447290 331356
rect 436738 331236 436744 331288
rect 436796 331276 436802 331288
rect 447594 331276 447600 331288
rect 436796 331248 447600 331276
rect 436796 331236 436802 331248
rect 447594 331236 447600 331248
rect 447652 331236 447658 331288
rect 444190 330556 444196 330608
rect 444248 330596 444254 330608
rect 445754 330596 445760 330608
rect 444248 330568 445760 330596
rect 444248 330556 444254 330568
rect 445754 330556 445760 330568
rect 445812 330596 445818 330608
rect 447226 330596 447232 330608
rect 445812 330568 447232 330596
rect 445812 330556 445818 330568
rect 447226 330556 447232 330568
rect 447284 330556 447290 330608
rect 432598 330488 432604 330540
rect 432656 330528 432662 330540
rect 442350 330528 442356 330540
rect 432656 330500 442356 330528
rect 432656 330488 432662 330500
rect 442350 330488 442356 330500
rect 442408 330488 442414 330540
rect 442902 330080 442908 330132
rect 442960 330120 442966 330132
rect 445846 330120 445852 330132
rect 442960 330092 445852 330120
rect 442960 330080 442966 330092
rect 445846 330080 445852 330092
rect 445904 330120 445910 330132
rect 447226 330120 447232 330132
rect 445904 330092 447232 330120
rect 445904 330080 445910 330092
rect 447226 330080 447232 330092
rect 447284 330080 447290 330132
rect 438762 329740 438768 329792
rect 438820 329780 438826 329792
rect 444098 329780 444104 329792
rect 438820 329752 444104 329780
rect 438820 329740 438826 329752
rect 444098 329740 444104 329752
rect 444156 329780 444162 329792
rect 447226 329780 447232 329792
rect 444156 329752 447232 329780
rect 444156 329740 444162 329752
rect 447226 329740 447232 329752
rect 447284 329740 447290 329792
rect 432414 329672 432420 329724
rect 432472 329712 432478 329724
rect 436922 329712 436928 329724
rect 432472 329684 436928 329712
rect 432472 329672 432478 329684
rect 436922 329672 436928 329684
rect 436980 329672 436986 329724
rect 435358 329060 435364 329112
rect 435416 329100 435422 329112
rect 447226 329100 447232 329112
rect 435416 329072 447232 329100
rect 435416 329060 435422 329072
rect 447226 329060 447232 329072
rect 447284 329060 447290 329112
rect 432782 328856 432788 328908
rect 432840 328896 432846 328908
rect 435542 328896 435548 328908
rect 432840 328868 435548 328896
rect 432840 328856 432846 328868
rect 435542 328856 435548 328868
rect 435600 328856 435606 328908
rect 431862 327700 431868 327752
rect 431920 327740 431926 327752
rect 447226 327740 447232 327752
rect 431920 327712 447232 327740
rect 431920 327700 431926 327712
rect 447226 327700 447232 327712
rect 447284 327700 447290 327752
rect 435726 327020 435732 327072
rect 435784 327060 435790 327072
rect 447226 327060 447232 327072
rect 435784 327032 447232 327060
rect 435784 327020 435790 327032
rect 447226 327020 447232 327032
rect 447284 327060 447290 327072
rect 447870 327060 447876 327072
rect 447284 327032 447876 327060
rect 447284 327020 447290 327032
rect 447870 327020 447876 327032
rect 447928 327020 447934 327072
rect 431402 326340 431408 326392
rect 431460 326380 431466 326392
rect 441614 326380 441620 326392
rect 431460 326352 441620 326380
rect 431460 326340 431466 326352
rect 441614 326340 441620 326352
rect 441672 326380 441678 326392
rect 448146 326380 448152 326392
rect 441672 326352 448152 326380
rect 441672 326340 441678 326352
rect 448146 326340 448152 326352
rect 448204 326340 448210 326392
rect 429930 325592 429936 325644
rect 429988 325632 429994 325644
rect 447778 325632 447784 325644
rect 429988 325604 447784 325632
rect 429988 325592 429994 325604
rect 447778 325592 447784 325604
rect 447836 325632 447842 325644
rect 448054 325632 448060 325644
rect 447836 325604 448060 325632
rect 447836 325592 447842 325604
rect 448054 325592 448060 325604
rect 448112 325592 448118 325644
rect 439774 325524 439780 325576
rect 439832 325564 439838 325576
rect 447962 325564 447968 325576
rect 439832 325536 447968 325564
rect 439832 325524 439838 325536
rect 447962 325524 447968 325536
rect 448020 325524 448026 325576
rect 431310 323552 431316 323604
rect 431368 323592 431374 323604
rect 447318 323592 447324 323604
rect 431368 323564 447324 323592
rect 431368 323552 431374 323564
rect 447318 323552 447324 323564
rect 447376 323552 447382 323604
rect 512914 322940 512920 322992
rect 512972 322980 512978 322992
rect 519538 322980 519544 322992
rect 512972 322952 519544 322980
rect 512972 322940 512978 322952
rect 519538 322940 519544 322952
rect 519596 322940 519602 322992
rect 442626 322872 442632 322924
rect 442684 322912 442690 322924
rect 449894 322912 449900 322924
rect 442684 322884 449900 322912
rect 442684 322872 442690 322884
rect 449894 322872 449900 322884
rect 449952 322872 449958 322924
rect 514018 322464 514024 322516
rect 514076 322504 514082 322516
rect 514294 322504 514300 322516
rect 514076 322476 514300 322504
rect 514076 322464 514082 322476
rect 514294 322464 514300 322476
rect 514352 322464 514358 322516
rect 510522 322396 510528 322448
rect 510580 322436 510586 322448
rect 580626 322436 580632 322448
rect 510580 322408 580632 322436
rect 510580 322396 510586 322408
rect 580626 322396 580632 322408
rect 580684 322396 580690 322448
rect 510062 322328 510068 322380
rect 510120 322368 510126 322380
rect 580534 322368 580540 322380
rect 510120 322340 580540 322368
rect 510120 322328 510126 322340
rect 580534 322328 580540 322340
rect 580592 322328 580598 322380
rect 514018 322260 514024 322312
rect 514076 322300 514082 322312
rect 580350 322300 580356 322312
rect 514076 322272 580356 322300
rect 514076 322260 514082 322272
rect 580350 322260 580356 322272
rect 580408 322260 580414 322312
rect 509142 322192 509148 322244
rect 509200 322232 509206 322244
rect 580166 322232 580172 322244
rect 509200 322204 580172 322232
rect 509200 322192 509206 322204
rect 580166 322192 580172 322204
rect 580224 322192 580230 322244
rect 507210 321852 507216 321904
rect 507268 321892 507274 321904
rect 509234 321892 509240 321904
rect 507268 321864 509240 321892
rect 507268 321852 507274 321864
rect 509234 321852 509240 321864
rect 509292 321852 509298 321904
rect 444006 321784 444012 321836
rect 444064 321824 444070 321836
rect 462130 321824 462136 321836
rect 444064 321796 462136 321824
rect 444064 321784 444070 321796
rect 462130 321784 462136 321796
rect 462188 321784 462194 321836
rect 507578 321784 507584 321836
rect 507636 321824 507642 321836
rect 509878 321824 509884 321836
rect 507636 321796 509884 321824
rect 507636 321784 507642 321796
rect 509878 321784 509884 321796
rect 509936 321784 509942 321836
rect 450722 321716 450728 321768
rect 450780 321756 450786 321768
rect 482554 321756 482560 321768
rect 450780 321728 482560 321756
rect 450780 321716 450786 321728
rect 482554 321716 482560 321728
rect 482612 321716 482618 321768
rect 507946 321716 507952 321768
rect 508004 321756 508010 321768
rect 510062 321756 510068 321768
rect 508004 321728 510068 321756
rect 508004 321716 508010 321728
rect 510062 321716 510068 321728
rect 510120 321716 510126 321768
rect 448974 321648 448980 321700
rect 449032 321688 449038 321700
rect 472342 321688 472348 321700
rect 449032 321660 472348 321688
rect 449032 321648 449038 321660
rect 472342 321648 472348 321660
rect 472400 321648 472406 321700
rect 507854 321648 507860 321700
rect 507912 321688 507918 321700
rect 514018 321688 514024 321700
rect 507912 321660 514024 321688
rect 507912 321648 507918 321660
rect 514018 321648 514024 321660
rect 514076 321648 514082 321700
rect 442534 321580 442540 321632
rect 442592 321620 442598 321632
rect 482278 321620 482284 321632
rect 442592 321592 482284 321620
rect 442592 321580 442598 321592
rect 482278 321580 482284 321592
rect 482336 321580 482342 321632
rect 456610 321512 456616 321564
rect 456668 321552 456674 321564
rect 580902 321552 580908 321564
rect 456668 321524 580908 321552
rect 456668 321512 456674 321524
rect 580902 321512 580908 321524
rect 580960 321512 580966 321564
rect 456334 321444 456340 321496
rect 456392 321484 456398 321496
rect 580074 321484 580080 321496
rect 456392 321456 580080 321484
rect 456392 321444 456398 321456
rect 580074 321444 580080 321456
rect 580132 321444 580138 321496
rect 457990 321376 457996 321428
rect 458048 321416 458054 321428
rect 580442 321416 580448 321428
rect 458048 321388 580448 321416
rect 458048 321376 458054 321388
rect 580442 321376 580448 321388
rect 580500 321376 580506 321428
rect 449158 321308 449164 321360
rect 449216 321348 449222 321360
rect 459370 321348 459376 321360
rect 449216 321320 459376 321348
rect 449216 321308 449222 321320
rect 459370 321308 459376 321320
rect 459428 321308 459434 321360
rect 466822 321308 466828 321360
rect 466880 321348 466886 321360
rect 569494 321348 569500 321360
rect 466880 321320 569500 321348
rect 466880 321308 466886 321320
rect 569494 321308 569500 321320
rect 569552 321308 569558 321360
rect 445018 321240 445024 321292
rect 445076 321280 445082 321292
rect 459094 321280 459100 321292
rect 445076 321252 459100 321280
rect 445076 321240 445082 321252
rect 459094 321240 459100 321252
rect 459152 321240 459158 321292
rect 468202 321240 468208 321292
rect 468260 321280 468266 321292
rect 567838 321280 567844 321292
rect 468260 321252 567844 321280
rect 468260 321240 468266 321252
rect 567838 321240 567844 321252
rect 567896 321240 567902 321292
rect 445110 321172 445116 321224
rect 445168 321212 445174 321224
rect 458818 321212 458824 321224
rect 445168 321184 458824 321212
rect 445168 321172 445174 321184
rect 458818 321172 458824 321184
rect 458876 321172 458882 321224
rect 477586 321172 477592 321224
rect 477644 321212 477650 321224
rect 569402 321212 569408 321224
rect 477644 321184 569408 321212
rect 477644 321172 477650 321184
rect 569402 321172 569408 321184
rect 569460 321172 569466 321224
rect 449250 321104 449256 321156
rect 449308 321144 449314 321156
rect 460474 321144 460480 321156
rect 449308 321116 460480 321144
rect 449308 321104 449314 321116
rect 460474 321104 460480 321116
rect 460532 321104 460538 321156
rect 467650 321104 467656 321156
rect 467708 321144 467714 321156
rect 515398 321144 515404 321156
rect 467708 321116 515404 321144
rect 467708 321104 467714 321116
rect 515398 321104 515404 321116
rect 515456 321104 515462 321156
rect 445202 321036 445208 321088
rect 445260 321076 445266 321088
rect 460198 321076 460204 321088
rect 445260 321048 460204 321076
rect 445260 321036 445266 321048
rect 460198 321036 460204 321048
rect 460256 321036 460262 321088
rect 467374 321036 467380 321088
rect 467432 321076 467438 321088
rect 511258 321076 511264 321088
rect 467432 321048 511264 321076
rect 467432 321036 467438 321048
rect 511258 321036 511264 321048
rect 511316 321036 511322 321088
rect 449066 320968 449072 321020
rect 449124 321008 449130 321020
rect 479794 321008 479800 321020
rect 449124 320980 479800 321008
rect 449124 320968 449130 320980
rect 479794 320968 479800 320980
rect 479852 320968 479858 321020
rect 445662 320900 445668 320952
rect 445720 320940 445726 320952
rect 469030 320940 469036 320952
rect 445720 320912 469036 320940
rect 445720 320900 445726 320912
rect 469030 320900 469036 320912
rect 469088 320900 469094 320952
rect 507394 320900 507400 320952
rect 507452 320940 507458 320952
rect 513374 320940 513380 320952
rect 507452 320912 513380 320940
rect 507452 320900 507458 320912
rect 513374 320900 513380 320912
rect 513432 320900 513438 320952
rect 449894 320832 449900 320884
rect 449952 320872 449958 320884
rect 469214 320872 469220 320884
rect 449952 320844 469220 320872
rect 449952 320832 449958 320844
rect 469214 320832 469220 320844
rect 469272 320832 469278 320884
rect 506934 320832 506940 320884
rect 506992 320872 506998 320884
rect 516778 320872 516784 320884
rect 506992 320844 516784 320872
rect 506992 320832 506998 320844
rect 516778 320832 516784 320844
rect 516836 320832 516842 320884
rect 446490 320764 446496 320816
rect 446548 320804 446554 320816
rect 480070 320804 480076 320816
rect 446548 320776 480076 320804
rect 446548 320764 446554 320776
rect 480070 320764 480076 320776
rect 480128 320764 480134 320816
rect 447042 320696 447048 320748
rect 447100 320736 447106 320748
rect 482830 320736 482836 320748
rect 447100 320708 482836 320736
rect 447100 320696 447106 320708
rect 482830 320696 482836 320708
rect 482888 320696 482894 320748
rect 446398 320628 446404 320680
rect 446456 320668 446462 320680
rect 469858 320668 469864 320680
rect 446456 320640 469864 320668
rect 446456 320628 446462 320640
rect 469858 320628 469864 320640
rect 469916 320628 469922 320680
rect 507026 320492 507032 320544
rect 507084 320532 507090 320544
rect 509970 320532 509976 320544
rect 507084 320504 509976 320532
rect 507084 320492 507090 320504
rect 509970 320492 509976 320504
rect 510028 320492 510034 320544
rect 444282 320084 444288 320136
rect 444340 320124 444346 320136
rect 458542 320124 458548 320136
rect 444340 320096 458548 320124
rect 444340 320084 444346 320096
rect 458542 320084 458548 320096
rect 458600 320084 458606 320136
rect 469214 320084 469220 320136
rect 469272 320124 469278 320136
rect 472618 320124 472624 320136
rect 469272 320096 472624 320124
rect 469272 320084 469278 320096
rect 472618 320084 472624 320096
rect 472676 320084 472682 320136
rect 477034 320084 477040 320136
rect 477092 320124 477098 320136
rect 509142 320124 509148 320136
rect 477092 320096 509148 320124
rect 477092 320084 477098 320096
rect 509142 320084 509148 320096
rect 509200 320084 509206 320136
rect 445386 320016 445392 320068
rect 445444 320056 445450 320068
rect 461026 320056 461032 320068
rect 445444 320028 461032 320056
rect 445444 320016 445450 320028
rect 461026 320016 461032 320028
rect 461084 320016 461090 320068
rect 467098 320016 467104 320068
rect 467156 320056 467162 320068
rect 580810 320056 580816 320068
rect 467156 320028 580816 320056
rect 467156 320016 467162 320028
rect 580810 320016 580816 320028
rect 580868 320016 580874 320068
rect 449526 319948 449532 320000
rect 449584 319988 449590 320000
rect 461854 319988 461860 320000
rect 449584 319960 461860 319988
rect 449584 319948 449590 319960
rect 461854 319948 461860 319960
rect 461912 319948 461918 320000
rect 477862 319948 477868 320000
rect 477920 319988 477926 320000
rect 569310 319988 569316 320000
rect 477920 319960 569316 319988
rect 477920 319948 477926 319960
rect 569310 319948 569316 319960
rect 569368 319948 569374 320000
rect 443914 319880 443920 319932
rect 443972 319920 443978 319932
rect 461578 319920 461584 319932
rect 443972 319892 461584 319920
rect 443972 319880 443978 319892
rect 461578 319880 461584 319892
rect 461636 319880 461642 319932
rect 478690 319880 478696 319932
rect 478748 319920 478754 319932
rect 569218 319920 569224 319932
rect 478748 319892 569224 319920
rect 478748 319880 478754 319892
rect 569218 319880 569224 319892
rect 569276 319880 569282 319932
rect 442442 319812 442448 319864
rect 442500 319852 442506 319864
rect 471790 319852 471796 319864
rect 442500 319824 471796 319852
rect 442500 319812 442506 319824
rect 471790 319812 471796 319824
rect 471848 319812 471854 319864
rect 478414 319812 478420 319864
rect 478472 319852 478478 319864
rect 567930 319852 567936 319864
rect 478472 319824 567936 319852
rect 478472 319812 478478 319824
rect 567930 319812 567936 319824
rect 567988 319812 567994 319864
rect 468754 319744 468760 319796
rect 468812 319784 468818 319796
rect 515490 319784 515496 319796
rect 468812 319756 515496 319784
rect 468812 319744 468818 319756
rect 515490 319744 515496 319756
rect 515548 319744 515554 319796
rect 467926 319676 467932 319728
rect 467984 319716 467990 319728
rect 507946 319716 507952 319728
rect 467984 319688 507952 319716
rect 467984 319676 467990 319688
rect 507946 319676 507952 319688
rect 508004 319676 508010 319728
rect 468478 319608 468484 319660
rect 468536 319648 468542 319660
rect 507854 319648 507860 319660
rect 468536 319620 507860 319648
rect 468536 319608 468542 319620
rect 507854 319608 507860 319620
rect 507912 319608 507918 319660
rect 446674 319540 446680 319592
rect 446732 319580 446738 319592
rect 469582 319580 469588 319592
rect 446732 319552 469588 319580
rect 446732 319540 446738 319552
rect 469582 319540 469588 319552
rect 469640 319540 469646 319592
rect 477310 319540 477316 319592
rect 477368 319580 477374 319592
rect 514294 319580 514300 319592
rect 477368 319552 514300 319580
rect 477368 319540 477374 319552
rect 514294 319540 514300 319552
rect 514352 319540 514358 319592
rect 435634 319472 435640 319524
rect 435692 319512 435698 319524
rect 469122 319512 469128 319524
rect 435692 319484 469128 319512
rect 435692 319472 435698 319484
rect 469122 319472 469128 319484
rect 469180 319472 469186 319524
rect 469214 319472 469220 319524
rect 469272 319512 469278 319524
rect 472894 319512 472900 319524
rect 469272 319484 472900 319512
rect 469272 319472 469278 319484
rect 472894 319472 472900 319484
rect 472952 319472 472958 319524
rect 478966 319472 478972 319524
rect 479024 319512 479030 319524
rect 511350 319512 511356 319524
rect 479024 319484 511356 319512
rect 479024 319472 479030 319484
rect 511350 319472 511356 319484
rect 511408 319472 511414 319524
rect 460198 319404 460204 319456
rect 460256 319444 460262 319456
rect 474550 319444 474556 319456
rect 460256 319416 474556 319444
rect 460256 319404 460262 319416
rect 474550 319404 474556 319416
rect 474608 319404 474614 319456
rect 480806 319404 480812 319456
rect 480864 319444 480870 319456
rect 483106 319444 483112 319456
rect 480864 319416 483112 319444
rect 480864 319404 480870 319416
rect 483106 319404 483112 319416
rect 483164 319404 483170 319456
rect 502150 319404 502156 319456
rect 502208 319444 502214 319456
rect 543734 319444 543740 319456
rect 502208 319416 543740 319444
rect 502208 319404 502214 319416
rect 543734 319404 543740 319416
rect 543792 319404 543798 319456
rect 445294 319336 445300 319388
rect 445352 319376 445358 319388
rect 471514 319376 471520 319388
rect 445352 319348 471520 319376
rect 445352 319336 445358 319348
rect 471514 319336 471520 319348
rect 471572 319336 471578 319388
rect 478138 319336 478144 319388
rect 478196 319376 478202 319388
rect 510522 319376 510528 319388
rect 478196 319348 510528 319376
rect 478196 319336 478202 319348
rect 510522 319336 510528 319348
rect 510580 319336 510586 319388
rect 457162 319268 457168 319320
rect 457220 319308 457226 319320
rect 580718 319308 580724 319320
rect 457220 319280 580724 319308
rect 457220 319268 457226 319280
rect 580718 319268 580724 319280
rect 580776 319268 580782 319320
rect 446858 319200 446864 319252
rect 446916 319240 446922 319252
rect 480346 319240 480352 319252
rect 446916 319212 480352 319240
rect 446916 319200 446922 319212
rect 480346 319200 480352 319212
rect 480404 319200 480410 319252
rect 450538 319132 450544 319184
rect 450596 319172 450602 319184
rect 482002 319172 482008 319184
rect 450596 319144 482008 319172
rect 450596 319132 450602 319144
rect 482002 319132 482008 319144
rect 482060 319132 482066 319184
rect 450630 319064 450636 319116
rect 450688 319104 450694 319116
rect 479518 319104 479524 319116
rect 450688 319076 479524 319104
rect 450688 319064 450694 319076
rect 479518 319064 479524 319076
rect 479576 319064 479582 319116
rect 446582 318996 446588 319048
rect 446640 319036 446646 319048
rect 470134 319036 470140 319048
rect 446640 319008 470140 319036
rect 446640 318996 446646 319008
rect 470134 318996 470140 319008
rect 470192 318996 470198 319048
rect 454310 318928 454316 318980
rect 454368 318968 454374 318980
rect 454678 318968 454684 318980
rect 454368 318940 454684 318968
rect 454368 318928 454374 318940
rect 454678 318928 454684 318940
rect 454736 318928 454742 318980
rect 456886 318724 456892 318776
rect 456944 318764 456950 318776
rect 578878 318764 578884 318776
rect 456944 318736 578884 318764
rect 456944 318724 456950 318736
rect 578878 318724 578884 318736
rect 578936 318724 578942 318776
rect 457438 318656 457444 318708
rect 457496 318696 457502 318708
rect 577498 318696 577504 318708
rect 457496 318668 577504 318696
rect 457496 318656 457502 318668
rect 577498 318656 577504 318668
rect 577556 318656 577562 318708
rect 457714 318588 457720 318640
rect 457772 318628 457778 318640
rect 571978 318628 571984 318640
rect 457772 318600 571984 318628
rect 457772 318588 457778 318600
rect 571978 318588 571984 318600
rect 572036 318588 572042 318640
rect 438210 318520 438216 318572
rect 438268 318560 438274 318572
rect 470686 318560 470692 318572
rect 438268 318532 470692 318560
rect 438268 318520 438274 318532
rect 470686 318520 470692 318532
rect 470744 318520 470750 318572
rect 441154 318452 441160 318504
rect 441212 318492 441218 318504
rect 470410 318492 470416 318504
rect 441212 318464 470416 318492
rect 441212 318452 441218 318464
rect 470410 318452 470416 318464
rect 470468 318452 470474 318504
rect 449434 318384 449440 318436
rect 449492 318424 449498 318436
rect 472066 318424 472072 318436
rect 449492 318396 472072 318424
rect 449492 318384 449498 318396
rect 472066 318384 472072 318396
rect 472124 318384 472130 318436
rect 458818 318112 458824 318164
rect 458876 318152 458882 318164
rect 486970 318152 486976 318164
rect 458876 318124 486976 318152
rect 458876 318112 458882 318124
rect 486970 318112 486976 318124
rect 487028 318112 487034 318164
rect 457438 318044 457444 318096
rect 457496 318084 457502 318096
rect 489178 318084 489184 318096
rect 457496 318056 489184 318084
rect 457496 318044 457502 318056
rect 489178 318044 489184 318056
rect 489236 318044 489242 318096
rect 494422 318044 494428 318096
rect 494480 318084 494486 318096
rect 540974 318084 540980 318096
rect 494480 318056 540980 318084
rect 494480 318044 494486 318056
rect 540974 318044 540980 318056
rect 541032 318044 541038 318096
rect 443822 317364 443828 317416
rect 443880 317404 443886 317416
rect 481726 317404 481732 317416
rect 443880 317376 481732 317404
rect 443880 317364 443886 317376
rect 481726 317364 481732 317376
rect 481784 317364 481790 317416
rect 446950 317296 446956 317348
rect 447008 317336 447014 317348
rect 481174 317336 481180 317348
rect 447008 317308 481180 317336
rect 447008 317296 447014 317308
rect 481174 317296 481180 317308
rect 481232 317296 481238 317348
rect 480254 317228 480260 317280
rect 480312 317268 480318 317280
rect 483382 317268 483388 317280
rect 480312 317240 483388 317268
rect 480312 317228 480318 317240
rect 483382 317228 483388 317240
rect 483440 317228 483446 317280
rect 467098 317160 467104 317212
rect 467156 317200 467162 317212
rect 469214 317200 469220 317212
rect 467156 317172 469220 317200
rect 467156 317160 467162 317172
rect 469214 317160 469220 317172
rect 469272 317160 469278 317212
rect 473446 317160 473452 317212
rect 473504 317200 473510 317212
rect 473906 317200 473912 317212
rect 473504 317172 473912 317200
rect 473504 317160 473510 317172
rect 473906 317160 473912 317172
rect 473964 317160 473970 317212
rect 501598 317024 501604 317076
rect 501656 317064 501662 317076
rect 539134 317064 539140 317076
rect 501656 317036 539140 317064
rect 501656 317024 501662 317036
rect 539134 317024 539140 317036
rect 539192 317024 539198 317076
rect 499666 316956 499672 317008
rect 499724 316996 499730 317008
rect 542446 316996 542452 317008
rect 499724 316968 542452 316996
rect 499724 316956 499730 316968
rect 542446 316956 542452 316968
rect 542504 316956 542510 317008
rect 472618 316888 472624 316940
rect 472676 316928 472682 316940
rect 480806 316928 480812 316940
rect 472676 316900 480812 316928
rect 472676 316888 472682 316900
rect 480806 316888 480812 316900
rect 480864 316888 480870 316940
rect 497182 316888 497188 316940
rect 497240 316928 497246 316940
rect 541066 316928 541072 316940
rect 497240 316900 541072 316928
rect 497240 316888 497246 316900
rect 541066 316888 541072 316900
rect 541124 316888 541130 316940
rect 459002 316820 459008 316872
rect 459060 316860 459066 316872
rect 492214 316860 492220 316872
rect 459060 316832 492220 316860
rect 459060 316820 459066 316832
rect 492214 316820 492220 316832
rect 492272 316820 492278 316872
rect 496078 316820 496084 316872
rect 496136 316860 496142 316872
rect 543182 316860 543188 316872
rect 496136 316832 543188 316860
rect 496136 316820 496142 316832
rect 543182 316820 543188 316832
rect 543240 316820 543246 316872
rect 454770 316752 454776 316804
rect 454828 316792 454834 316804
rect 502426 316792 502432 316804
rect 454828 316764 502432 316792
rect 454828 316752 454834 316764
rect 502426 316752 502432 316764
rect 502484 316752 502490 316804
rect 456058 316684 456064 316736
rect 456116 316724 456122 316736
rect 461578 316724 461584 316736
rect 456116 316696 461584 316724
rect 456116 316684 456122 316696
rect 461578 316684 461584 316696
rect 461636 316684 461642 316736
rect 502978 316724 502984 316736
rect 470566 316696 502984 316724
rect 454678 316616 454684 316668
rect 454736 316656 454742 316668
rect 470566 316656 470594 316696
rect 502978 316684 502984 316696
rect 503036 316684 503042 316736
rect 454736 316628 470594 316656
rect 454736 316616 454742 316628
rect 361758 315936 361764 315988
rect 361816 315976 361822 315988
rect 399478 315976 399484 315988
rect 361816 315948 399484 315976
rect 361816 315936 361822 315948
rect 399478 315936 399484 315948
rect 399536 315936 399542 315988
rect 447778 315528 447784 315580
rect 447836 315568 447842 315580
rect 456886 315568 456892 315580
rect 447836 315540 456892 315568
rect 447836 315528 447842 315540
rect 456886 315528 456892 315540
rect 456944 315528 456950 315580
rect 501046 315528 501052 315580
rect 501104 315568 501110 315580
rect 542722 315568 542728 315580
rect 501104 315540 542728 315568
rect 501104 315528 501110 315540
rect 542722 315528 542728 315540
rect 542780 315528 542786 315580
rect 453390 315460 453396 315512
rect 453448 315500 453454 315512
rect 494146 315500 494152 315512
rect 453448 315472 494152 315500
rect 453448 315460 453454 315472
rect 494146 315460 494152 315472
rect 494204 315460 494210 315512
rect 498286 315460 498292 315512
rect 498344 315500 498350 315512
rect 541158 315500 541164 315512
rect 498344 315472 541164 315500
rect 498344 315460 498350 315472
rect 541158 315460 541164 315472
rect 541216 315460 541222 315512
rect 450630 315392 450636 315444
rect 450688 315432 450694 315444
rect 504082 315432 504088 315444
rect 450688 315404 504088 315432
rect 450688 315392 450694 315404
rect 504082 315392 504088 315404
rect 504140 315392 504146 315444
rect 450538 315324 450544 315376
rect 450596 315364 450602 315376
rect 503806 315364 503812 315376
rect 450596 315336 503812 315364
rect 450596 315324 450602 315336
rect 503806 315324 503812 315336
rect 503864 315324 503870 315376
rect 455506 315256 455512 315308
rect 455564 315296 455570 315308
rect 570598 315296 570604 315308
rect 455564 315268 570604 315296
rect 455564 315256 455570 315268
rect 570598 315256 570604 315268
rect 570656 315256 570662 315308
rect 457622 314644 457628 314696
rect 457680 314684 457686 314696
rect 462406 314684 462412 314696
rect 457680 314656 462412 314684
rect 457680 314644 457686 314656
rect 462406 314644 462412 314656
rect 462464 314644 462470 314696
rect 433242 314508 433248 314560
rect 433300 314548 433306 314560
rect 441062 314548 441068 314560
rect 433300 314520 441068 314548
rect 433300 314508 433306 314520
rect 441062 314508 441068 314520
rect 441120 314508 441126 314560
rect 451918 313964 451924 314016
rect 451976 314004 451982 314016
rect 487246 314004 487252 314016
rect 451976 313976 487252 314004
rect 451976 313964 451982 313976
rect 487246 313964 487252 313976
rect 487304 313964 487310 314016
rect 496630 313964 496636 314016
rect 496688 314004 496694 314016
rect 539594 314004 539600 314016
rect 496688 313976 539600 314004
rect 496688 313964 496694 313976
rect 539594 313964 539600 313976
rect 539652 313964 539658 314016
rect 485590 313896 485596 313948
rect 485648 313936 485654 313948
rect 529934 313936 529940 313948
rect 485648 313908 529940 313936
rect 485648 313896 485654 313908
rect 529934 313896 529940 313908
rect 529992 313896 529998 313948
rect 466546 313216 466552 313268
rect 466604 313256 466610 313268
rect 580166 313256 580172 313268
rect 466604 313228 580172 313256
rect 466604 313216 466610 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 465166 312536 465172 312588
rect 465224 312576 465230 312588
rect 551278 312576 551284 312588
rect 465224 312548 551284 312576
rect 465224 312536 465230 312548
rect 551278 312536 551284 312548
rect 551336 312536 551342 312588
rect 478138 312400 478144 312452
rect 478196 312440 478202 312452
rect 480254 312440 480260 312452
rect 478196 312412 480260 312440
rect 478196 312400 478202 312412
rect 480254 312400 480260 312412
rect 480312 312400 480318 312452
rect 452102 311176 452108 311228
rect 452160 311216 452166 311228
rect 492766 311216 492772 311228
rect 452160 311188 492772 311216
rect 452160 311176 452166 311188
rect 492766 311176 492772 311188
rect 492824 311176 492830 311228
rect 475378 311108 475384 311160
rect 475436 311148 475442 311160
rect 544378 311148 544384 311160
rect 475436 311120 544384 311148
rect 475436 311108 475442 311120
rect 544378 311108 544384 311120
rect 544436 311108 544442 311160
rect 453298 309816 453304 309868
rect 453356 309856 453362 309868
rect 488350 309856 488356 309868
rect 453356 309828 488356 309856
rect 453356 309816 453362 309828
rect 488350 309816 488356 309828
rect 488408 309816 488414 309868
rect 475102 309748 475108 309800
rect 475160 309788 475166 309800
rect 563698 309788 563704 309800
rect 475160 309760 563704 309788
rect 475160 309748 475166 309760
rect 563698 309748 563704 309760
rect 563756 309748 563762 309800
rect 458910 308456 458916 308508
rect 458968 308496 458974 308508
rect 488626 308496 488632 308508
rect 458968 308468 488632 308496
rect 458968 308456 458974 308468
rect 488626 308456 488632 308468
rect 488684 308456 488690 308508
rect 464614 308388 464620 308440
rect 464672 308428 464678 308440
rect 562318 308428 562324 308440
rect 464672 308400 562324 308428
rect 464672 308388 464678 308400
rect 562318 308388 562324 308400
rect 562376 308388 562382 308440
rect 432230 307708 432236 307760
rect 432288 307748 432294 307760
rect 436830 307748 436836 307760
rect 432288 307720 436836 307748
rect 432288 307708 432294 307720
rect 436830 307708 436836 307720
rect 436888 307708 436894 307760
rect 381630 306280 381636 306332
rect 381688 306320 381694 306332
rect 463510 306320 463516 306332
rect 381688 306292 463516 306320
rect 381688 306280 381694 306292
rect 463510 306280 463516 306292
rect 463568 306280 463574 306332
rect 385862 306212 385868 306264
rect 385920 306252 385926 306264
rect 474274 306252 474280 306264
rect 385920 306224 474280 306252
rect 385920 306212 385926 306224
rect 474274 306212 474280 306224
rect 474332 306212 474338 306264
rect 384574 306144 384580 306196
rect 384632 306184 384638 306196
rect 473998 306184 474004 306196
rect 384632 306156 474004 306184
rect 384632 306144 384638 306156
rect 473998 306144 474004 306156
rect 474056 306144 474062 306196
rect 381722 306076 381728 306128
rect 381780 306116 381786 306128
rect 473722 306116 473728 306128
rect 381780 306088 473728 306116
rect 381780 306076 381786 306088
rect 473722 306076 473728 306088
rect 473780 306076 473786 306128
rect 384758 306008 384764 306060
rect 384816 306048 384822 306060
rect 484762 306048 484768 306060
rect 384816 306020 484768 306048
rect 384816 306008 384822 306020
rect 484762 306008 484768 306020
rect 484820 306008 484826 306060
rect 384850 305940 384856 305992
rect 384908 305980 384914 305992
rect 484486 305980 484492 305992
rect 384908 305952 484492 305980
rect 384908 305940 384914 305952
rect 484486 305940 484492 305952
rect 484544 305940 484550 305992
rect 381538 305872 381544 305924
rect 381596 305912 381602 305924
rect 484210 305912 484216 305924
rect 381596 305884 484216 305912
rect 381596 305872 381602 305884
rect 484210 305872 484216 305884
rect 484268 305872 484274 305924
rect 374638 305804 374644 305856
rect 374696 305844 374702 305856
rect 485314 305844 485320 305856
rect 374696 305816 485320 305844
rect 374696 305804 374702 305816
rect 485314 305804 485320 305816
rect 485372 305804 485378 305856
rect 426342 305736 426348 305788
rect 426400 305776 426406 305788
rect 441614 305776 441620 305788
rect 426400 305748 441620 305776
rect 426400 305736 426406 305748
rect 441614 305736 441620 305748
rect 441672 305736 441678 305788
rect 454218 305736 454224 305788
rect 454276 305776 454282 305788
rect 565078 305776 565084 305788
rect 454276 305748 565084 305776
rect 454276 305736 454282 305748
rect 565078 305736 565084 305748
rect 565136 305736 565142 305788
rect 360930 305668 360936 305720
rect 360988 305708 360994 305720
rect 512178 305708 512184 305720
rect 360988 305680 512184 305708
rect 360988 305668 360994 305680
rect 512178 305668 512184 305680
rect 512236 305668 512242 305720
rect 359458 305600 359464 305652
rect 359516 305640 359522 305652
rect 512546 305640 512552 305652
rect 359516 305612 512552 305640
rect 359516 305600 359522 305612
rect 512546 305600 512552 305612
rect 512604 305600 512610 305652
rect 384390 305532 384396 305584
rect 384448 305572 384454 305584
rect 464062 305572 464068 305584
rect 384448 305544 464068 305572
rect 384448 305532 384454 305544
rect 464062 305532 464068 305544
rect 464120 305532 464126 305584
rect 385770 305464 385776 305516
rect 385828 305504 385834 305516
rect 463786 305504 463792 305516
rect 385828 305476 463792 305504
rect 385828 305464 385834 305476
rect 463786 305464 463792 305476
rect 463844 305464 463850 305516
rect 457530 305396 457536 305448
rect 457588 305436 457594 305448
rect 490006 305436 490012 305448
rect 457588 305408 490012 305436
rect 457588 305396 457594 305408
rect 490006 305396 490012 305408
rect 490064 305396 490070 305448
rect 3418 304988 3424 305040
rect 3476 305028 3482 305040
rect 4798 305028 4804 305040
rect 3476 305000 4804 305028
rect 3476 304988 3482 305000
rect 4798 304988 4804 305000
rect 4856 304988 4862 305040
rect 361758 304920 361764 304972
rect 361816 304960 361822 304972
rect 443730 304960 443736 304972
rect 361816 304932 443736 304960
rect 361816 304920 361822 304932
rect 443730 304920 443736 304932
rect 443788 304920 443794 304972
rect 455782 304444 455788 304496
rect 455840 304484 455846 304496
rect 573358 304484 573364 304496
rect 455840 304456 573364 304484
rect 455840 304444 455846 304456
rect 573358 304444 573364 304456
rect 573416 304444 573422 304496
rect 385678 304376 385684 304428
rect 385736 304416 385742 304428
rect 519722 304416 519728 304428
rect 385736 304388 519728 304416
rect 385736 304376 385742 304388
rect 519722 304376 519728 304388
rect 519780 304376 519786 304428
rect 361022 304308 361028 304360
rect 361080 304348 361086 304360
rect 512822 304348 512828 304360
rect 361080 304320 512828 304348
rect 361080 304308 361086 304320
rect 512822 304308 512828 304320
rect 512880 304308 512886 304360
rect 359550 304240 359556 304292
rect 359608 304280 359614 304292
rect 512362 304280 512368 304292
rect 359608 304252 512368 304280
rect 359608 304240 359614 304252
rect 512362 304240 512368 304252
rect 512420 304240 512426 304292
rect 378686 303560 378692 303612
rect 378744 303600 378750 303612
rect 483934 303600 483940 303612
rect 378744 303572 483940 303600
rect 378744 303560 378750 303572
rect 483934 303560 483940 303572
rect 483992 303560 483998 303612
rect 485866 303560 485872 303612
rect 485924 303600 485930 303612
rect 530026 303600 530032 303612
rect 485924 303572 530032 303600
rect 485924 303560 485930 303572
rect 530026 303560 530032 303572
rect 530084 303560 530090 303612
rect 381998 303492 382004 303544
rect 382056 303532 382062 303544
rect 511442 303532 511448 303544
rect 382056 303504 511448 303532
rect 382056 303492 382062 303504
rect 511442 303492 511448 303504
rect 511500 303492 511506 303544
rect 379054 303424 379060 303476
rect 379112 303464 379118 303476
rect 509510 303464 509516 303476
rect 379112 303436 509516 303464
rect 379112 303424 379118 303436
rect 509510 303424 509516 303436
rect 509568 303424 509574 303476
rect 376018 303356 376024 303408
rect 376076 303396 376082 303408
rect 506934 303396 506940 303408
rect 376076 303368 506940 303396
rect 376076 303356 376082 303368
rect 506934 303356 506940 303368
rect 506992 303356 506998 303408
rect 379238 303288 379244 303340
rect 379296 303328 379302 303340
rect 511074 303328 511080 303340
rect 379296 303300 511080 303328
rect 379296 303288 379302 303300
rect 511074 303288 511080 303300
rect 511132 303288 511138 303340
rect 382090 303220 382096 303272
rect 382148 303260 382154 303272
rect 515306 303260 515312 303272
rect 382148 303232 515312 303260
rect 382148 303220 382154 303232
rect 515306 303220 515312 303232
rect 515364 303220 515370 303272
rect 376202 303152 376208 303204
rect 376260 303192 376266 303204
rect 509418 303192 509424 303204
rect 376260 303164 509424 303192
rect 376260 303152 376266 303164
rect 509418 303152 509424 303164
rect 509476 303152 509482 303204
rect 379330 303084 379336 303136
rect 379388 303124 379394 303136
rect 513926 303124 513932 303136
rect 379388 303096 513932 303124
rect 379388 303084 379394 303096
rect 513926 303084 513932 303096
rect 513984 303084 513990 303136
rect 379146 303016 379152 303068
rect 379204 303056 379210 303068
rect 515122 303056 515128 303068
rect 379204 303028 515128 303056
rect 379204 303016 379210 303028
rect 515122 303016 515128 303028
rect 515180 303016 515186 303068
rect 378962 302948 378968 303000
rect 379020 302988 379026 303000
rect 515214 302988 515220 303000
rect 379020 302960 515220 302988
rect 379020 302948 379026 302960
rect 515214 302948 515220 302960
rect 515272 302948 515278 303000
rect 373258 302880 373264 302932
rect 373316 302920 373322 302932
rect 513558 302920 513564 302932
rect 373316 302892 513564 302920
rect 373316 302880 373322 302892
rect 513558 302880 513564 302892
rect 513616 302880 513622 302932
rect 379422 302812 379428 302864
rect 379480 302852 379486 302864
rect 473906 302852 473912 302864
rect 379480 302824 473912 302852
rect 379480 302812 379486 302824
rect 473906 302812 473912 302824
rect 473964 302812 473970 302864
rect 381446 302744 381452 302796
rect 381504 302784 381510 302796
rect 463234 302784 463240 302796
rect 381504 302756 463240 302784
rect 381504 302744 381510 302756
rect 463234 302744 463240 302756
rect 463292 302744 463298 302796
rect 386138 302676 386144 302728
rect 386196 302716 386202 302728
rect 462958 302716 462964 302728
rect 386196 302688 462964 302716
rect 386196 302676 386202 302688
rect 462958 302676 462964 302688
rect 463016 302676 463022 302728
rect 486418 301588 486424 301640
rect 486476 301628 486482 301640
rect 529198 301628 529204 301640
rect 486476 301600 529204 301628
rect 486476 301588 486482 301600
rect 529198 301588 529204 301600
rect 529256 301588 529262 301640
rect 378778 301520 378784 301572
rect 378836 301560 378842 301572
rect 464338 301560 464344 301572
rect 378836 301532 464344 301560
rect 378836 301520 378842 301532
rect 464338 301520 464344 301532
rect 464396 301520 464402 301572
rect 465718 301520 465724 301572
rect 465776 301560 465782 301572
rect 537478 301560 537484 301572
rect 465776 301532 537484 301560
rect 465776 301520 465782 301532
rect 537478 301520 537484 301532
rect 537536 301520 537542 301572
rect 407114 301452 407120 301504
rect 407172 301492 407178 301504
rect 502702 301492 502708 301504
rect 407172 301464 502708 301492
rect 407172 301452 407178 301464
rect 502702 301452 502708 301464
rect 502760 301452 502766 301504
rect 376294 300772 376300 300824
rect 376352 300812 376358 300824
rect 510982 300812 510988 300824
rect 376352 300784 510988 300812
rect 376352 300772 376358 300784
rect 510982 300772 510988 300784
rect 511040 300772 511046 300824
rect 373626 300704 373632 300756
rect 373684 300744 373690 300756
rect 511534 300744 511540 300756
rect 373684 300716 511540 300744
rect 373684 300704 373690 300716
rect 511534 300704 511540 300716
rect 511592 300704 511598 300756
rect 376386 300636 376392 300688
rect 376444 300676 376450 300688
rect 513742 300676 513748 300688
rect 376444 300648 513748 300676
rect 376444 300636 376450 300648
rect 513742 300636 513748 300648
rect 513800 300636 513806 300688
rect 368290 300568 368296 300620
rect 368348 300608 368354 300620
rect 507026 300608 507032 300620
rect 368348 300580 507032 300608
rect 368348 300568 368354 300580
rect 507026 300568 507032 300580
rect 507084 300568 507090 300620
rect 373534 300500 373540 300552
rect 373592 300540 373598 300552
rect 513466 300540 513472 300552
rect 373592 300512 513472 300540
rect 373592 300500 373598 300512
rect 513466 300500 513472 300512
rect 513524 300500 513530 300552
rect 373442 300432 373448 300484
rect 373500 300472 373506 300484
rect 514938 300472 514944 300484
rect 373500 300444 514944 300472
rect 373500 300432 373506 300444
rect 514938 300432 514944 300444
rect 514996 300432 515002 300484
rect 370866 300364 370872 300416
rect 370924 300404 370930 300416
rect 514846 300404 514852 300416
rect 370924 300376 514852 300404
rect 370924 300364 370930 300376
rect 514846 300364 514852 300376
rect 514904 300364 514910 300416
rect 371050 300296 371056 300348
rect 371108 300336 371114 300348
rect 516134 300336 516140 300348
rect 371108 300308 516140 300336
rect 371108 300296 371114 300308
rect 516134 300296 516140 300308
rect 516192 300296 516198 300348
rect 370958 300228 370964 300280
rect 371016 300268 371022 300280
rect 517698 300268 517704 300280
rect 371016 300240 517704 300268
rect 371016 300228 371022 300240
rect 517698 300228 517704 300240
rect 517756 300228 517762 300280
rect 370774 300160 370780 300212
rect 370832 300200 370838 300212
rect 517514 300200 517520 300212
rect 370832 300172 517520 300200
rect 370832 300160 370838 300172
rect 517514 300160 517520 300172
rect 517572 300160 517578 300212
rect 368106 300092 368112 300144
rect 368164 300132 368170 300144
rect 518342 300132 518348 300144
rect 368164 300104 518348 300132
rect 368164 300092 368170 300104
rect 518342 300092 518348 300104
rect 518400 300092 518406 300144
rect 376478 300024 376484 300076
rect 376536 300064 376542 300076
rect 509326 300064 509332 300076
rect 376536 300036 509332 300064
rect 376536 300024 376542 300036
rect 509326 300024 509332 300036
rect 509384 300024 509390 300076
rect 378594 299956 378600 300008
rect 378652 299996 378658 300008
rect 483658 299996 483664 300008
rect 378652 299968 483664 299996
rect 378652 299956 378658 299968
rect 483658 299956 483664 299968
rect 483716 299956 483722 300008
rect 376662 299888 376668 299940
rect 376720 299928 376726 299940
rect 473170 299928 473176 299940
rect 376720 299900 473176 299928
rect 376720 299888 376726 299900
rect 473170 299888 473176 299900
rect 473228 299888 473234 299940
rect 461578 299412 461584 299464
rect 461636 299452 461642 299464
rect 580166 299452 580172 299464
rect 461636 299424 580172 299452
rect 461636 299412 461642 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 376570 298800 376576 298852
rect 376628 298840 376634 298852
rect 485038 298840 485044 298852
rect 376628 298812 485044 298840
rect 376628 298800 376634 298812
rect 485038 298800 485044 298812
rect 485096 298800 485102 298852
rect 371970 298732 371976 298784
rect 372028 298772 372034 298784
rect 513190 298772 513196 298784
rect 372028 298744 513196 298772
rect 372028 298732 372034 298744
rect 513190 298732 513196 298744
rect 513248 298732 513254 298784
rect 365162 298052 365168 298104
rect 365220 298092 365226 298104
rect 507578 298092 507584 298104
rect 365220 298064 507584 298092
rect 365220 298052 365226 298064
rect 507578 298052 507584 298064
rect 507636 298052 507642 298104
rect 367830 297984 367836 298036
rect 367888 298024 367894 298036
rect 514110 298024 514116 298036
rect 367888 297996 514116 298024
rect 367888 297984 367894 297996
rect 514110 297984 514116 297996
rect 514168 297984 514174 298036
rect 363598 297916 363604 297968
rect 363656 297956 363662 297968
rect 512270 297956 512276 297968
rect 363656 297928 512276 297956
rect 363656 297916 363662 297928
rect 512270 297916 512276 297928
rect 512328 297916 512334 297968
rect 367922 297848 367928 297900
rect 367980 297888 367986 297900
rect 516962 297888 516968 297900
rect 367980 297860 516968 297888
rect 367980 297848 367986 297860
rect 516962 297848 516968 297860
rect 517020 297848 517026 297900
rect 365070 297780 365076 297832
rect 365128 297820 365134 297832
rect 515582 297820 515588 297832
rect 365128 297792 515588 297820
rect 365128 297780 365134 297792
rect 515582 297780 515588 297792
rect 515640 297780 515646 297832
rect 361206 297712 361212 297764
rect 361264 297752 361270 297764
rect 512086 297752 512092 297764
rect 361264 297724 512092 297752
rect 361264 297712 361270 297724
rect 512086 297712 512092 297724
rect 512144 297712 512150 297764
rect 365530 297644 365536 297696
rect 365588 297684 365594 297696
rect 516870 297684 516876 297696
rect 365588 297656 516876 297684
rect 365588 297644 365594 297656
rect 516870 297644 516876 297656
rect 516928 297644 516934 297696
rect 365254 297576 365260 297628
rect 365312 297616 365318 297628
rect 516686 297616 516692 297628
rect 365312 297588 516692 297616
rect 365312 297576 365318 297588
rect 516686 297576 516692 297588
rect 516744 297576 516750 297628
rect 362310 297508 362316 297560
rect 362368 297548 362374 297560
rect 513834 297548 513840 297560
rect 362368 297520 513840 297548
rect 362368 297508 362374 297520
rect 513834 297508 513840 297520
rect 513892 297508 513898 297560
rect 365438 297440 365444 297492
rect 365496 297480 365502 297492
rect 518250 297480 518256 297492
rect 365496 297452 518256 297480
rect 365496 297440 365502 297452
rect 518250 297440 518256 297452
rect 518308 297440 518314 297492
rect 362218 297372 362224 297424
rect 362276 297412 362282 297424
rect 518066 297412 518072 297424
rect 362276 297384 518072 297412
rect 362276 297372 362282 297384
rect 518066 297372 518072 297384
rect 518124 297372 518130 297424
rect 365346 297304 365352 297356
rect 365404 297344 365410 297356
rect 507762 297344 507768 297356
rect 365404 297316 507768 297344
rect 365404 297304 365410 297316
rect 507762 297304 507768 297316
rect 507820 297304 507826 297356
rect 382918 297236 382924 297288
rect 382976 297276 382982 297288
rect 518158 297276 518164 297288
rect 382976 297248 518164 297276
rect 382976 297236 382982 297248
rect 518158 297236 518164 297248
rect 518216 297236 518222 297288
rect 464338 297168 464344 297220
rect 464396 297208 464402 297220
rect 467098 297208 467104 297220
rect 464396 297180 467104 297208
rect 464396 297168 464402 297180
rect 467098 297168 467104 297180
rect 467156 297168 467162 297220
rect 476206 297168 476212 297220
rect 476264 297208 476270 297220
rect 548518 297208 548524 297220
rect 476264 297180 548524 297208
rect 476264 297168 476270 297180
rect 548518 297168 548524 297180
rect 548576 297168 548582 297220
rect 454402 295944 454408 295996
rect 454460 295984 454466 295996
rect 578878 295984 578884 295996
rect 454460 295956 578884 295984
rect 454460 295944 454466 295956
rect 578878 295944 578884 295956
rect 578936 295944 578942 295996
rect 369210 295264 369216 295316
rect 369268 295304 369274 295316
rect 514754 295304 514760 295316
rect 369268 295276 514760 295304
rect 369268 295264 369274 295276
rect 514754 295264 514760 295276
rect 514812 295264 514818 295316
rect 366634 295196 366640 295248
rect 366692 295236 366698 295248
rect 514202 295236 514208 295248
rect 366692 295208 514208 295236
rect 366692 295196 366698 295208
rect 514202 295196 514208 295208
rect 514260 295196 514266 295248
rect 369118 295128 369124 295180
rect 369176 295168 369182 295180
rect 516226 295168 516232 295180
rect 369176 295140 516232 295168
rect 369176 295128 369182 295140
rect 516226 295128 516232 295140
rect 516284 295128 516290 295180
rect 366450 295060 366456 295112
rect 366508 295100 366514 295112
rect 513650 295100 513656 295112
rect 366508 295072 513656 295100
rect 366508 295060 366514 295072
rect 513650 295060 513656 295072
rect 513708 295060 513714 295112
rect 361298 294992 361304 295044
rect 361356 295032 361362 295044
rect 510890 295032 510896 295044
rect 361356 295004 510896 295032
rect 361356 294992 361362 295004
rect 510890 294992 510896 295004
rect 510948 294992 510954 295044
rect 369302 294924 369308 294976
rect 369360 294964 369366 294976
rect 518986 294964 518992 294976
rect 369360 294936 518992 294964
rect 369360 294924 369366 294936
rect 518986 294924 518992 294936
rect 519044 294924 519050 294976
rect 366726 294856 366732 294908
rect 366784 294896 366790 294908
rect 517790 294896 517796 294908
rect 366784 294868 517796 294896
rect 366784 294856 366790 294868
rect 517790 294856 517796 294868
rect 517848 294856 517854 294908
rect 363966 294788 363972 294840
rect 364024 294828 364030 294840
rect 516410 294828 516416 294840
rect 364024 294800 516416 294828
rect 364024 294788 364030 294800
rect 516410 294788 516416 294800
rect 516468 294788 516474 294840
rect 363874 294720 363880 294772
rect 363932 294760 363938 294772
rect 517882 294760 517888 294772
rect 363932 294732 517888 294760
rect 363932 294720 363938 294732
rect 517882 294720 517888 294732
rect 517940 294720 517946 294772
rect 362402 294652 362408 294704
rect 362460 294692 362466 294704
rect 516594 294692 516600 294704
rect 362460 294664 516600 294692
rect 362460 294652 362466 294664
rect 516594 294652 516600 294664
rect 516652 294652 516658 294704
rect 362494 294584 362500 294636
rect 362552 294624 362558 294636
rect 517974 294624 517980 294636
rect 362552 294596 517980 294624
rect 362552 294584 362558 294596
rect 517974 294584 517980 294596
rect 518032 294584 518038 294636
rect 366542 294516 366548 294568
rect 366600 294556 366606 294568
rect 510706 294556 510712 294568
rect 366600 294528 510712 294556
rect 366600 294516 366606 294528
rect 510706 294516 510712 294528
rect 510764 294516 510770 294568
rect 368198 294448 368204 294500
rect 368256 294488 368262 294500
rect 509786 294488 509792 294500
rect 368256 294460 509792 294488
rect 368256 294448 368262 294460
rect 509786 294448 509792 294460
rect 509844 294448 509850 294500
rect 454310 294380 454316 294432
rect 454368 294420 454374 294432
rect 576118 294420 576124 294432
rect 454368 294392 576124 294420
rect 454368 294380 454374 294392
rect 576118 294380 576124 294392
rect 576176 294380 576182 294432
rect 361758 293904 361764 293956
rect 361816 293944 361822 293956
rect 385954 293944 385960 293956
rect 361816 293916 385960 293944
rect 361816 293904 361822 293916
rect 385954 293904 385960 293916
rect 386012 293904 386018 293956
rect 459094 293292 459100 293344
rect 459152 293332 459158 293344
rect 488902 293332 488908 293344
rect 459152 293304 488908 293332
rect 459152 293292 459158 293304
rect 488902 293292 488908 293304
rect 488960 293292 488966 293344
rect 475930 293224 475936 293276
rect 475988 293264 475994 293276
rect 536098 293264 536104 293276
rect 475988 293236 536104 293264
rect 475988 293224 475994 293236
rect 536098 293224 536104 293236
rect 536156 293224 536162 293276
rect 3510 292748 3516 292800
rect 3568 292788 3574 292800
rect 4890 292788 4896 292800
rect 3568 292760 4896 292788
rect 3568 292748 3574 292760
rect 4890 292748 4896 292760
rect 4948 292748 4954 292800
rect 375098 292476 375104 292528
rect 375156 292516 375162 292528
rect 507394 292516 507400 292528
rect 375156 292488 507400 292516
rect 375156 292476 375162 292488
rect 507394 292476 507400 292488
rect 507452 292476 507458 292528
rect 381814 292408 381820 292460
rect 381872 292448 381878 292460
rect 519170 292448 519176 292460
rect 381872 292420 519176 292448
rect 381872 292408 381878 292420
rect 519170 292408 519176 292420
rect 519228 292408 519234 292460
rect 380158 292340 380164 292392
rect 380216 292380 380222 292392
rect 520642 292380 520648 292392
rect 380216 292352 520648 292380
rect 380216 292340 380222 292352
rect 520642 292340 520648 292352
rect 520700 292340 520706 292392
rect 380250 292272 380256 292324
rect 380308 292312 380314 292324
rect 520734 292312 520740 292324
rect 380308 292284 520740 292312
rect 380308 292272 380314 292284
rect 520734 292272 520740 292284
rect 520792 292272 520798 292324
rect 377582 292204 377588 292256
rect 377640 292244 377646 292256
rect 519262 292244 519268 292256
rect 377640 292216 519268 292244
rect 377640 292204 377646 292216
rect 519262 292204 519268 292216
rect 519320 292204 519326 292256
rect 377398 292136 377404 292188
rect 377456 292176 377462 292188
rect 520826 292176 520832 292188
rect 377456 292148 520832 292176
rect 377456 292136 377462 292148
rect 520826 292136 520832 292148
rect 520884 292136 520890 292188
rect 375006 292068 375012 292120
rect 375064 292108 375070 292120
rect 519446 292108 519452 292120
rect 375064 292080 519452 292108
rect 375064 292068 375070 292080
rect 519446 292068 519452 292080
rect 519504 292068 519510 292120
rect 374730 292000 374736 292052
rect 374788 292040 374794 292052
rect 519630 292040 519636 292052
rect 374788 292012 519636 292040
rect 374788 292000 374794 292012
rect 519630 292000 519636 292012
rect 519688 292000 519694 292052
rect 374914 291932 374920 291984
rect 374972 291972 374978 291984
rect 520918 291972 520924 291984
rect 374972 291944 520924 291972
rect 374972 291932 374978 291944
rect 520918 291932 520924 291944
rect 520976 291932 520982 291984
rect 372246 291864 372252 291916
rect 372304 291904 372310 291916
rect 518894 291904 518900 291916
rect 372304 291876 518900 291904
rect 372304 291864 372310 291876
rect 518894 291864 518900 291876
rect 518952 291864 518958 291916
rect 372338 291796 372344 291848
rect 372396 291836 372402 291848
rect 520274 291836 520280 291848
rect 372396 291808 520280 291836
rect 372396 291796 372402 291808
rect 520274 291796 520280 291808
rect 520332 291796 520338 291848
rect 377674 291728 377680 291780
rect 377732 291768 377738 291780
rect 507670 291768 507676 291780
rect 377732 291740 507676 291768
rect 377732 291728 377738 291740
rect 507670 291728 507676 291740
rect 507728 291728 507734 291780
rect 454954 291660 454960 291712
rect 455012 291700 455018 291712
rect 574738 291700 574744 291712
rect 455012 291672 574744 291700
rect 455012 291660 455018 291672
rect 574738 291660 574744 291672
rect 574796 291660 574802 291712
rect 455230 290436 455236 290488
rect 455288 290476 455294 290488
rect 533338 290476 533344 290488
rect 455288 290448 533344 290476
rect 455288 290436 455294 290448
rect 533338 290436 533344 290448
rect 533396 290436 533402 290488
rect 383194 289756 383200 289808
rect 383252 289796 383258 289808
rect 516318 289796 516324 289808
rect 383252 289768 516324 289796
rect 383252 289756 383258 289768
rect 516318 289756 516324 289768
rect 516376 289756 516382 289808
rect 386230 289688 386236 289740
rect 386288 289728 386294 289740
rect 520458 289728 520464 289740
rect 386288 289700 520464 289728
rect 386288 289688 386294 289700
rect 520458 289688 520464 289700
rect 520516 289688 520522 289740
rect 380434 289620 380440 289672
rect 380492 289660 380498 289672
rect 515030 289660 515036 289672
rect 380492 289632 515036 289660
rect 380492 289620 380498 289632
rect 515030 289620 515036 289632
rect 515088 289620 515094 289672
rect 383286 289552 383292 289604
rect 383344 289592 383350 289604
rect 519078 289592 519084 289604
rect 383344 289564 519084 289592
rect 383344 289552 383350 289564
rect 519078 289552 519084 289564
rect 519136 289552 519142 289604
rect 380342 289484 380348 289536
rect 380400 289524 380406 289536
rect 516502 289524 516508 289536
rect 380400 289496 516508 289524
rect 380400 289484 380406 289496
rect 516502 289484 516508 289496
rect 516560 289484 516566 289536
rect 383010 289416 383016 289468
rect 383068 289456 383074 289468
rect 519354 289456 519360 289468
rect 383068 289428 519360 289456
rect 383068 289416 383074 289428
rect 519354 289416 519360 289428
rect 519412 289416 519418 289468
rect 383102 289348 383108 289400
rect 383160 289388 383166 289400
rect 520550 289388 520556 289400
rect 383160 289360 520556 289388
rect 383160 289348 383166 289360
rect 520550 289348 520556 289360
rect 520608 289348 520614 289400
rect 378870 289280 378876 289332
rect 378928 289320 378934 289332
rect 517606 289320 517612 289332
rect 378928 289292 517612 289320
rect 378928 289280 378934 289292
rect 517606 289280 517612 289292
rect 517664 289280 517670 289332
rect 363782 289212 363788 289264
rect 363840 289252 363846 289264
rect 507302 289252 507308 289264
rect 363840 289224 507308 289252
rect 363840 289212 363846 289224
rect 507302 289212 507308 289224
rect 507360 289212 507366 289264
rect 373350 289144 373356 289196
rect 373408 289184 373414 289196
rect 520366 289184 520372 289196
rect 373408 289156 520372 289184
rect 373408 289144 373414 289156
rect 520366 289144 520372 289156
rect 520424 289144 520430 289196
rect 370590 289076 370596 289128
rect 370648 289116 370654 289128
rect 523034 289116 523040 289128
rect 370648 289088 523040 289116
rect 370648 289076 370654 289088
rect 523034 289076 523040 289088
rect 523092 289076 523098 289128
rect 385954 289008 385960 289060
rect 386012 289048 386018 289060
rect 507486 289048 507492 289060
rect 386012 289020 507492 289048
rect 386012 289008 386018 289020
rect 507486 289008 507492 289020
rect 507544 289008 507550 289060
rect 386046 288940 386052 288992
rect 386104 288980 386110 288992
rect 507210 288980 507216 288992
rect 386104 288952 507216 288980
rect 386104 288940 386110 288952
rect 507210 288940 507216 288952
rect 507268 288940 507274 288992
rect 446582 288872 446588 288924
rect 446640 288912 446646 288924
rect 464338 288912 464344 288924
rect 446640 288884 464344 288912
rect 446640 288872 446646 288884
rect 464338 288872 464344 288884
rect 464396 288872 464402 288924
rect 473998 288804 474004 288856
rect 474056 288844 474062 288856
rect 478138 288844 478144 288856
rect 474056 288816 478144 288844
rect 474056 288804 474062 288816
rect 478138 288804 478144 288816
rect 478196 288804 478202 288856
rect 465994 287648 466000 287700
rect 466052 287688 466058 287700
rect 569218 287688 569224 287700
rect 466052 287660 569224 287688
rect 466052 287648 466058 287660
rect 569218 287648 569224 287660
rect 569276 287648 569282 287700
rect 452010 286764 452016 286816
rect 452068 286804 452074 286816
rect 487522 286804 487528 286816
rect 452068 286776 487528 286804
rect 452068 286764 452074 286776
rect 487522 286764 487528 286776
rect 487580 286764 487586 286816
rect 456794 286696 456800 286748
rect 456852 286736 456858 286748
rect 504910 286736 504916 286748
rect 456852 286708 504916 286736
rect 456852 286696 456858 286708
rect 504910 286696 504916 286708
rect 504968 286696 504974 286748
rect 439682 286628 439688 286680
rect 439740 286668 439746 286680
rect 446582 286668 446588 286680
rect 439740 286640 446588 286668
rect 439740 286628 439746 286640
rect 446582 286628 446588 286640
rect 446640 286628 446646 286680
rect 475654 286628 475660 286680
rect 475712 286668 475718 286680
rect 571978 286668 571984 286680
rect 475712 286640 571984 286668
rect 475712 286628 475718 286640
rect 571978 286628 571984 286640
rect 572036 286628 572042 286680
rect 377490 286560 377496 286612
rect 377548 286600 377554 286612
rect 507118 286600 507124 286612
rect 377548 286572 507124 286600
rect 377548 286560 377554 286572
rect 507118 286560 507124 286572
rect 507176 286560 507182 286612
rect 384942 286492 384948 286544
rect 385000 286532 385006 286544
rect 521838 286532 521844 286544
rect 385000 286504 521844 286532
rect 385000 286492 385006 286504
rect 521838 286492 521844 286504
rect 521896 286492 521902 286544
rect 374822 286424 374828 286476
rect 374880 286464 374886 286476
rect 521654 286464 521660 286476
rect 374880 286436 521660 286464
rect 374880 286424 374886 286436
rect 521654 286424 521660 286436
rect 521712 286424 521718 286476
rect 372062 286356 372068 286408
rect 372120 286396 372126 286408
rect 521746 286396 521752 286408
rect 372120 286368 521752 286396
rect 372120 286356 372126 286368
rect 521746 286356 521752 286368
rect 521804 286356 521810 286408
rect 369394 286288 369400 286340
rect 369452 286328 369458 286340
rect 523126 286328 523132 286340
rect 369452 286300 523132 286328
rect 369452 286288 369458 286300
rect 523126 286288 523132 286300
rect 523184 286288 523190 286340
rect 460382 285676 460388 285728
rect 460440 285716 460446 285728
rect 462682 285716 462688 285728
rect 460440 285688 462688 285716
rect 460440 285676 460446 285688
rect 462682 285676 462688 285688
rect 462740 285676 462746 285728
rect 453574 285064 453580 285116
rect 453632 285104 453638 285116
rect 493870 285104 493876 285116
rect 453632 285076 493876 285104
rect 453632 285064 453638 285076
rect 493870 285064 493876 285076
rect 493928 285064 493934 285116
rect 464890 284996 464896 285048
rect 464948 285036 464954 285048
rect 547138 285036 547144 285048
rect 464948 285008 547144 285036
rect 464948 284996 464954 285008
rect 547138 284996 547144 285008
rect 547196 284996 547202 285048
rect 363690 284928 363696 284980
rect 363748 284968 363754 284980
rect 474826 284968 474832 284980
rect 363748 284940 474832 284968
rect 363748 284928 363754 284940
rect 474826 284928 474832 284940
rect 474884 284928 474890 284980
rect 486142 284928 486148 284980
rect 486200 284968 486206 284980
rect 531314 284968 531320 284980
rect 486200 284940 531320 284968
rect 486200 284928 486206 284940
rect 531314 284928 531320 284940
rect 531372 284928 531378 284980
rect 452286 283704 452292 283756
rect 452344 283744 452350 283756
rect 493042 283744 493048 283756
rect 452344 283716 493048 283744
rect 452344 283704 452350 283716
rect 493042 283704 493048 283716
rect 493100 283704 493106 283756
rect 501874 283704 501880 283756
rect 501932 283744 501938 283756
rect 539226 283744 539232 283756
rect 501932 283716 539232 283744
rect 501932 283704 501938 283716
rect 539226 283704 539232 283716
rect 539284 283704 539290 283756
rect 449894 283636 449900 283688
rect 449952 283676 449958 283688
rect 504634 283676 504640 283688
rect 449952 283648 504640 283676
rect 449952 283636 449958 283648
rect 504634 283636 504640 283648
rect 504692 283636 504698 283688
rect 446398 283568 446404 283620
rect 446456 283608 446462 283620
rect 457622 283608 457628 283620
rect 446456 283580 457628 283608
rect 446456 283568 446462 283580
rect 457622 283568 457628 283580
rect 457680 283568 457686 283620
rect 476482 283568 476488 283620
rect 476540 283608 476546 283620
rect 566458 283608 566464 283620
rect 476540 283580 566464 283608
rect 476540 283568 476546 283580
rect 566458 283568 566464 283580
rect 566516 283568 566522 283620
rect 361758 282820 361764 282872
rect 361816 282860 361822 282872
rect 431218 282860 431224 282872
rect 361816 282832 431224 282860
rect 361816 282820 361822 282832
rect 431218 282820 431224 282832
rect 431276 282820 431282 282872
rect 471238 282208 471244 282260
rect 471296 282248 471302 282260
rect 473998 282248 474004 282260
rect 471296 282220 474004 282248
rect 471296 282208 471302 282220
rect 473998 282208 474004 282220
rect 474056 282208 474062 282260
rect 456242 282140 456248 282192
rect 456300 282180 456306 282192
rect 492490 282180 492496 282192
rect 456300 282152 492496 282180
rect 456300 282140 456306 282152
rect 492490 282140 492496 282152
rect 492548 282140 492554 282192
rect 459278 280780 459284 280832
rect 459336 280820 459342 280832
rect 491386 280820 491392 280832
rect 459336 280792 491392 280820
rect 459336 280780 459342 280792
rect 491386 280780 491392 280792
rect 491444 280780 491450 280832
rect 459186 279420 459192 279472
rect 459244 279460 459250 279472
rect 490558 279460 490564 279472
rect 459244 279432 490564 279460
rect 459244 279420 459250 279432
rect 490558 279420 490564 279432
rect 490616 279420 490622 279472
rect 452378 277992 452384 278044
rect 452436 278032 452442 278044
rect 493318 278032 493324 278044
rect 452436 278004 493324 278032
rect 452436 277992 452442 278004
rect 493318 277992 493324 278004
rect 493376 277992 493382 278044
rect 498838 277992 498844 278044
rect 498896 278032 498902 278044
rect 541526 278032 541532 278044
rect 498896 278004 541532 278032
rect 498896 277992 498902 278004
rect 541526 277992 541532 278004
rect 541584 277992 541590 278044
rect 460290 276768 460296 276820
rect 460348 276808 460354 276820
rect 489454 276808 489460 276820
rect 460348 276780 489460 276808
rect 460348 276768 460354 276780
rect 489454 276768 489460 276780
rect 489512 276768 489518 276820
rect 498010 276768 498016 276820
rect 498068 276808 498074 276820
rect 539870 276808 539876 276820
rect 498068 276780 539876 276808
rect 498068 276768 498074 276780
rect 539870 276768 539876 276780
rect 539928 276768 539934 276820
rect 457714 276700 457720 276752
rect 457772 276740 457778 276752
rect 491662 276740 491668 276752
rect 457772 276712 491668 276740
rect 457772 276700 457778 276712
rect 491662 276700 491668 276712
rect 491720 276700 491726 276752
rect 496906 276700 496912 276752
rect 496964 276740 496970 276752
rect 539778 276740 539784 276752
rect 496964 276712 539784 276740
rect 496964 276700 496970 276712
rect 539778 276700 539784 276712
rect 539836 276700 539842 276752
rect 359642 276632 359648 276684
rect 359700 276672 359706 276684
rect 511994 276672 512000 276684
rect 359700 276644 512000 276672
rect 359700 276632 359706 276644
rect 511994 276632 512000 276644
rect 512052 276632 512058 276684
rect 497734 275408 497740 275460
rect 497792 275448 497798 275460
rect 541434 275448 541440 275460
rect 497792 275420 541440 275448
rect 497792 275408 497798 275420
rect 541434 275408 541440 275420
rect 541492 275408 541498 275460
rect 457622 275340 457628 275392
rect 457680 275380 457686 275392
rect 490834 275380 490840 275392
rect 457680 275352 490840 275380
rect 457680 275340 457686 275352
rect 490834 275340 490840 275352
rect 490892 275340 490898 275392
rect 495250 275340 495256 275392
rect 495308 275380 495314 275392
rect 541250 275380 541256 275392
rect 495308 275352 541256 275380
rect 495308 275340 495314 275352
rect 541250 275340 541256 275352
rect 541308 275340 541314 275392
rect 453482 275272 453488 275324
rect 453540 275312 453546 275324
rect 488074 275312 488080 275324
rect 453540 275284 488080 275312
rect 453540 275272 453546 275284
rect 488074 275272 488080 275284
rect 488132 275272 488138 275324
rect 495802 275272 495808 275324
rect 495860 275312 495866 275324
rect 542814 275312 542820 275324
rect 495860 275284 542820 275312
rect 495860 275272 495866 275284
rect 542814 275272 542820 275284
rect 542872 275272 542878 275324
rect 456978 274660 456984 274712
rect 457036 274700 457042 274712
rect 460382 274700 460388 274712
rect 457036 274672 460388 274700
rect 457036 274660 457042 274672
rect 460382 274660 460388 274672
rect 460440 274660 460446 274712
rect 499114 274048 499120 274100
rect 499172 274088 499178 274100
rect 540054 274088 540060 274100
rect 499172 274060 540060 274088
rect 499172 274048 499178 274060
rect 540054 274048 540060 274060
rect 540112 274048 540118 274100
rect 456150 273980 456156 274032
rect 456208 274020 456214 274032
rect 490374 274020 490380 274032
rect 456208 273992 490380 274020
rect 456208 273980 456214 273992
rect 490374 273980 490380 273992
rect 490432 273980 490438 274032
rect 497458 273980 497464 274032
rect 497516 274020 497522 274032
rect 541342 274020 541348 274032
rect 497516 273992 541348 274020
rect 497516 273980 497522 273992
rect 541342 273980 541348 273992
rect 541400 273980 541406 274032
rect 453666 273912 453672 273964
rect 453724 273952 453730 273964
rect 493594 273952 493600 273964
rect 453724 273924 493600 273952
rect 453724 273912 453730 273924
rect 493594 273912 493600 273924
rect 493652 273912 493658 273964
rect 495526 273912 495532 273964
rect 495584 273952 495590 273964
rect 542630 273952 542636 273964
rect 495584 273924 542636 273952
rect 495584 273912 495590 273924
rect 542630 273912 542636 273924
rect 542688 273912 542694 273964
rect 476758 273164 476764 273216
rect 476816 273204 476822 273216
rect 580166 273204 580172 273216
rect 476816 273176 580172 273204
rect 476816 273164 476822 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 456058 272552 456064 272604
rect 456116 272592 456122 272604
rect 489730 272592 489736 272604
rect 456116 272564 489736 272592
rect 456116 272552 456122 272564
rect 489730 272552 489736 272564
rect 489788 272552 489794 272604
rect 498562 272552 498568 272604
rect 498620 272592 498626 272604
rect 539962 272592 539968 272604
rect 498620 272564 539968 272592
rect 498620 272552 498626 272564
rect 539962 272552 539968 272564
rect 540020 272552 540026 272604
rect 454954 272484 454960 272536
rect 455012 272524 455018 272536
rect 491938 272524 491944 272536
rect 455012 272496 491944 272524
rect 455012 272484 455018 272496
rect 491938 272484 491944 272496
rect 491996 272484 492002 272536
rect 496354 272484 496360 272536
rect 496412 272524 496418 272536
rect 542906 272524 542912 272536
rect 496412 272496 542912 272524
rect 496412 272484 496418 272496
rect 542906 272484 542912 272496
rect 542964 272484 542970 272536
rect 361758 271804 361764 271856
rect 361816 271844 361822 271856
rect 439590 271844 439596 271856
rect 361816 271816 439596 271844
rect 361816 271804 361822 271816
rect 439590 271804 439596 271816
rect 439648 271804 439654 271856
rect 501322 271396 501328 271448
rect 501380 271436 501386 271448
rect 540330 271436 540336 271448
rect 501380 271408 540336 271436
rect 501380 271396 501386 271408
rect 540330 271396 540336 271408
rect 540388 271396 540394 271448
rect 456334 271328 456340 271380
rect 456392 271368 456398 271380
rect 491110 271368 491116 271380
rect 456392 271340 491116 271368
rect 456392 271328 456398 271340
rect 491110 271328 491116 271340
rect 491168 271328 491174 271380
rect 494974 271328 494980 271380
rect 495032 271368 495038 271380
rect 539686 271368 539692 271380
rect 495032 271340 539692 271368
rect 495032 271328 495038 271340
rect 539686 271328 539692 271340
rect 539744 271328 539750 271380
rect 436830 271260 436836 271312
rect 436888 271300 436894 271312
rect 439682 271300 439688 271312
rect 436888 271272 439688 271300
rect 436888 271260 436894 271272
rect 439682 271260 439688 271272
rect 439740 271260 439746 271312
rect 454862 271260 454868 271312
rect 454920 271300 454926 271312
rect 504358 271300 504364 271312
rect 454920 271272 504364 271300
rect 454920 271260 454926 271272
rect 504358 271260 504364 271272
rect 504416 271260 504422 271312
rect 450722 271192 450728 271244
rect 450780 271232 450786 271244
rect 503530 271232 503536 271244
rect 450780 271204 503536 271232
rect 450780 271192 450786 271204
rect 503530 271192 503536 271204
rect 503588 271192 503594 271244
rect 466270 271124 466276 271176
rect 466328 271164 466334 271176
rect 580258 271164 580264 271176
rect 466328 271136 580264 271164
rect 466328 271124 466334 271136
rect 580258 271124 580264 271136
rect 580316 271124 580322 271176
rect 500494 270036 500500 270088
rect 500552 270076 500558 270088
rect 540238 270076 540244 270088
rect 500552 270048 540244 270076
rect 500552 270036 500558 270048
rect 540238 270036 540244 270048
rect 540296 270036 540302 270088
rect 455046 269968 455052 270020
rect 455104 270008 455110 270020
rect 486694 270008 486700 270020
rect 455104 269980 486700 270008
rect 455104 269968 455110 269980
rect 486694 269968 486700 269980
rect 486752 269968 486758 270020
rect 499942 269968 499948 270020
rect 500000 270008 500006 270020
rect 543090 270008 543096 270020
rect 500000 269980 543096 270008
rect 500000 269968 500006 269980
rect 543090 269968 543096 269980
rect 543148 269968 543154 270020
rect 450814 269900 450820 269952
rect 450872 269940 450878 269952
rect 503254 269940 503260 269952
rect 450872 269912 503260 269940
rect 450872 269900 450878 269912
rect 503254 269900 503260 269912
rect 503312 269900 503318 269952
rect 465442 269832 465448 269884
rect 465500 269872 465506 269884
rect 554038 269872 554044 269884
rect 465500 269844 554044 269872
rect 465500 269832 465506 269844
rect 554038 269832 554044 269844
rect 554096 269832 554102 269884
rect 445662 269764 445668 269816
rect 445720 269804 445726 269816
rect 510614 269804 510620 269816
rect 445720 269776 510620 269804
rect 445720 269764 445726 269776
rect 510614 269764 510620 269776
rect 510672 269764 510678 269816
rect 442994 269288 443000 269340
rect 443052 269328 443058 269340
rect 446398 269328 446404 269340
rect 443052 269300 446404 269328
rect 443052 269288 443058 269300
rect 446398 269288 446404 269300
rect 446456 269288 446462 269340
rect 447778 268540 447784 268592
rect 447836 268580 447842 268592
rect 456978 268580 456984 268592
rect 447836 268552 456984 268580
rect 447836 268540 447842 268552
rect 456978 268540 456984 268552
rect 457036 268540 457042 268592
rect 453758 268472 453764 268524
rect 453816 268512 453822 268524
rect 472618 268512 472624 268524
rect 453816 268484 472624 268512
rect 453816 268472 453822 268484
rect 472618 268472 472624 268484
rect 472676 268472 472682 268524
rect 500218 268472 500224 268524
rect 500276 268512 500282 268524
rect 540146 268512 540152 268524
rect 500276 268484 540152 268512
rect 500276 268472 500282 268484
rect 540146 268472 540152 268484
rect 540204 268472 540210 268524
rect 450078 268404 450084 268456
rect 450136 268444 450142 268456
rect 471238 268444 471244 268456
rect 450136 268416 471244 268444
rect 450136 268404 450142 268416
rect 471238 268404 471244 268416
rect 471296 268404 471302 268456
rect 499390 268404 499396 268456
rect 499448 268444 499454 268456
rect 542998 268444 543004 268456
rect 499448 268416 543004 268444
rect 499448 268404 499454 268416
rect 542998 268404 543004 268416
rect 543056 268404 543062 268456
rect 452194 268336 452200 268388
rect 452252 268376 452258 268388
rect 487798 268376 487804 268388
rect 452252 268348 487804 268376
rect 452252 268336 452258 268348
rect 487798 268336 487804 268348
rect 487856 268336 487862 268388
rect 494698 268336 494704 268388
rect 494756 268376 494762 268388
rect 542538 268376 542544 268388
rect 494756 268348 542544 268376
rect 494756 268336 494762 268348
rect 542538 268336 542544 268348
rect 542596 268336 542602 268388
rect 449618 263508 449624 263560
rect 449676 263548 449682 263560
rect 456978 263548 456984 263560
rect 449676 263520 456984 263548
rect 449676 263508 449682 263520
rect 456978 263508 456984 263520
rect 457036 263508 457042 263560
rect 440234 262760 440240 262812
rect 440292 262800 440298 262812
rect 442994 262800 443000 262812
rect 440292 262772 443000 262800
rect 440292 262760 440298 262772
rect 442994 262760 443000 262772
rect 443052 262760 443058 262812
rect 445018 262760 445024 262812
rect 445076 262800 445082 262812
rect 450078 262800 450084 262812
rect 445076 262772 450084 262800
rect 445076 262760 445082 262772
rect 450078 262760 450084 262772
rect 450136 262760 450142 262812
rect 361758 260788 361764 260840
rect 361816 260828 361822 260840
rect 440970 260828 440976 260840
rect 361816 260800 440976 260828
rect 361816 260788 361822 260800
rect 440970 260788 440976 260800
rect 441028 260788 441034 260840
rect 431954 260312 431960 260364
rect 432012 260352 432018 260364
rect 440234 260352 440240 260364
rect 432012 260324 440240 260352
rect 432012 260312 432018 260324
rect 440234 260312 440240 260324
rect 440292 260312 440298 260364
rect 429930 254872 429936 254924
rect 429988 254912 429994 254924
rect 431954 254912 431960 254924
rect 429988 254884 431960 254912
rect 429988 254872 429994 254884
rect 431954 254872 431960 254884
rect 432012 254872 432018 254924
rect 3786 253920 3792 253972
rect 3844 253960 3850 253972
rect 4982 253960 4988 253972
rect 3844 253932 4988 253960
rect 3844 253920 3850 253932
rect 4982 253920 4988 253932
rect 5040 253920 5046 253972
rect 442442 252424 442448 252476
rect 442500 252464 442506 252476
rect 447778 252464 447784 252476
rect 442500 252436 447784 252464
rect 442500 252424 442506 252436
rect 447778 252424 447784 252436
rect 447836 252424 447842 252476
rect 361758 249704 361764 249756
rect 361816 249744 361822 249756
rect 435450 249744 435456 249756
rect 361816 249716 435456 249744
rect 361816 249704 361822 249716
rect 435450 249704 435456 249716
rect 435508 249704 435514 249756
rect 442350 249704 442356 249756
rect 442408 249744 442414 249756
rect 445018 249744 445024 249756
rect 442408 249716 445024 249744
rect 442408 249704 442414 249716
rect 445018 249704 445024 249716
rect 445076 249704 445082 249756
rect 449710 249024 449716 249076
rect 449768 249064 449774 249076
rect 458082 249064 458088 249076
rect 449768 249036 458088 249064
rect 449768 249024 449774 249036
rect 458082 249024 458088 249036
rect 458140 249024 458146 249076
rect 573358 245556 573364 245608
rect 573416 245596 573422 245608
rect 580166 245596 580172 245608
rect 573416 245568 580172 245596
rect 573416 245556 573422 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 439590 244944 439596 244996
rect 439648 244984 439654 244996
rect 442442 244984 442448 244996
rect 439648 244956 442448 244984
rect 439648 244944 439654 244956
rect 442442 244944 442448 244956
rect 442500 244944 442506 244996
rect 3878 241408 3884 241460
rect 3936 241448 3942 241460
rect 5074 241448 5080 241460
rect 3936 241420 5080 241448
rect 3936 241408 3942 241420
rect 5074 241408 5080 241420
rect 5132 241408 5138 241460
rect 361758 238688 361764 238740
rect 361816 238728 361822 238740
rect 442258 238728 442264 238740
rect 361816 238700 442264 238728
rect 361816 238688 361822 238700
rect 442258 238688 442264 238700
rect 442316 238688 442322 238740
rect 419442 233860 419448 233912
rect 419500 233900 419506 233912
rect 456702 233900 456708 233912
rect 419500 233872 456708 233900
rect 419500 233860 419506 233872
rect 456702 233860 456708 233872
rect 456760 233860 456766 233912
rect 566458 233180 566464 233232
rect 566516 233220 566522 233232
rect 579982 233220 579988 233232
rect 566516 233192 579988 233220
rect 566516 233180 566522 233192
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 448238 232568 448244 232620
rect 448296 232608 448302 232620
rect 454034 232608 454040 232620
rect 448296 232580 454040 232608
rect 448296 232568 448302 232580
rect 454034 232568 454040 232580
rect 454092 232568 454098 232620
rect 428458 232500 428464 232552
rect 428516 232540 428522 232552
rect 453758 232540 453764 232552
rect 428516 232512 453764 232540
rect 428516 232500 428522 232512
rect 453758 232500 453764 232512
rect 453816 232500 453822 232552
rect 433978 230936 433984 230988
rect 434036 230976 434042 230988
rect 439590 230976 439596 230988
rect 434036 230948 439596 230976
rect 434036 230936 434042 230948
rect 439590 230936 439596 230948
rect 439648 230936 439654 230988
rect 424318 227740 424324 227792
rect 424376 227780 424382 227792
rect 429930 227780 429936 227792
rect 424376 227752 429936 227780
rect 424376 227740 424382 227752
rect 429930 227740 429936 227752
rect 429988 227740 429994 227792
rect 361758 227672 361764 227724
rect 361816 227712 361822 227724
rect 443638 227712 443644 227724
rect 361816 227684 443644 227712
rect 361816 227672 361822 227684
rect 443638 227672 443644 227684
rect 443696 227672 443702 227724
rect 416038 221416 416044 221468
rect 416096 221456 416102 221468
rect 454034 221456 454040 221468
rect 416096 221428 454040 221456
rect 416096 221416 416102 221428
rect 454034 221416 454040 221428
rect 454092 221456 454098 221468
rect 457898 221456 457904 221468
rect 454092 221428 457904 221456
rect 454092 221416 454098 221428
rect 457898 221416 457904 221428
rect 457956 221416 457962 221468
rect 569218 219376 569224 219428
rect 569276 219416 569282 219428
rect 580166 219416 580172 219428
rect 569276 219388 580172 219416
rect 569276 219376 569282 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 427814 217540 427820 217592
rect 427872 217580 427878 217592
rect 433978 217580 433984 217592
rect 427872 217552 433984 217580
rect 427872 217540 427878 217552
rect 433978 217540 433984 217552
rect 434036 217540 434042 217592
rect 423030 216656 423036 216708
rect 423088 216696 423094 216708
rect 428458 216696 428464 216708
rect 423088 216668 428464 216696
rect 423088 216656 423094 216668
rect 428458 216656 428464 216668
rect 428516 216656 428522 216708
rect 361666 216316 361672 216368
rect 361724 216356 361730 216368
rect 364058 216356 364064 216368
rect 361724 216328 364064 216356
rect 361724 216316 361730 216328
rect 364058 216316 364064 216328
rect 364116 216316 364122 216368
rect 3970 214752 3976 214804
rect 4028 214792 4034 214804
rect 5166 214792 5172 214804
rect 4028 214764 5172 214792
rect 4028 214752 4034 214764
rect 5166 214752 5172 214764
rect 5224 214752 5230 214804
rect 422938 213120 422944 213172
rect 422996 213160 423002 213172
rect 427814 213160 427820 213172
rect 422996 213132 427820 213160
rect 422996 213120 423002 213132
rect 427814 213120 427820 213132
rect 427872 213120 427878 213172
rect 434254 212984 434260 213036
rect 434312 213024 434318 213036
rect 436830 213024 436836 213036
rect 434312 212996 436836 213024
rect 434312 212984 434318 212996
rect 436830 212984 436836 212996
rect 436888 212984 436894 213036
rect 406378 211760 406384 211812
rect 406436 211800 406442 211812
rect 423030 211800 423036 211812
rect 406436 211772 423036 211800
rect 406436 211760 406442 211772
rect 423030 211760 423036 211772
rect 423088 211760 423094 211812
rect 420178 209788 420184 209840
rect 420236 209828 420242 209840
rect 424318 209828 424324 209840
rect 420236 209800 424324 209828
rect 420236 209788 420242 209800
rect 424318 209788 424324 209800
rect 424376 209788 424382 209840
rect 428458 209788 428464 209840
rect 428516 209828 428522 209840
rect 434254 209828 434260 209840
rect 428516 209800 434260 209828
rect 428516 209788 428522 209800
rect 434254 209788 434260 209800
rect 434312 209788 434318 209840
rect 570598 206932 570604 206984
rect 570656 206972 570662 206984
rect 579798 206972 579804 206984
rect 570656 206944 579804 206972
rect 570656 206932 570662 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 411254 206252 411260 206304
rect 411312 206292 411318 206304
rect 448330 206292 448336 206304
rect 411312 206264 448336 206292
rect 411312 206252 411318 206264
rect 448330 206252 448336 206264
rect 448388 206292 448394 206304
rect 456702 206292 456708 206304
rect 448388 206264 456708 206292
rect 448388 206252 448394 206264
rect 456702 206252 456708 206264
rect 456760 206252 456766 206304
rect 361758 205572 361764 205624
rect 361816 205612 361822 205624
rect 439498 205612 439504 205624
rect 361816 205584 439504 205612
rect 361816 205572 361822 205584
rect 439498 205572 439504 205584
rect 439556 205572 439562 205624
rect 433242 203532 433248 203584
rect 433300 203572 433306 203584
rect 442350 203572 442356 203584
rect 433300 203544 442356 203572
rect 433300 203532 433306 203544
rect 442350 203532 442356 203544
rect 442408 203532 442414 203584
rect 419534 201492 419540 201544
rect 419592 201532 419598 201544
rect 422938 201532 422944 201544
rect 419592 201504 422944 201532
rect 419592 201492 419598 201504
rect 422938 201492 422944 201504
rect 422996 201492 423002 201544
rect 417418 200744 417424 200796
rect 417476 200784 417482 200796
rect 433242 200784 433248 200796
rect 417476 200756 433248 200784
rect 417476 200744 417482 200756
rect 433242 200744 433248 200756
rect 433300 200744 433306 200796
rect 459462 200744 459468 200796
rect 459520 200784 459526 200796
rect 485774 200784 485780 200796
rect 459520 200756 485780 200784
rect 459520 200744 459526 200756
rect 485774 200744 485780 200756
rect 485832 200744 485838 200796
rect 458082 200132 458088 200184
rect 458140 200172 458146 200184
rect 462958 200172 462964 200184
rect 458140 200144 462964 200172
rect 458140 200132 458146 200144
rect 462958 200132 462964 200144
rect 463016 200132 463022 200184
rect 459370 199384 459376 199436
rect 459428 199424 459434 199436
rect 481634 199424 481640 199436
rect 459428 199396 481640 199424
rect 459428 199384 459434 199396
rect 481634 199384 481640 199396
rect 481692 199384 481698 199436
rect 398098 196664 398104 196716
rect 398156 196704 398162 196716
rect 419534 196704 419540 196716
rect 398156 196676 419540 196704
rect 398156 196664 398162 196676
rect 419534 196664 419540 196676
rect 419592 196664 419598 196716
rect 367738 196596 367744 196648
rect 367796 196636 367802 196648
rect 406378 196636 406384 196648
rect 367796 196608 406384 196636
rect 367796 196596 367802 196608
rect 406378 196596 406384 196608
rect 406436 196596 406442 196648
rect 448422 196596 448428 196648
rect 448480 196636 448486 196648
rect 461578 196636 461584 196648
rect 448480 196608 461584 196636
rect 448480 196596 448486 196608
rect 461578 196596 461584 196608
rect 461636 196596 461642 196648
rect 449986 195236 449992 195288
rect 450044 195276 450050 195288
rect 528554 195276 528560 195288
rect 450044 195248 528560 195276
rect 450044 195236 450050 195248
rect 528554 195236 528560 195248
rect 528612 195236 528618 195288
rect 416130 194692 416136 194744
rect 416188 194732 416194 194744
rect 420178 194732 420184 194744
rect 416188 194704 420184 194732
rect 416188 194692 416194 194704
rect 420178 194692 420184 194704
rect 420236 194692 420242 194744
rect 361758 194488 361764 194540
rect 361816 194528 361822 194540
rect 429838 194528 429844 194540
rect 361816 194500 429844 194528
rect 361816 194488 361822 194500
rect 429838 194488 429844 194500
rect 429896 194488 429902 194540
rect 392578 193808 392584 193860
rect 392636 193848 392642 193860
rect 398098 193848 398104 193860
rect 392636 193820 398104 193848
rect 392636 193808 392642 193820
rect 398098 193808 398104 193820
rect 398156 193808 398162 193860
rect 548518 193128 548524 193180
rect 548576 193168 548582 193180
rect 580166 193168 580172 193180
rect 548576 193140 580172 193168
rect 548576 193128 548582 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 404998 189728 405004 189780
rect 405056 189768 405062 189780
rect 416130 189768 416136 189780
rect 405056 189740 416136 189768
rect 405056 189728 405062 189740
rect 416130 189728 416136 189740
rect 416188 189728 416194 189780
rect 361758 183472 361764 183524
rect 361816 183512 361822 183524
rect 436738 183512 436744 183524
rect 361816 183484 436744 183512
rect 361816 183472 361822 183484
rect 436738 183472 436744 183484
rect 436796 183472 436802 183524
rect 389910 182112 389916 182164
rect 389968 182152 389974 182164
rect 392578 182152 392584 182164
rect 389968 182124 392584 182152
rect 389968 182112 389974 182124
rect 392578 182112 392584 182124
rect 392636 182112 392642 182164
rect 361574 180072 361580 180124
rect 361632 180112 361638 180124
rect 417418 180112 417424 180124
rect 361632 180084 417424 180112
rect 361632 180072 361638 180084
rect 417418 180072 417424 180084
rect 417476 180072 417482 180124
rect 537478 179324 537484 179376
rect 537536 179364 537542 179376
rect 580166 179364 580172 179376
rect 537536 179336 580172 179364
rect 537536 179324 537542 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 401594 172524 401600 172576
rect 401652 172564 401658 172576
rect 404998 172564 405004 172576
rect 401652 172536 405004 172564
rect 401652 172524 401658 172536
rect 404998 172524 405004 172536
rect 405056 172524 405062 172576
rect 361758 171776 361764 171828
rect 361816 171816 361822 171828
rect 440878 171816 440884 171828
rect 361816 171788 440884 171816
rect 361816 171776 361822 171788
rect 440878 171776 440884 171788
rect 440936 171816 440942 171828
rect 524414 171816 524420 171828
rect 440936 171788 524420 171816
rect 440936 171776 440942 171788
rect 524414 171776 524420 171788
rect 524472 171776 524478 171828
rect 397454 169736 397460 169788
rect 397512 169776 397518 169788
rect 401594 169776 401600 169788
rect 397512 169748 401600 169776
rect 397512 169736 397518 169748
rect 401594 169736 401600 169748
rect 401652 169736 401658 169788
rect 362678 167628 362684 167680
rect 362736 167668 362742 167680
rect 389910 167668 389916 167680
rect 362736 167640 389916 167668
rect 362736 167628 362742 167640
rect 389910 167628 389916 167640
rect 389968 167628 389974 167680
rect 533338 166948 533344 167000
rect 533396 166988 533402 167000
rect 580166 166988 580172 167000
rect 533396 166960 580172 166988
rect 533396 166948 533402 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 390554 164840 390560 164892
rect 390612 164880 390618 164892
rect 397454 164880 397460 164892
rect 390612 164852 397460 164880
rect 390612 164840 390618 164852
rect 397454 164840 397460 164852
rect 397512 164840 397518 164892
rect 414750 163888 414756 163940
rect 414808 163928 414814 163940
rect 416038 163928 416044 163940
rect 414808 163900 416044 163928
rect 414808 163888 414814 163900
rect 416038 163888 416044 163900
rect 416096 163888 416102 163940
rect 434898 162800 434904 162852
rect 434956 162840 434962 162852
rect 435358 162840 435364 162852
rect 434956 162812 435364 162840
rect 434956 162800 434962 162812
rect 435358 162800 435364 162812
rect 435416 162800 435422 162852
rect 365714 162188 365720 162240
rect 365772 162228 365778 162240
rect 390554 162228 390560 162240
rect 365772 162200 390560 162228
rect 365772 162188 365778 162200
rect 390554 162188 390560 162200
rect 390612 162188 390618 162240
rect 389818 162120 389824 162172
rect 389876 162160 389882 162172
rect 444926 162160 444932 162172
rect 389876 162132 444932 162160
rect 389876 162120 389882 162132
rect 444926 162120 444932 162132
rect 444984 162120 444990 162172
rect 425054 161848 425060 161900
rect 425112 161888 425118 161900
rect 426342 161888 426348 161900
rect 425112 161860 426348 161888
rect 425112 161848 425118 161860
rect 426342 161848 426348 161860
rect 426400 161888 426406 161900
rect 496814 161888 496820 161900
rect 426400 161860 496820 161888
rect 426400 161848 426406 161860
rect 496814 161848 496820 161860
rect 496872 161848 496878 161900
rect 428642 161780 428648 161832
rect 428700 161820 428706 161832
rect 500954 161820 500960 161832
rect 428700 161792 500960 161820
rect 428700 161780 428706 161792
rect 500954 161780 500960 161792
rect 501012 161780 501018 161832
rect 421742 161712 421748 161764
rect 421800 161752 421806 161764
rect 494054 161752 494060 161764
rect 421800 161724 494060 161752
rect 421800 161712 421806 161724
rect 494054 161712 494060 161724
rect 494112 161712 494118 161764
rect 410518 161644 410524 161696
rect 410576 161684 410582 161696
rect 425054 161684 425060 161696
rect 410576 161656 425060 161684
rect 410576 161644 410582 161656
rect 425054 161644 425060 161656
rect 425112 161644 425118 161696
rect 431862 161644 431868 161696
rect 431920 161684 431926 161696
rect 505094 161684 505100 161696
rect 431920 161656 505100 161684
rect 431920 161644 431926 161656
rect 505094 161644 505100 161656
rect 505152 161644 505158 161696
rect 407758 161576 407764 161628
rect 407816 161616 407822 161628
rect 434898 161616 434904 161628
rect 407816 161588 434904 161616
rect 407816 161576 407822 161588
rect 434898 161576 434904 161588
rect 434956 161576 434962 161628
rect 438762 161576 438768 161628
rect 438820 161616 438826 161628
rect 513374 161616 513380 161628
rect 438820 161588 513380 161616
rect 438820 161576 438826 161588
rect 513374 161576 513380 161588
rect 513432 161576 513438 161628
rect 403618 161508 403624 161560
rect 403676 161548 403682 161560
rect 438780 161548 438808 161576
rect 442902 161548 442908 161560
rect 403676 161520 438808 161548
rect 441586 161520 442908 161548
rect 403676 161508 403682 161520
rect 441586 161492 441614 161520
rect 442902 161508 442908 161520
rect 442960 161548 442966 161560
rect 517514 161548 517520 161560
rect 442960 161520 517520 161548
rect 442960 161508 442966 161520
rect 517514 161508 517520 161520
rect 517572 161508 517578 161560
rect 362586 161440 362592 161492
rect 362644 161480 362650 161492
rect 441586 161480 441620 161492
rect 362644 161452 441620 161480
rect 362644 161440 362650 161452
rect 441614 161440 441620 161452
rect 441672 161440 441678 161492
rect 444926 161440 444932 161492
rect 444984 161480 444990 161492
rect 445662 161480 445668 161492
rect 444984 161452 445668 161480
rect 444984 161440 444990 161452
rect 445662 161440 445668 161452
rect 445720 161480 445726 161492
rect 532694 161480 532700 161492
rect 445720 161452 532700 161480
rect 445720 161440 445726 161452
rect 532694 161440 532700 161452
rect 532752 161440 532758 161492
rect 361758 161372 361764 161424
rect 361816 161412 361822 161424
rect 444190 161412 444196 161424
rect 361816 161384 444196 161412
rect 361816 161372 361822 161384
rect 444190 161372 444196 161384
rect 444248 161372 444254 161424
rect 359826 160692 359832 160744
rect 359884 160732 359890 160744
rect 367738 160732 367744 160744
rect 359884 160704 367744 160732
rect 359884 160692 359890 160704
rect 367738 160692 367744 160704
rect 367796 160692 367802 160744
rect 420914 160692 420920 160744
rect 420972 160732 420978 160744
rect 428458 160732 428464 160744
rect 420972 160704 428464 160732
rect 420972 160692 420978 160704
rect 428458 160692 428464 160704
rect 428516 160692 428522 160744
rect 444190 160692 444196 160744
rect 444248 160732 444254 160744
rect 521654 160732 521660 160744
rect 444248 160704 521660 160732
rect 444248 160692 444254 160704
rect 521654 160692 521660 160704
rect 521712 160692 521718 160744
rect 410610 160352 410616 160404
rect 410668 160392 410674 160404
rect 427998 160392 428004 160404
rect 410668 160364 428004 160392
rect 410668 160352 410674 160364
rect 427998 160352 428004 160364
rect 428056 160352 428062 160404
rect 406378 160284 406384 160336
rect 406436 160324 406442 160336
rect 431310 160324 431316 160336
rect 406436 160296 431316 160324
rect 406436 160284 406442 160296
rect 431310 160284 431316 160296
rect 431368 160284 431374 160336
rect 386322 160216 386328 160268
rect 386380 160256 386386 160268
rect 414750 160256 414756 160268
rect 386380 160228 414756 160256
rect 386380 160216 386386 160228
rect 414750 160216 414756 160228
rect 414808 160216 414814 160268
rect 381354 160148 381360 160200
rect 381412 160188 381418 160200
rect 421374 160188 421380 160200
rect 381412 160160 421380 160188
rect 381412 160148 381418 160160
rect 421374 160148 421380 160160
rect 421432 160188 421438 160200
rect 421742 160188 421748 160200
rect 421432 160160 421748 160188
rect 421432 160148 421438 160160
rect 421742 160148 421748 160160
rect 421800 160148 421806 160200
rect 434898 160148 434904 160200
rect 434956 160188 434962 160200
rect 435266 160188 435272 160200
rect 434956 160160 435272 160188
rect 434956 160148 434962 160160
rect 435266 160148 435272 160160
rect 435324 160188 435330 160200
rect 450906 160188 450912 160200
rect 435324 160160 450912 160188
rect 435324 160148 435330 160160
rect 450906 160148 450912 160160
rect 450964 160148 450970 160200
rect 359734 160080 359740 160132
rect 359792 160120 359798 160132
rect 362678 160120 362684 160132
rect 359792 160092 362684 160120
rect 359792 160080 359798 160092
rect 362678 160080 362684 160092
rect 362736 160080 362742 160132
rect 383378 160080 383384 160132
rect 383436 160120 383442 160132
rect 418384 160120 418390 160132
rect 383436 160092 418390 160120
rect 383436 160080 383442 160092
rect 418384 160080 418390 160092
rect 418442 160120 418448 160132
rect 419442 160120 419448 160132
rect 418442 160092 419448 160120
rect 418442 160080 418448 160092
rect 419442 160080 419448 160092
rect 419500 160120 419506 160132
rect 461670 160120 461676 160132
rect 419500 160092 461676 160120
rect 419500 160080 419506 160092
rect 461670 160080 461676 160092
rect 461728 160080 461734 160132
rect 420914 159508 420920 159520
rect 412606 159480 420920 159508
rect 407390 159400 407396 159452
rect 407448 159440 407454 159452
rect 412606 159440 412634 159480
rect 420914 159468 420920 159480
rect 420972 159468 420978 159520
rect 407448 159412 412634 159440
rect 407448 159400 407454 159412
rect 449802 159332 449808 159384
rect 449860 159372 449866 159384
rect 536834 159372 536840 159384
rect 449860 159344 536840 159372
rect 449860 159332 449866 159344
rect 536834 159332 536840 159344
rect 536892 159332 536898 159384
rect 452562 158380 452568 158432
rect 452620 158420 452626 158432
rect 455046 158420 455052 158432
rect 452620 158392 455052 158420
rect 452620 158380 452626 158392
rect 455046 158380 455052 158392
rect 455104 158380 455110 158432
rect 452378 157292 452384 157344
rect 452436 157332 452442 157344
rect 453390 157332 453396 157344
rect 452436 157304 453396 157332
rect 452436 157292 452442 157304
rect 453390 157292 453396 157304
rect 453448 157292 453454 157344
rect 405642 156068 405648 156120
rect 405700 156108 405706 156120
rect 407390 156108 407396 156120
rect 405700 156080 407396 156108
rect 405700 156068 405706 156080
rect 407390 156068 407396 156080
rect 407448 156068 407454 156120
rect 359918 155864 359924 155916
rect 359976 155904 359982 155916
rect 365714 155904 365720 155916
rect 359976 155876 365720 155904
rect 359976 155864 359982 155876
rect 365714 155864 365720 155876
rect 365772 155864 365778 155916
rect 452378 155796 452384 155848
rect 452436 155836 452442 155848
rect 453574 155836 453580 155848
rect 452436 155808 453580 155836
rect 452436 155796 452442 155808
rect 453574 155796 453580 155808
rect 453632 155796 453638 155848
rect 452378 154300 452384 154352
rect 452436 154340 452442 154352
rect 453666 154340 453672 154352
rect 452436 154312 453672 154340
rect 452436 154300 452442 154312
rect 453666 154300 453672 154312
rect 453724 154300 453730 154352
rect 402330 153212 402336 153264
rect 402388 153252 402394 153264
rect 405642 153252 405648 153264
rect 402388 153224 405648 153252
rect 402388 153212 402394 153224
rect 405642 153212 405648 153224
rect 405700 153212 405706 153264
rect 536098 153144 536104 153196
rect 536156 153184 536162 153196
rect 580166 153184 580172 153196
rect 536156 153156 580172 153184
rect 536156 153144 536162 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 452562 148996 452568 149048
rect 452620 149036 452626 149048
rect 456242 149036 456248 149048
rect 452620 149008 456248 149036
rect 452620 148996 452626 149008
rect 456242 148996 456248 149008
rect 456300 148996 456306 149048
rect 399478 147636 399484 147688
rect 399536 147676 399542 147688
rect 402330 147676 402336 147688
rect 399536 147648 402336 147676
rect 399536 147636 399542 147648
rect 402330 147636 402336 147648
rect 402388 147636 402394 147688
rect 452562 147500 452568 147552
rect 452620 147540 452626 147552
rect 459002 147540 459008 147552
rect 452620 147512 459008 147540
rect 452620 147500 452626 147512
rect 459002 147500 459008 147512
rect 459060 147500 459066 147552
rect 452562 146140 452568 146192
rect 452620 146180 452626 146192
rect 454954 146180 454960 146192
rect 452620 146152 454960 146180
rect 452620 146140 452626 146152
rect 454954 146140 454960 146152
rect 455012 146140 455018 146192
rect 452562 144780 452568 144832
rect 452620 144820 452626 144832
rect 457714 144820 457720 144832
rect 452620 144792 457720 144820
rect 452620 144780 452626 144792
rect 457714 144780 457720 144792
rect 457772 144780 457778 144832
rect 452562 143420 452568 143472
rect 452620 143460 452626 143472
rect 459278 143460 459284 143472
rect 452620 143432 459284 143460
rect 452620 143420 452626 143432
rect 459278 143420 459284 143432
rect 459336 143420 459342 143472
rect 461670 142876 461676 142928
rect 461728 142916 461734 142928
rect 489914 142916 489920 142928
rect 461728 142888 489920 142916
rect 461728 142876 461734 142888
rect 489914 142876 489920 142888
rect 489972 142876 489978 142928
rect 450906 142808 450912 142860
rect 450964 142848 450970 142860
rect 509602 142848 509608 142860
rect 450964 142820 509608 142848
rect 450964 142808 450970 142820
rect 509602 142808 509608 142820
rect 509660 142808 509666 142860
rect 452562 142060 452568 142112
rect 452620 142100 452626 142112
rect 456334 142100 456340 142112
rect 452620 142072 456340 142100
rect 452620 142060 452626 142072
rect 456334 142060 456340 142072
rect 456392 142060 456398 142112
rect 464338 140768 464344 140820
rect 464396 140808 464402 140820
rect 481634 140808 481640 140820
rect 464396 140780 481640 140808
rect 464396 140768 464402 140780
rect 481634 140768 481640 140780
rect 481692 140768 481698 140820
rect 452562 140700 452568 140752
rect 452620 140740 452626 140752
rect 457622 140740 457628 140752
rect 452620 140712 457628 140740
rect 452620 140700 452626 140712
rect 457622 140700 457628 140712
rect 457680 140700 457686 140752
rect 388438 140020 388444 140072
rect 388496 140060 388502 140072
rect 399478 140060 399484 140072
rect 388496 140032 399484 140060
rect 388496 140020 388502 140032
rect 399478 140020 399484 140032
rect 399536 140020 399542 140072
rect 361758 139340 361764 139392
rect 361816 139380 361822 139392
rect 403618 139380 403624 139392
rect 361816 139352 403624 139380
rect 361816 139340 361822 139352
rect 403618 139340 403624 139352
rect 403676 139340 403682 139392
rect 452562 139340 452568 139392
rect 452620 139380 452626 139392
rect 459186 139380 459192 139392
rect 452620 139352 459192 139380
rect 452620 139340 452626 139352
rect 459186 139340 459192 139352
rect 459244 139340 459250 139392
rect 554038 139340 554044 139392
rect 554096 139380 554102 139392
rect 580166 139380 580172 139392
rect 554096 139352 580172 139380
rect 554096 139340 554102 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 452562 137844 452568 137896
rect 452620 137884 452626 137896
rect 456150 137884 456156 137896
rect 452620 137856 456156 137884
rect 452620 137844 452626 137856
rect 456150 137844 456156 137856
rect 456208 137844 456214 137896
rect 451550 136484 451556 136536
rect 451608 136524 451614 136536
rect 457530 136524 457536 136536
rect 451608 136496 457536 136524
rect 451608 136484 451614 136496
rect 457530 136484 457536 136496
rect 457588 136484 457594 136536
rect 452562 135124 452568 135176
rect 452620 135164 452626 135176
rect 456058 135164 456064 135176
rect 452620 135136 456064 135164
rect 452620 135124 452626 135136
rect 456058 135124 456064 135136
rect 456116 135124 456122 135176
rect 452562 133764 452568 133816
rect 452620 133804 452626 133816
rect 460290 133804 460296 133816
rect 452620 133776 460296 133804
rect 452620 133764 452626 133776
rect 460290 133764 460296 133776
rect 460348 133764 460354 133816
rect 452562 132404 452568 132456
rect 452620 132444 452626 132456
rect 457438 132444 457444 132456
rect 452620 132416 457444 132444
rect 452620 132404 452626 132416
rect 457438 132404 457444 132416
rect 457496 132404 457502 132456
rect 452562 131044 452568 131096
rect 452620 131084 452626 131096
rect 459094 131084 459100 131096
rect 452620 131056 459100 131084
rect 452620 131044 452626 131056
rect 459094 131044 459100 131056
rect 459152 131044 459158 131096
rect 452562 129684 452568 129736
rect 452620 129724 452626 129736
rect 458910 129724 458916 129736
rect 452620 129696 458916 129724
rect 452620 129684 452626 129696
rect 458910 129684 458916 129696
rect 458968 129684 458974 129736
rect 361758 128256 361764 128308
rect 361816 128296 361822 128308
rect 407758 128296 407764 128308
rect 361816 128268 407764 128296
rect 361816 128256 361822 128268
rect 407758 128256 407764 128268
rect 407816 128256 407822 128308
rect 452286 128256 452292 128308
rect 452344 128296 452350 128308
rect 453298 128296 453304 128308
rect 452344 128268 453304 128296
rect 452344 128256 452350 128268
rect 453298 128256 453304 128268
rect 453356 128256 453362 128308
rect 452378 126896 452384 126948
rect 452436 126936 452442 126948
rect 453482 126936 453488 126948
rect 452436 126908 453488 126936
rect 452436 126896 452442 126908
rect 453482 126896 453488 126908
rect 453540 126896 453546 126948
rect 574738 126896 574744 126948
rect 574796 126936 574802 126948
rect 580166 126936 580172 126948
rect 574796 126908 580172 126936
rect 574796 126896 574802 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 362586 124856 362592 124908
rect 362644 124896 362650 124908
rect 388438 124896 388444 124908
rect 362644 124868 388444 124896
rect 362644 124856 362650 124868
rect 388438 124856 388444 124868
rect 388496 124856 388502 124908
rect 451918 122136 451924 122188
rect 451976 122176 451982 122188
rect 458818 122176 458824 122188
rect 451976 122148 458824 122176
rect 451976 122136 451982 122148
rect 458818 122136 458824 122148
rect 458876 122136 458882 122188
rect 361758 117240 361764 117292
rect 361816 117280 361822 117292
rect 406378 117280 406384 117292
rect 361816 117252 406384 117280
rect 361816 117240 361822 117252
rect 406378 117240 406384 117252
rect 406436 117240 406442 117292
rect 571978 113092 571984 113144
rect 572036 113132 572042 113144
rect 579798 113132 579804 113144
rect 572036 113104 579804 113132
rect 572036 113092 572042 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 445294 107312 445300 107364
rect 445352 107352 445358 107364
rect 454862 107352 454868 107364
rect 445352 107324 454868 107352
rect 445352 107312 445358 107324
rect 454862 107312 454868 107324
rect 454920 107312 454926 107364
rect 439130 107244 439136 107296
rect 439188 107284 439194 107296
rect 450630 107284 450636 107296
rect 439188 107256 450636 107284
rect 439188 107244 439194 107256
rect 450630 107244 450636 107256
rect 450688 107244 450694 107296
rect 432966 107176 432972 107228
rect 433024 107216 433030 107228
rect 450538 107216 450544 107228
rect 433024 107188 450544 107216
rect 433024 107176 433030 107188
rect 450538 107176 450544 107188
rect 450596 107176 450602 107228
rect 426802 107108 426808 107160
rect 426860 107148 426866 107160
rect 450722 107148 450728 107160
rect 426860 107120 450728 107148
rect 426860 107108 426866 107120
rect 450722 107108 450728 107120
rect 450780 107108 450786 107160
rect 420638 107040 420644 107092
rect 420696 107080 420702 107092
rect 450814 107080 450820 107092
rect 420696 107052 450820 107080
rect 420696 107040 420702 107052
rect 450814 107040 450820 107052
rect 450872 107040 450878 107092
rect 414474 106972 414480 107024
rect 414532 107012 414538 107024
rect 454678 107012 454684 107024
rect 414532 106984 454684 107012
rect 414532 106972 414538 106984
rect 454678 106972 454684 106984
rect 454736 106972 454742 107024
rect 402146 106904 402152 106956
rect 402204 106944 402210 106956
rect 454770 106944 454776 106956
rect 402204 106916 454776 106944
rect 402204 106904 402210 106916
rect 454770 106904 454776 106916
rect 454828 106904 454834 106956
rect 367738 106292 367744 106344
rect 367796 106332 367802 106344
rect 389818 106332 389824 106344
rect 367796 106304 389824 106332
rect 367796 106292 367802 106304
rect 389818 106292 389824 106304
rect 389876 106292 389882 106344
rect 361758 106224 361764 106276
rect 361816 106264 361822 106276
rect 410610 106264 410616 106276
rect 361816 106236 410616 106264
rect 361816 106224 361822 106236
rect 410610 106224 410616 106236
rect 410668 106224 410674 106276
rect 362678 105544 362684 105596
rect 362736 105584 362742 105596
rect 410518 105584 410524 105596
rect 362736 105556 410524 105584
rect 362736 105544 362742 105556
rect 410518 105544 410524 105556
rect 410576 105544 410582 105596
rect 551278 100648 551284 100700
rect 551336 100688 551342 100700
rect 580166 100688 580172 100700
rect 551336 100660 580172 100688
rect 551336 100648 551342 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 3694 98608 3700 98660
rect 3752 98648 3758 98660
rect 19978 98648 19984 98660
rect 3752 98620 19984 98648
rect 3752 98608 3758 98620
rect 19978 98608 19984 98620
rect 20036 98608 20042 98660
rect 4890 97996 4896 98048
rect 4948 98036 4954 98048
rect 4948 98008 6914 98036
rect 4948 97996 4954 98008
rect 6886 97968 6914 98008
rect 8938 97968 8944 97980
rect 6886 97940 8944 97968
rect 8938 97928 8944 97940
rect 8996 97928 9002 97980
rect 576118 86912 576124 86964
rect 576176 86952 576182 86964
rect 580166 86952 580172 86964
rect 576176 86924 580172 86952
rect 576176 86912 576182 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 3142 84192 3148 84244
rect 3200 84232 3206 84244
rect 20898 84232 20904 84244
rect 3200 84204 20904 84232
rect 3200 84192 3206 84204
rect 20898 84192 20904 84204
rect 20956 84192 20962 84244
rect 361758 84124 361764 84176
rect 361816 84164 361822 84176
rect 381354 84164 381360 84176
rect 361816 84136 381360 84164
rect 361816 84124 361822 84136
rect 381354 84124 381360 84136
rect 381412 84124 381418 84176
rect 361758 73108 361764 73160
rect 361816 73148 361822 73160
rect 383378 73148 383384 73160
rect 361816 73120 383384 73148
rect 361816 73108 361822 73120
rect 383378 73108 383384 73120
rect 383436 73108 383442 73160
rect 544378 73108 544384 73160
rect 544436 73148 544442 73160
rect 580166 73148 580172 73160
rect 544436 73120 580172 73148
rect 544436 73108 544442 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 4982 71204 4988 71256
rect 5040 71244 5046 71256
rect 6178 71244 6184 71256
rect 5040 71216 6184 71244
rect 5040 71204 5046 71216
rect 6178 71204 6184 71216
rect 6236 71204 6242 71256
rect 3142 70388 3148 70440
rect 3200 70428 3206 70440
rect 20070 70428 20076 70440
rect 3200 70400 20076 70428
rect 3200 70388 3206 70400
rect 20070 70388 20076 70400
rect 20128 70388 20134 70440
rect 8938 67532 8944 67584
rect 8996 67572 9002 67584
rect 10962 67572 10968 67584
rect 8996 67544 10968 67572
rect 8996 67532 9002 67544
rect 10962 67532 10968 67544
rect 11020 67532 11026 67584
rect 462498 67532 462504 67584
rect 462556 67572 462562 67584
rect 464338 67572 464344 67584
rect 462556 67544 464344 67572
rect 462556 67532 462562 67544
rect 464338 67532 464344 67544
rect 464396 67532 464402 67584
rect 4798 66852 4804 66904
rect 4856 66892 4862 66904
rect 7282 66892 7288 66904
rect 4856 66864 7288 66892
rect 4856 66852 4862 66864
rect 7282 66852 7288 66864
rect 7340 66852 7346 66904
rect 7282 63656 7288 63708
rect 7340 63696 7346 63708
rect 9674 63696 9680 63708
rect 7340 63668 9680 63696
rect 7340 63656 7346 63668
rect 9674 63656 9680 63668
rect 9732 63656 9738 63708
rect 361758 62024 361764 62076
rect 361816 62064 361822 62076
rect 386322 62064 386328 62076
rect 361816 62036 386328 62064
rect 361816 62024 361822 62036
rect 386322 62024 386328 62036
rect 386380 62024 386386 62076
rect 5074 60664 5080 60716
rect 5132 60704 5138 60716
rect 5994 60704 6000 60716
rect 5132 60676 6000 60704
rect 5132 60664 5138 60676
rect 5994 60664 6000 60676
rect 6052 60664 6058 60716
rect 547138 60664 547144 60716
rect 547196 60704 547202 60716
rect 580166 60704 580172 60716
rect 547196 60676 580172 60704
rect 547196 60664 547202 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 11054 59372 11060 59424
rect 11112 59412 11118 59424
rect 11112 59384 12480 59412
rect 11112 59372 11118 59384
rect 12452 59344 12480 59384
rect 13814 59344 13820 59356
rect 12452 59316 13820 59344
rect 13814 59304 13820 59316
rect 13872 59304 13878 59356
rect 5994 58624 6000 58676
rect 6052 58664 6058 58676
rect 11698 58664 11704 58676
rect 6052 58636 11704 58664
rect 6052 58624 6058 58636
rect 11698 58624 11704 58636
rect 11756 58624 11762 58676
rect 5166 57196 5172 57248
rect 5224 57236 5230 57248
rect 8202 57236 8208 57248
rect 5224 57208 8208 57236
rect 5224 57196 5230 57208
rect 8202 57196 8208 57208
rect 8260 57196 8266 57248
rect 13814 56516 13820 56568
rect 13872 56556 13878 56568
rect 16482 56556 16488 56568
rect 13872 56528 16488 56556
rect 13872 56516 13878 56528
rect 16482 56516 16488 56528
rect 16540 56516 16546 56568
rect 9674 55224 9680 55276
rect 9732 55264 9738 55276
rect 9732 55236 11100 55264
rect 9732 55224 9738 55236
rect 11072 55196 11100 55236
rect 13722 55196 13728 55208
rect 11072 55168 13728 55196
rect 13722 55156 13728 55168
rect 13780 55156 13786 55208
rect 6178 53796 6184 53848
rect 6236 53836 6242 53848
rect 6236 53808 6914 53836
rect 6236 53796 6242 53808
rect 6886 53768 6914 53808
rect 8386 53768 8392 53780
rect 6886 53740 8392 53768
rect 8386 53728 8392 53740
rect 8444 53728 8450 53780
rect 11698 53388 11704 53440
rect 11756 53428 11762 53440
rect 13722 53428 13728 53440
rect 11756 53400 13728 53428
rect 11756 53388 11762 53400
rect 13722 53388 13728 53400
rect 13780 53388 13786 53440
rect 8202 52436 8208 52488
rect 8260 52476 8266 52488
rect 8260 52448 8340 52476
rect 8260 52436 8266 52448
rect 8312 52408 8340 52448
rect 11054 52408 11060 52420
rect 8312 52380 11060 52408
rect 11054 52368 11060 52380
rect 11112 52368 11118 52420
rect 8386 51688 8392 51740
rect 8444 51728 8450 51740
rect 19242 51728 19248 51740
rect 8444 51700 19248 51728
rect 8444 51688 8450 51700
rect 19242 51688 19248 51700
rect 19300 51688 19306 51740
rect 13722 51076 13728 51128
rect 13780 51116 13786 51128
rect 13780 51088 13952 51116
rect 13780 51076 13786 51088
rect 13924 51048 13952 51088
rect 361758 51076 361764 51128
rect 361816 51116 361822 51128
rect 384206 51116 384212 51128
rect 361816 51088 384212 51116
rect 361816 51076 361822 51088
rect 384206 51076 384212 51088
rect 384264 51076 384270 51128
rect 540606 51076 540612 51128
rect 540664 51116 540670 51128
rect 543734 51116 543740 51128
rect 540664 51088 543740 51116
rect 540664 51076 540670 51088
rect 543734 51076 543740 51088
rect 543792 51076 543798 51128
rect 17862 51048 17868 51060
rect 13924 51020 17868 51048
rect 17862 51008 17868 51020
rect 17920 51008 17926 51060
rect 13814 50940 13820 50992
rect 13872 50980 13878 50992
rect 18598 50980 18604 50992
rect 13872 50952 18604 50980
rect 13872 50940 13878 50952
rect 18598 50940 18604 50952
rect 18656 50940 18662 50992
rect 16574 50124 16580 50176
rect 16632 50164 16638 50176
rect 19334 50164 19340 50176
rect 16632 50136 19340 50164
rect 16632 50124 16638 50136
rect 19334 50124 19340 50136
rect 19392 50124 19398 50176
rect 11054 49716 11060 49768
rect 11112 49756 11118 49768
rect 11112 49728 16574 49756
rect 11112 49716 11118 49728
rect 16546 49688 16574 49728
rect 18230 49688 18236 49700
rect 16546 49660 18236 49688
rect 18230 49648 18236 49660
rect 18288 49648 18294 49700
rect 18598 48288 18604 48340
rect 18656 48328 18662 48340
rect 18656 48300 19380 48328
rect 18656 48288 18662 48300
rect 19352 48260 19380 48300
rect 20898 48260 20904 48272
rect 19352 48232 20904 48260
rect 20898 48220 20904 48232
rect 20956 48220 20962 48272
rect 17862 48152 17868 48204
rect 17920 48192 17926 48204
rect 20714 48192 20720 48204
rect 17920 48164 20720 48192
rect 17920 48152 17926 48164
rect 20714 48152 20720 48164
rect 20772 48152 20778 48204
rect 18230 47880 18236 47932
rect 18288 47920 18294 47932
rect 20806 47920 20812 47932
rect 18288 47892 20812 47920
rect 18288 47880 18294 47892
rect 20806 47880 20812 47892
rect 20864 47880 20870 47932
rect 19334 46996 19340 47048
rect 19392 47036 19398 47048
rect 21266 47036 21272 47048
rect 19392 47008 21272 47036
rect 19392 46996 19398 47008
rect 21266 46996 21272 47008
rect 21324 46996 21330 47048
rect 3510 46860 3516 46912
rect 3568 46900 3574 46912
rect 386138 46900 386144 46912
rect 3568 46872 386144 46900
rect 3568 46860 3574 46872
rect 386138 46860 386144 46872
rect 386196 46860 386202 46912
rect 3694 46792 3700 46844
rect 3752 46832 3758 46844
rect 385862 46832 385868 46844
rect 3752 46804 385868 46832
rect 3752 46792 3758 46804
rect 385862 46792 385868 46804
rect 385920 46792 385926 46844
rect 3234 46724 3240 46776
rect 3292 46764 3298 46776
rect 384574 46764 384580 46776
rect 3292 46736 384580 46764
rect 3292 46724 3298 46736
rect 384574 46724 384580 46736
rect 384632 46724 384638 46776
rect 3326 46656 3332 46708
rect 3384 46696 3390 46708
rect 381630 46696 381636 46708
rect 3384 46668 381636 46696
rect 3384 46656 3390 46668
rect 381630 46656 381636 46668
rect 381688 46656 381694 46708
rect 3970 46588 3976 46640
rect 4028 46628 4034 46640
rect 381722 46628 381728 46640
rect 4028 46600 381728 46628
rect 4028 46588 4034 46600
rect 381722 46588 381728 46600
rect 381780 46588 381786 46640
rect 3878 46520 3884 46572
rect 3936 46560 3942 46572
rect 381446 46560 381452 46572
rect 3936 46532 381452 46560
rect 3936 46520 3942 46532
rect 381446 46520 381452 46532
rect 381504 46520 381510 46572
rect 3602 46452 3608 46504
rect 3660 46492 3666 46504
rect 379422 46492 379428 46504
rect 3660 46464 379428 46492
rect 3660 46452 3666 46464
rect 379422 46452 379428 46464
rect 379480 46452 379486 46504
rect 3786 46384 3792 46436
rect 3844 46424 3850 46436
rect 378686 46424 378692 46436
rect 3844 46396 378692 46424
rect 3844 46384 3850 46396
rect 378686 46384 378692 46396
rect 378744 46384 378750 46436
rect 20070 46316 20076 46368
rect 20128 46356 20134 46368
rect 384390 46356 384396 46368
rect 20128 46328 384396 46356
rect 20128 46316 20134 46328
rect 384390 46316 384396 46328
rect 384448 46316 384454 46368
rect 19978 46248 19984 46300
rect 20036 46288 20042 46300
rect 376662 46288 376668 46300
rect 20036 46260 376668 46288
rect 20036 46248 20042 46260
rect 376662 46248 376668 46260
rect 376720 46248 376726 46300
rect 20806 46180 20812 46232
rect 20864 46220 20870 46232
rect 359918 46220 359924 46232
rect 20864 46192 359924 46220
rect 20864 46180 20870 46192
rect 359918 46180 359924 46192
rect 359976 46180 359982 46232
rect 20714 46112 20720 46164
rect 20772 46152 20778 46164
rect 359826 46152 359832 46164
rect 20772 46124 359832 46152
rect 20772 46112 20778 46124
rect 359826 46112 359832 46124
rect 359884 46112 359890 46164
rect 21266 46044 21272 46096
rect 21324 46084 21330 46096
rect 359734 46084 359740 46096
rect 21324 46056 359740 46084
rect 21324 46044 21330 46056
rect 359734 46044 359740 46056
rect 359792 46044 359798 46096
rect 358170 45772 358176 45824
rect 358228 45812 358234 45824
rect 362586 45812 362592 45824
rect 358228 45784 362592 45812
rect 358228 45772 358234 45784
rect 362586 45772 362592 45784
rect 362644 45772 362650 45824
rect 4062 45568 4068 45620
rect 4120 45568 4126 45620
rect 4080 45540 4108 45568
rect 381538 45540 381544 45552
rect 4080 45512 381544 45540
rect 381538 45500 381544 45512
rect 381596 45500 381602 45552
rect 3510 45432 3516 45484
rect 3568 45472 3574 45484
rect 376570 45472 376576 45484
rect 3568 45444 376576 45472
rect 3568 45432 3574 45444
rect 376570 45432 376576 45444
rect 376628 45432 376634 45484
rect 20898 45364 20904 45416
rect 20956 45404 20962 45416
rect 358170 45404 358176 45416
rect 20956 45376 358176 45404
rect 20956 45364 20962 45376
rect 358170 45364 358176 45376
rect 358228 45364 358234 45416
rect 71774 45296 71780 45348
rect 71832 45336 71838 45348
rect 378962 45336 378968 45348
rect 71832 45308 378968 45336
rect 71832 45296 71838 45308
rect 378962 45296 378968 45308
rect 379020 45296 379026 45348
rect 69014 45228 69020 45280
rect 69072 45268 69078 45280
rect 379238 45268 379244 45280
rect 69072 45240 379244 45268
rect 69072 45228 69078 45240
rect 379238 45228 379244 45240
rect 379296 45228 379302 45280
rect 64874 45160 64880 45212
rect 64932 45200 64938 45212
rect 379330 45200 379336 45212
rect 64932 45172 379336 45200
rect 64932 45160 64938 45172
rect 379330 45160 379336 45172
rect 379388 45160 379394 45212
rect 60734 45092 60740 45144
rect 60792 45132 60798 45144
rect 382090 45132 382096 45144
rect 60792 45104 382096 45132
rect 60792 45092 60798 45104
rect 382090 45092 382096 45104
rect 382148 45092 382154 45144
rect 57974 45024 57980 45076
rect 58032 45064 58038 45076
rect 381998 45064 382004 45076
rect 58032 45036 382004 45064
rect 58032 45024 58038 45036
rect 381998 45024 382004 45036
rect 382056 45024 382062 45076
rect 53834 44956 53840 45008
rect 53892 44996 53898 45008
rect 381906 44996 381912 45008
rect 53892 44968 381912 44996
rect 53892 44956 53898 44968
rect 381906 44956 381912 44968
rect 381964 44956 381970 45008
rect 51074 44888 51080 44940
rect 51132 44928 51138 44940
rect 382182 44928 382188 44940
rect 51132 44900 382188 44928
rect 51132 44888 51138 44900
rect 382182 44888 382188 44900
rect 382240 44888 382246 44940
rect 6914 44820 6920 44872
rect 6972 44860 6978 44872
rect 384666 44860 384672 44872
rect 6972 44832 384672 44860
rect 6972 44820 6978 44832
rect 384666 44820 384672 44832
rect 384724 44820 384730 44872
rect 75914 44752 75920 44804
rect 75972 44792 75978 44804
rect 379146 44792 379152 44804
rect 75972 44764 379152 44792
rect 75972 44752 75978 44764
rect 379146 44752 379152 44764
rect 379204 44752 379210 44804
rect 78674 44684 78680 44736
rect 78732 44724 78738 44736
rect 379054 44724 379060 44736
rect 78732 44696 379060 44724
rect 78732 44684 78738 44696
rect 379054 44684 379060 44696
rect 379112 44684 379118 44736
rect 85574 44616 85580 44668
rect 85632 44656 85638 44668
rect 376478 44656 376484 44668
rect 85632 44628 376484 44656
rect 85632 44616 85638 44628
rect 376478 44616 376484 44628
rect 376536 44616 376542 44668
rect 114554 42712 114560 42764
rect 114612 42752 114618 42764
rect 370958 42752 370964 42764
rect 114612 42724 370964 42752
rect 114612 42712 114618 42724
rect 370958 42712 370964 42724
rect 371016 42712 371022 42764
rect 110414 42644 110420 42696
rect 110472 42684 110478 42696
rect 370866 42684 370872 42696
rect 110472 42656 370872 42684
rect 110472 42644 110478 42656
rect 370866 42644 370872 42656
rect 370924 42644 370930 42696
rect 107654 42576 107660 42628
rect 107712 42616 107718 42628
rect 373258 42616 373264 42628
rect 107712 42588 373264 42616
rect 107712 42576 107718 42588
rect 373258 42576 373264 42588
rect 373316 42576 373322 42628
rect 103514 42508 103520 42560
rect 103572 42548 103578 42560
rect 373442 42548 373448 42560
rect 103572 42520 373448 42548
rect 103572 42508 103578 42520
rect 373442 42508 373448 42520
rect 373500 42508 373506 42560
rect 100754 42440 100760 42492
rect 100812 42480 100818 42492
rect 373534 42480 373540 42492
rect 100812 42452 373540 42480
rect 100812 42440 100818 42452
rect 373534 42440 373540 42452
rect 373592 42440 373598 42492
rect 96614 42372 96620 42424
rect 96672 42412 96678 42424
rect 373626 42412 373632 42424
rect 96672 42384 373632 42412
rect 96672 42372 96678 42384
rect 373626 42372 373632 42384
rect 373684 42372 373690 42424
rect 93854 42304 93860 42356
rect 93912 42344 93918 42356
rect 376386 42344 376392 42356
rect 93912 42316 376392 42344
rect 93912 42304 93918 42316
rect 376386 42304 376392 42316
rect 376444 42304 376450 42356
rect 89714 42236 89720 42288
rect 89772 42276 89778 42288
rect 376294 42276 376300 42288
rect 89772 42248 376300 42276
rect 89772 42236 89778 42248
rect 376294 42236 376300 42248
rect 376352 42236 376358 42288
rect 82814 42168 82820 42220
rect 82872 42208 82878 42220
rect 376202 42208 376208 42220
rect 82872 42180 376208 42208
rect 82872 42168 82878 42180
rect 376202 42168 376208 42180
rect 376260 42168 376266 42220
rect 20714 42100 20720 42152
rect 20772 42140 20778 42152
rect 368290 42140 368296 42152
rect 20772 42112 368296 42140
rect 20772 42100 20778 42112
rect 368290 42100 368296 42112
rect 368348 42100 368354 42152
rect 11054 42032 11060 42084
rect 11112 42072 11118 42084
rect 376110 42072 376116 42084
rect 11112 42044 376116 42072
rect 11112 42032 11118 42044
rect 376110 42032 376116 42044
rect 376168 42032 376174 42084
rect 118694 41964 118700 42016
rect 118752 42004 118758 42016
rect 371050 42004 371056 42016
rect 118752 41976 371056 42004
rect 118752 41964 118758 41976
rect 371050 41964 371056 41976
rect 371108 41964 371114 42016
rect 121454 41896 121460 41948
rect 121512 41936 121518 41948
rect 370774 41936 370780 41948
rect 121512 41908 370780 41936
rect 121512 41896 121518 41908
rect 370774 41896 370780 41908
rect 370832 41896 370838 41948
rect 461578 41352 461584 41404
rect 461636 41392 461642 41404
rect 536834 41392 536840 41404
rect 461636 41364 536840 41392
rect 461636 41352 461642 41364
rect 536834 41352 536840 41364
rect 536892 41352 536898 41404
rect 77294 39992 77300 40044
rect 77352 40032 77358 40044
rect 361298 40032 361304 40044
rect 77352 40004 361304 40032
rect 77352 39992 77358 40004
rect 361298 39992 361304 40004
rect 361356 39992 361362 40044
rect 73154 39924 73160 39976
rect 73212 39964 73218 39976
rect 362494 39964 362500 39976
rect 73212 39936 362500 39964
rect 73212 39924 73218 39936
rect 362494 39924 362500 39936
rect 362552 39924 362558 39976
rect 69106 39856 69112 39908
rect 69164 39896 69170 39908
rect 362402 39896 362408 39908
rect 69164 39868 362408 39896
rect 69164 39856 69170 39868
rect 362402 39856 362408 39868
rect 362460 39856 362466 39908
rect 66254 39788 66260 39840
rect 66312 39828 66318 39840
rect 362218 39828 362224 39840
rect 66312 39800 362224 39828
rect 66312 39788 66318 39800
rect 362218 39788 362224 39800
rect 362276 39788 362282 39840
rect 62114 39720 62120 39772
rect 62172 39760 62178 39772
rect 362310 39760 362316 39772
rect 62172 39732 362316 39760
rect 62172 39720 62178 39732
rect 362310 39720 362316 39732
rect 362368 39720 362374 39772
rect 59354 39652 59360 39704
rect 59412 39692 59418 39704
rect 365254 39692 365260 39704
rect 59412 39664 365260 39692
rect 59412 39652 59418 39664
rect 365254 39652 365260 39664
rect 365312 39652 365318 39704
rect 44174 39584 44180 39636
rect 44232 39624 44238 39636
rect 365530 39624 365536 39636
rect 44232 39596 365536 39624
rect 44232 39584 44238 39596
rect 365530 39584 365536 39596
rect 365588 39584 365594 39636
rect 40034 39516 40040 39568
rect 40092 39556 40098 39568
rect 365438 39556 365444 39568
rect 40092 39528 365444 39556
rect 40092 39516 40098 39528
rect 365438 39516 365444 39528
rect 365496 39516 365502 39568
rect 33134 39448 33140 39500
rect 33192 39488 33198 39500
rect 368106 39488 368112 39500
rect 33192 39460 368112 39488
rect 33192 39448 33198 39460
rect 368106 39448 368112 39460
rect 368164 39448 368170 39500
rect 26234 39380 26240 39432
rect 26292 39420 26298 39432
rect 368014 39420 368020 39432
rect 26292 39392 368020 39420
rect 26292 39380 26298 39392
rect 368014 39380 368020 39392
rect 368072 39380 368078 39432
rect 2774 39312 2780 39364
rect 2832 39352 2838 39364
rect 365346 39352 365352 39364
rect 2832 39324 365352 39352
rect 2832 39312 2838 39324
rect 365346 39312 365352 39324
rect 365404 39312 365410 39364
rect 80054 39244 80060 39296
rect 80112 39284 80118 39296
rect 363874 39284 363880 39296
rect 80112 39256 363880 39284
rect 80112 39244 80118 39256
rect 363874 39244 363880 39256
rect 363932 39244 363938 39296
rect 84194 39176 84200 39228
rect 84252 39216 84258 39228
rect 363966 39216 363972 39228
rect 84252 39188 363972 39216
rect 84252 39176 84258 39188
rect 363966 39176 363972 39188
rect 364024 39176 364030 39228
rect 115934 37204 115940 37256
rect 115992 37244 115998 37256
rect 372246 37244 372252 37256
rect 115992 37216 372252 37244
rect 115992 37204 115998 37216
rect 372246 37204 372252 37216
rect 372304 37204 372310 37256
rect 111794 37136 111800 37188
rect 111852 37176 111858 37188
rect 369302 37176 369308 37188
rect 111852 37148 369308 37176
rect 111852 37136 111858 37148
rect 369302 37136 369308 37148
rect 369360 37136 369366 37188
rect 109034 37068 109040 37120
rect 109092 37108 109098 37120
rect 369210 37108 369216 37120
rect 109092 37080 369216 37108
rect 109092 37068 109098 37080
rect 369210 37068 369216 37080
rect 369268 37068 369274 37120
rect 104894 37000 104900 37052
rect 104952 37040 104958 37052
rect 369118 37040 369124 37052
rect 104952 37012 369124 37040
rect 104952 37000 104958 37012
rect 369118 37000 369124 37012
rect 369176 37000 369182 37052
rect 102134 36932 102140 36984
rect 102192 36972 102198 36984
rect 366634 36972 366640 36984
rect 102192 36944 366640 36972
rect 102192 36932 102198 36944
rect 366634 36932 366640 36944
rect 366692 36932 366698 36984
rect 97994 36864 98000 36916
rect 98052 36904 98058 36916
rect 366726 36904 366732 36916
rect 98052 36876 366732 36904
rect 98052 36864 98058 36876
rect 366726 36864 366732 36876
rect 366784 36864 366790 36916
rect 93946 36796 93952 36848
rect 94004 36836 94010 36848
rect 366542 36836 366548 36848
rect 94004 36808 366548 36836
rect 94004 36796 94010 36808
rect 366542 36796 366548 36808
rect 366600 36796 366606 36848
rect 91094 36728 91100 36780
rect 91152 36768 91158 36780
rect 368198 36768 368204 36780
rect 91152 36740 368204 36768
rect 91152 36728 91158 36740
rect 368198 36728 368204 36740
rect 368256 36728 368262 36780
rect 86954 36660 86960 36712
rect 87012 36700 87018 36712
rect 366450 36700 366456 36712
rect 87012 36672 366456 36700
rect 87012 36660 87018 36672
rect 366450 36660 366456 36672
rect 366508 36660 366514 36712
rect 22094 36592 22100 36644
rect 22152 36632 22158 36644
rect 375098 36632 375104 36644
rect 22152 36604 375104 36632
rect 22152 36592 22158 36604
rect 375098 36592 375104 36604
rect 375156 36592 375162 36644
rect 17954 36524 17960 36576
rect 18012 36564 18018 36576
rect 372154 36564 372160 36576
rect 18012 36536 372160 36564
rect 18012 36524 18018 36536
rect 372154 36524 372160 36536
rect 372212 36524 372218 36576
rect 118786 36456 118792 36508
rect 118844 36496 118850 36508
rect 372338 36496 372344 36508
rect 118844 36468 372344 36496
rect 118844 36456 118850 36468
rect 372338 36456 372344 36468
rect 372396 36456 372402 36508
rect 122834 36388 122840 36440
rect 122892 36428 122898 36440
rect 371878 36428 371884 36440
rect 122892 36400 371884 36428
rect 122892 36388 122898 36400
rect 371878 36388 371884 36400
rect 371936 36388 371942 36440
rect 74534 34416 74540 34468
rect 74592 34456 74598 34468
rect 383102 34456 383108 34468
rect 74592 34428 383108 34456
rect 74592 34416 74598 34428
rect 383102 34416 383108 34428
rect 383160 34416 383166 34468
rect 462958 34416 462964 34468
rect 463016 34456 463022 34468
rect 536834 34456 536840 34468
rect 463016 34428 536840 34456
rect 463016 34416 463022 34428
rect 536834 34416 536840 34428
rect 536892 34416 536898 34468
rect 67634 34348 67640 34400
rect 67692 34388 67698 34400
rect 380434 34388 380440 34400
rect 67692 34360 380440 34388
rect 67692 34348 67698 34360
rect 380434 34348 380440 34360
rect 380492 34348 380498 34400
rect 70394 34280 70400 34332
rect 70452 34320 70458 34332
rect 383194 34320 383200 34332
rect 70452 34292 383200 34320
rect 70452 34280 70458 34292
rect 383194 34280 383200 34292
rect 383252 34280 383258 34332
rect 63494 34212 63500 34264
rect 63552 34252 63558 34264
rect 380342 34252 380348 34264
rect 63552 34224 380348 34252
rect 63552 34212 63558 34224
rect 380342 34212 380348 34224
rect 380400 34212 380406 34264
rect 60826 34144 60832 34196
rect 60884 34184 60890 34196
rect 381814 34184 381820 34196
rect 60884 34156 381820 34184
rect 60884 34144 60890 34156
rect 381814 34144 381820 34156
rect 381872 34144 381878 34196
rect 52454 34076 52460 34128
rect 52512 34116 52518 34128
rect 380158 34116 380164 34128
rect 52512 34088 380164 34116
rect 52512 34076 52518 34088
rect 380158 34076 380164 34088
rect 380216 34076 380222 34128
rect 49694 34008 49700 34060
rect 49752 34048 49758 34060
rect 380250 34048 380256 34060
rect 49752 34020 380256 34048
rect 49752 34008 49758 34020
rect 380250 34008 380256 34020
rect 380308 34008 380314 34060
rect 44266 33940 44272 33992
rect 44324 33980 44330 33992
rect 377582 33980 377588 33992
rect 44324 33952 377588 33980
rect 44324 33940 44330 33952
rect 377582 33940 377588 33952
rect 377640 33940 377646 33992
rect 34514 33872 34520 33924
rect 34572 33912 34578 33924
rect 374914 33912 374920 33924
rect 34572 33884 374920 33912
rect 34572 33872 34578 33884
rect 374914 33872 374920 33884
rect 374972 33872 374978 33924
rect 30374 33804 30380 33856
rect 30432 33844 30438 33856
rect 375006 33844 375012 33856
rect 30432 33816 375012 33844
rect 30432 33804 30438 33816
rect 375006 33804 375012 33816
rect 375064 33804 375070 33856
rect 9674 33736 9680 33788
rect 9732 33776 9738 33788
rect 377674 33776 377680 33788
rect 9732 33748 377680 33776
rect 9732 33736 9738 33748
rect 377674 33736 377680 33748
rect 377732 33736 377738 33788
rect 77386 33668 77392 33720
rect 77444 33708 77450 33720
rect 383286 33708 383292 33720
rect 77444 33680 383292 33708
rect 77444 33668 77450 33680
rect 383286 33668 383292 33680
rect 383344 33668 383350 33720
rect 85666 33600 85672 33652
rect 85724 33640 85730 33652
rect 386230 33640 386236 33652
rect 85724 33612 386236 33640
rect 85724 33600 85730 33612
rect 386230 33600 386236 33612
rect 386288 33600 386294 33652
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 378778 33096 378784 33108
rect 3568 33068 378784 33096
rect 3568 33056 3574 33068
rect 378778 33056 378784 33068
rect 378836 33056 378842 33108
rect 563698 33056 563704 33108
rect 563756 33096 563762 33108
rect 580166 33096 580172 33108
rect 563756 33068 580172 33096
rect 563756 33056 563762 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 3418 31696 3424 31748
rect 3476 31736 3482 31748
rect 460198 31736 460204 31748
rect 3476 31708 460204 31736
rect 3476 31696 3482 31708
rect 460198 31696 460204 31708
rect 460256 31696 460262 31748
rect 120074 31628 120080 31680
rect 120132 31668 120138 31680
rect 364978 31668 364984 31680
rect 120132 31640 364984 31668
rect 120132 31628 120138 31640
rect 364978 31628 364984 31640
rect 365036 31628 365042 31680
rect 384206 31628 384212 31680
rect 384264 31668 384270 31680
rect 462314 31668 462320 31680
rect 384264 31640 462320 31668
rect 384264 31628 384270 31640
rect 462314 31628 462320 31640
rect 462372 31628 462378 31680
rect 113174 31560 113180 31612
rect 113232 31600 113238 31612
rect 370590 31600 370596 31612
rect 113232 31572 370596 31600
rect 113232 31560 113238 31572
rect 370590 31560 370596 31572
rect 370648 31560 370654 31612
rect 102226 31492 102232 31544
rect 102284 31532 102290 31544
rect 373350 31532 373356 31544
rect 102284 31504 373356 31532
rect 102284 31492 102290 31504
rect 373350 31492 373356 31504
rect 373408 31492 373414 31544
rect 111058 31424 111064 31476
rect 111116 31464 111122 31476
rect 386046 31464 386052 31476
rect 111116 31436 386052 31464
rect 111116 31424 111122 31436
rect 386046 31424 386052 31436
rect 386104 31424 386110 31476
rect 99374 31356 99380 31408
rect 99432 31396 99438 31408
rect 376018 31396 376024 31408
rect 99432 31368 376024 31396
rect 99432 31356 99438 31368
rect 376018 31356 376024 31368
rect 376076 31356 376082 31408
rect 92474 31288 92480 31340
rect 92532 31328 92538 31340
rect 378870 31328 378876 31340
rect 92532 31300 378876 31328
rect 92532 31288 92538 31300
rect 378870 31288 378876 31300
rect 378928 31288 378934 31340
rect 35894 31220 35900 31272
rect 35952 31260 35958 31272
rect 369394 31260 369400 31272
rect 35952 31232 369400 31260
rect 35952 31220 35958 31232
rect 369394 31220 369400 31232
rect 369452 31220 369458 31272
rect 19334 31152 19340 31204
rect 19392 31192 19398 31204
rect 363782 31192 363788 31204
rect 19392 31164 363788 31192
rect 19392 31152 19398 31164
rect 363782 31152 363788 31164
rect 363840 31152 363846 31204
rect 31754 31084 31760 31136
rect 31812 31124 31818 31136
rect 384942 31124 384948 31136
rect 31812 31096 384948 31124
rect 31812 31084 31818 31096
rect 384942 31084 384948 31096
rect 385000 31084 385006 31136
rect 13814 31016 13820 31068
rect 13872 31056 13878 31068
rect 385954 31056 385960 31068
rect 13872 31028 385960 31056
rect 13872 31016 13878 31028
rect 385954 31016 385960 31028
rect 386012 31016 386018 31068
rect 117314 30948 117320 31000
rect 117372 30988 117378 31000
rect 360838 30988 360844 31000
rect 117372 30960 360844 30988
rect 117372 30948 117378 30960
rect 360838 30948 360844 30960
rect 360896 30948 360902 31000
rect 124214 30880 124220 30932
rect 124272 30920 124278 30932
rect 366358 30920 366364 30932
rect 124272 30892 366364 30920
rect 124272 30880 124278 30892
rect 366358 30880 366364 30892
rect 366416 30880 366422 30932
rect 106918 28364 106924 28416
rect 106976 28404 106982 28416
rect 377490 28404 377496 28416
rect 106976 28376 377496 28404
rect 106976 28364 106982 28376
rect 377490 28364 377496 28376
rect 377548 28364 377554 28416
rect 45554 28296 45560 28348
rect 45612 28336 45618 28348
rect 374822 28336 374828 28348
rect 45612 28308 374828 28336
rect 45612 28296 45618 28308
rect 374822 28296 374828 28308
rect 374880 28296 374886 28348
rect 38654 28228 38660 28280
rect 38712 28268 38718 28280
rect 372062 28268 372068 28280
rect 38712 28240 372068 28268
rect 38712 28228 38718 28240
rect 372062 28228 372068 28240
rect 372120 28228 372126 28280
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 363690 20652 363696 20664
rect 3476 20624 363696 20652
rect 3476 20612 3482 20624
rect 363690 20612 363696 20624
rect 363748 20612 363754 20664
rect 562318 20612 562324 20664
rect 562376 20652 562382 20664
rect 579982 20652 579988 20664
rect 562376 20624 579988 20652
rect 562376 20612 562382 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 566 7556 572 7608
rect 624 7596 630 7608
rect 367738 7596 367744 7608
rect 624 7568 367744 7596
rect 624 7556 630 7568
rect 367738 7556 367744 7568
rect 367796 7556 367802 7608
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 374638 6848 374644 6860
rect 3476 6820 374644 6848
rect 3476 6808 3482 6820
rect 374638 6808 374644 6820
rect 374696 6808 374702 6860
rect 565078 6808 565084 6860
rect 565136 6848 565142 6860
rect 580166 6848 580172 6860
rect 565136 6820 580172 6848
rect 565136 6808 565142 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 89162 4088 89168 4140
rect 89220 4128 89226 4140
rect 363598 4128 363604 4140
rect 89220 4100 363604 4128
rect 89220 4088 89226 4100
rect 363598 4088 363604 4100
rect 363656 4088 363662 4140
rect 82078 4020 82084 4072
rect 82136 4060 82142 4072
rect 359642 4060 359648 4072
rect 82136 4032 359648 4060
rect 82136 4020 82142 4032
rect 359642 4020 359648 4032
rect 359700 4020 359706 4072
rect 56042 3952 56048 4004
rect 56100 3992 56106 4004
rect 359458 3992 359464 4004
rect 56100 3964 359464 3992
rect 56100 3952 56106 3964
rect 359458 3952 359464 3964
rect 359516 3952 359522 4004
rect 57238 3884 57244 3936
rect 57296 3924 57302 3936
rect 371970 3924 371976 3936
rect 57296 3896 371976 3924
rect 57296 3884 57302 3896
rect 371970 3884 371976 3896
rect 372028 3884 372034 3936
rect 48958 3816 48964 3868
rect 49016 3856 49022 3868
rect 365070 3856 365076 3868
rect 49016 3828 365076 3856
rect 49016 3816 49022 3828
rect 365070 3816 365076 3828
rect 365128 3816 365134 3868
rect 43070 3748 43076 3800
rect 43128 3788 43134 3800
rect 361114 3788 361120 3800
rect 43128 3760 361120 3788
rect 43128 3748 43134 3760
rect 361114 3748 361120 3760
rect 361172 3748 361178 3800
rect 52546 3680 52552 3732
rect 52604 3720 52610 3732
rect 382918 3720 382924 3732
rect 52604 3692 382924 3720
rect 52604 3680 52610 3692
rect 382918 3680 382924 3692
rect 382976 3680 382982 3732
rect 37182 3612 37188 3664
rect 37240 3652 37246 3664
rect 367922 3652 367928 3664
rect 37240 3624 367928 3652
rect 37240 3612 37246 3624
rect 367922 3612 367928 3624
rect 367980 3612 367986 3664
rect 41874 3544 41880 3596
rect 41932 3584 41938 3596
rect 377398 3584 377404 3596
rect 41932 3556 377404 3584
rect 41932 3544 41938 3556
rect 377398 3544 377404 3556
rect 377456 3544 377462 3596
rect 27706 3476 27712 3528
rect 27764 3516 27770 3528
rect 374730 3516 374736 3528
rect 27764 3488 374736 3516
rect 27764 3476 27770 3488
rect 374730 3476 374736 3488
rect 374788 3476 374794 3528
rect 38378 3408 38384 3460
rect 38436 3448 38442 3460
rect 385678 3448 385684 3460
rect 38436 3420 385684 3448
rect 38436 3408 38442 3420
rect 385678 3408 385684 3420
rect 385736 3408 385742 3460
rect 60734 3340 60740 3392
rect 60792 3380 60798 3392
rect 61654 3380 61660 3392
rect 60792 3352 61660 3380
rect 60792 3340 60798 3352
rect 61654 3340 61660 3352
rect 61712 3340 61718 3392
rect 85574 3340 85580 3392
rect 85632 3380 85638 3392
rect 86494 3380 86500 3392
rect 85632 3352 86500 3380
rect 85632 3340 85638 3352
rect 86494 3340 86500 3352
rect 86552 3340 86558 3392
rect 96246 3340 96252 3392
rect 96304 3380 96310 3392
rect 359550 3380 359556 3392
rect 96304 3352 359556 3380
rect 96304 3340 96310 3352
rect 359550 3340 359556 3352
rect 359608 3340 359614 3392
rect 110414 3272 110420 3324
rect 110472 3312 110478 3324
rect 111610 3312 111616 3324
rect 110472 3284 111616 3312
rect 110472 3272 110478 3284
rect 111610 3272 111616 3284
rect 111668 3272 111674 3324
rect 361206 3312 361212 3324
rect 111812 3284 361212 3312
rect 6454 3204 6460 3256
rect 6512 3244 6518 3256
rect 106826 3244 106832 3256
rect 6512 3216 106832 3244
rect 6512 3204 6518 3216
rect 106826 3204 106832 3216
rect 106884 3204 106890 3256
rect 28902 3136 28908 3188
rect 28960 3176 28966 3188
rect 28960 3148 103514 3176
rect 28960 3136 28966 3148
rect 103486 3108 103514 3148
rect 106918 3136 106924 3188
rect 106976 3176 106982 3188
rect 111812 3176 111840 3284
rect 361206 3272 361212 3284
rect 361264 3272 361270 3324
rect 360930 3244 360936 3256
rect 106976 3148 111840 3176
rect 113146 3216 360936 3244
rect 106976 3136 106982 3148
rect 111058 3108 111064 3120
rect 103486 3080 111064 3108
rect 111058 3068 111064 3080
rect 111116 3068 111122 3120
rect 110506 3000 110512 3052
rect 110564 3040 110570 3052
rect 113146 3040 113174 3216
rect 360930 3204 360936 3216
rect 360988 3204 360994 3256
rect 110564 3012 113174 3040
rect 110564 3000 110570 3012
rect 30098 2116 30104 2168
rect 30156 2156 30162 2168
rect 367830 2156 367836 2168
rect 30156 2128 367836 2156
rect 30156 2116 30162 2128
rect 367830 2116 367836 2128
rect 367888 2116 367894 2168
rect 2866 2048 2872 2100
rect 2924 2088 2930 2100
rect 384298 2088 384304 2100
rect 2924 2060 384304 2088
rect 2924 2048 2930 2060
rect 384298 2048 384304 2060
rect 384356 2048 384362 2100
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 429844 700748 429896 700800
rect 445116 700748 445168 700800
rect 364984 700680 365036 700732
rect 445024 700680 445076 700732
rect 332508 700612 332560 700664
rect 446496 700612 446548 700664
rect 300124 700544 300176 700596
rect 449164 700544 449216 700596
rect 283840 700476 283892 700528
rect 446404 700476 446456 700528
rect 154120 700408 154172 700460
rect 416044 700408 416096 700460
rect 444288 700408 444340 700460
rect 494796 700408 494848 700460
rect 105452 700340 105504 700392
rect 445208 700340 445260 700392
rect 445668 700340 445720 700392
rect 478512 700340 478564 700392
rect 40500 700272 40552 700324
rect 449256 700272 449308 700324
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 347780 685312 347832 685364
rect 446680 685312 446732 685364
rect 218060 685244 218112 685296
rect 446588 685244 446640 685296
rect 88340 685176 88392 685228
rect 416228 685176 416280 685228
rect 71780 685108 71832 685160
rect 419356 685108 419408 685160
rect 19984 684768 20036 684820
rect 419448 684768 419500 684820
rect 3976 684700 4028 684752
rect 418804 684700 418856 684752
rect 3608 684632 3660 684684
rect 418988 684632 419040 684684
rect 3424 684564 3476 684616
rect 419080 684564 419132 684616
rect 3332 684496 3384 684548
rect 418896 684496 418948 684548
rect 266360 683748 266412 683800
rect 446864 683748 446916 683800
rect 20812 683544 20864 683596
rect 359464 683544 359516 683596
rect 21364 683476 21416 683528
rect 416136 683476 416188 683528
rect 3884 683408 3936 683460
rect 419172 683408 419224 683460
rect 3516 683340 3568 683392
rect 419264 683340 419316 683392
rect 4068 683272 4120 683324
rect 420184 683272 420236 683324
rect 3792 683204 3844 683256
rect 445392 683204 445444 683256
rect 3240 683136 3292 683188
rect 445484 683136 445536 683188
rect 3148 682660 3200 682712
rect 420552 682660 420604 682712
rect 20076 681708 20128 681760
rect 20812 681708 20864 681760
rect 3516 679192 3568 679244
rect 3516 678988 3568 679040
rect 361764 678988 361816 679040
rect 365076 678988 365128 679040
rect 3700 678512 3752 678564
rect 3884 678172 3936 678224
rect 17684 670692 17736 670744
rect 20076 670692 20128 670744
rect 450636 669944 450688 669996
rect 462320 669944 462372 669996
rect 361764 667904 361816 667956
rect 381544 667904 381596 667956
rect 13820 667360 13872 667412
rect 17684 667360 17736 667412
rect 11796 665116 11848 665168
rect 13820 665184 13872 665236
rect 7564 659608 7616 659660
rect 11796 659676 11848 659728
rect 3148 658180 3200 658232
rect 19984 658180 20036 658232
rect 361764 656888 361816 656940
rect 406384 656888 406436 656940
rect 6184 655528 6236 655580
rect 7564 655528 7616 655580
rect 4804 652740 4856 652792
rect 6184 652740 6236 652792
rect 361764 645872 361816 645924
rect 378784 645872 378836 645924
rect 569224 643084 569276 643136
rect 579620 643084 579672 643136
rect 361580 634788 361632 634840
rect 407764 634788 407816 634840
rect 3700 631320 3752 631372
rect 20904 631320 20956 631372
rect 567844 630640 567896 630692
rect 580172 630640 580224 630692
rect 361580 623772 361632 623824
rect 376024 623772 376076 623824
rect 571984 616836 572036 616888
rect 580172 616836 580224 616888
rect 359464 616768 359516 616820
rect 360936 616768 360988 616820
rect 361580 612756 361632 612808
rect 410524 612756 410576 612808
rect 360936 611192 360988 611244
rect 362224 611192 362276 611244
rect 458732 603712 458784 603764
rect 459008 603712 459060 603764
rect 361764 601672 361816 601724
rect 374644 601672 374696 601724
rect 362224 600244 362276 600296
rect 362960 600244 363012 600296
rect 457628 600244 457680 600296
rect 461584 600244 461636 600296
rect 459008 599836 459060 599888
rect 463700 599836 463752 599888
rect 458824 599700 458876 599752
rect 465080 599700 465132 599752
rect 457536 599632 457588 599684
rect 469864 599632 469916 599684
rect 457444 599564 457496 599616
rect 469956 599564 470008 599616
rect 459928 598408 459980 598460
rect 463792 598408 463844 598460
rect 458640 598340 458692 598392
rect 465172 598340 465224 598392
rect 488632 598340 488684 598392
rect 494244 598340 494296 598392
rect 449900 598272 449952 598324
rect 526720 598272 526772 598324
rect 457904 598204 457956 598256
rect 468484 598204 468536 598256
rect 482284 598204 482336 598256
rect 494060 598204 494112 598256
rect 493324 598136 493376 598188
rect 494980 598136 495032 598188
rect 519544 598136 519596 598188
rect 520372 598136 520424 598188
rect 473268 598068 473320 598120
rect 475936 598068 475988 598120
rect 457352 596844 457404 596896
rect 465724 596844 465776 596896
rect 362960 596776 363012 596828
rect 368388 596776 368440 596828
rect 449808 596776 449860 596828
rect 469588 596776 469640 596828
rect 361764 590656 361816 590708
rect 371976 590656 372028 590708
rect 567936 590656 567988 590708
rect 580172 590656 580224 590708
rect 368480 589296 368532 589348
rect 372804 589228 372856 589280
rect 372804 584400 372856 584452
rect 379520 584400 379572 584452
rect 379520 582632 379572 582684
rect 381636 582632 381688 582684
rect 361764 579640 361816 579692
rect 370504 579640 370556 579692
rect 361764 568556 361816 568608
rect 367744 568556 367796 568608
rect 459652 564340 459704 564392
rect 462320 564340 462372 564392
rect 577504 563048 577556 563100
rect 579620 563048 579672 563100
rect 381636 559308 381688 559360
rect 383752 559308 383804 559360
rect 361580 557744 361632 557796
rect 363604 557744 363656 557796
rect 383752 554140 383804 554192
rect 385684 554140 385736 554192
rect 385684 550536 385736 550588
rect 387432 550536 387484 550588
rect 361580 546592 361632 546644
rect 363696 546592 363748 546644
rect 387432 546456 387484 546508
rect 388444 546456 388496 546508
rect 457720 543056 457772 543108
rect 464344 543056 464396 543108
rect 459836 542988 459888 543040
rect 466460 542988 466512 543040
rect 361580 535712 361632 535764
rect 363788 535712 363840 535764
rect 388444 535440 388496 535492
rect 389824 535440 389876 535492
rect 448336 526396 448388 526448
rect 500960 526396 501012 526448
rect 389824 524492 389876 524544
rect 391204 524492 391256 524544
rect 361764 524424 361816 524476
rect 411904 524424 411956 524476
rect 515404 524424 515456 524476
rect 580172 524424 580224 524476
rect 448244 522248 448296 522300
rect 493324 522248 493376 522300
rect 448428 520888 448480 520940
rect 506480 520888 506532 520940
rect 462964 520412 463016 520464
rect 488632 520412 488684 520464
rect 472900 520344 472952 520396
rect 473268 520344 473320 520396
rect 494244 520344 494296 520396
rect 458088 520004 458140 520056
rect 463056 520004 463108 520056
rect 457260 519596 457312 519648
rect 467932 519596 467984 519648
rect 448060 519528 448112 519580
rect 472900 519528 472952 519580
rect 459744 518712 459796 518764
rect 462504 518712 462556 518764
rect 457812 518372 457864 518424
rect 466552 518372 466604 518424
rect 459560 518304 459612 518356
rect 470692 518304 470744 518356
rect 459100 518236 459152 518288
rect 470876 518236 470928 518288
rect 447968 518168 448020 518220
rect 462412 518168 462464 518220
rect 457996 517964 458048 518016
rect 461676 517964 461728 518016
rect 391204 517488 391256 517540
rect 480168 517488 480220 517540
rect 482652 517488 482704 517540
rect 394608 517420 394660 517472
rect 448428 516128 448480 516180
rect 491852 516128 491904 516180
rect 494060 515380 494112 515432
rect 538220 515380 538272 515432
rect 3976 514768 4028 514820
rect 4804 514768 4856 514820
rect 361764 513340 361816 513392
rect 414664 513340 414716 513392
rect 494060 511980 494112 512032
rect 535460 511980 535512 512032
rect 394700 510620 394752 510672
rect 402244 510552 402296 510604
rect 494244 508512 494296 508564
rect 532700 508512 532752 508564
rect 494980 505112 495032 505164
rect 529940 505112 529992 505164
rect 361764 502324 361816 502376
rect 416320 502324 416372 502376
rect 448520 500216 448572 500268
rect 545120 500216 545172 500268
rect 450084 499808 450136 499860
rect 450728 499808 450780 499860
rect 447324 499536 447376 499588
rect 449716 499536 449768 499588
rect 447876 499468 447928 499520
rect 494060 499468 494112 499520
rect 447968 499400 448020 499452
rect 494152 499400 494204 499452
rect 448244 498856 448296 498908
rect 542452 498856 542504 498908
rect 449716 498788 449768 498840
rect 547880 498788 547932 498840
rect 452016 497564 452068 497616
rect 481640 497564 481692 497616
rect 449808 497496 449860 497548
rect 486240 497496 486292 497548
rect 451924 497428 451976 497480
rect 488632 497428 488684 497480
rect 454040 497088 454092 497140
rect 459560 497088 459612 497140
rect 454132 497020 454184 497072
rect 458088 497020 458140 497072
rect 455420 496952 455472 497004
rect 461032 496952 461084 497004
rect 452844 496884 452896 496936
rect 455144 496884 455196 496936
rect 451372 496816 451424 496868
rect 453672 496816 453724 496868
rect 454684 496816 454736 496868
rect 456616 496816 456668 496868
rect 569316 484372 569368 484424
rect 580172 484372 580224 484424
rect 361764 480224 361816 480276
rect 418712 480224 418764 480276
rect 511264 470568 511316 470620
rect 579988 470568 580040 470620
rect 402244 469276 402296 469328
rect 405004 469276 405056 469328
rect 361764 469208 361816 469260
rect 417424 469208 417476 469260
rect 494704 462476 494756 462528
rect 527640 462476 527692 462528
rect 436100 462408 436152 462460
rect 554136 462408 554188 462460
rect 433248 462340 433300 462392
rect 551192 462340 551244 462392
rect 515496 461660 515548 461712
rect 542360 461660 542412 461712
rect 480168 461592 480220 461644
rect 521752 461592 521804 461644
rect 449992 460912 450044 460964
rect 524420 460912 524472 460964
rect 361764 458192 361816 458244
rect 382924 458192 382976 458244
rect 449440 457444 449492 457496
rect 487160 457444 487212 457496
rect 473728 456764 473780 456816
rect 480168 456764 480220 456816
rect 449532 456016 449584 456068
rect 484400 456016 484452 456068
rect 488264 456016 488316 456068
rect 494704 456016 494756 456068
rect 450176 455472 450228 455524
rect 480996 455472 481048 455524
rect 422300 455404 422352 455456
rect 473728 455404 473780 455456
rect 405004 455336 405056 455388
rect 406476 455336 406528 455388
rect 450268 454792 450320 454844
rect 480260 454792 480312 454844
rect 449716 454724 449768 454776
rect 481916 454724 481968 454776
rect 449624 454656 449676 454708
rect 483112 454656 483164 454708
rect 406476 450916 406528 450968
rect 408500 450916 408552 450968
rect 427452 447108 427504 447160
rect 446956 447108 447008 447160
rect 432420 445748 432472 445800
rect 433248 445748 433300 445800
rect 444104 445748 444156 445800
rect 436100 445680 436152 445732
rect 437388 445680 437440 445732
rect 437296 444524 437348 444576
rect 445852 444524 445904 444576
rect 442632 444456 442684 444508
rect 445760 444456 445812 444508
rect 422760 444388 422812 444440
rect 445576 444388 445628 444440
rect 408500 441600 408552 441652
rect 413744 441532 413796 441584
rect 413744 437520 413796 437572
rect 414756 437520 414808 437572
rect 361764 436092 361816 436144
rect 418620 436092 418672 436144
rect 414756 431332 414808 431384
rect 416688 431332 416740 431384
rect 569408 430584 569460 430636
rect 580172 430584 580224 430636
rect 456892 429836 456944 429888
rect 474280 429836 474332 429888
rect 478144 429156 478196 429208
rect 479616 429156 479668 429208
rect 482284 429156 482336 429208
rect 484952 429156 485004 429208
rect 486424 429156 486476 429208
rect 487620 429156 487672 429208
rect 416688 429020 416740 429072
rect 420368 429020 420420 429072
rect 457444 428408 457496 428460
rect 471612 428408 471664 428460
rect 529204 423580 529256 423632
rect 530216 423580 530268 423632
rect 530584 423580 530636 423632
rect 532792 423580 532844 423632
rect 502984 423512 503036 423564
rect 523776 423512 523828 423564
rect 522304 423444 522356 423496
rect 549536 423444 549588 423496
rect 483020 423376 483072 423428
rect 522488 423376 522540 423428
rect 523684 423376 523736 423428
rect 552112 423376 552164 423428
rect 485780 423308 485832 423360
rect 526352 423308 526404 423360
rect 526444 423308 526496 423360
rect 554688 423308 554740 423360
rect 487160 423240 487212 423292
rect 528928 423240 528980 423292
rect 488540 423172 488592 423224
rect 531504 423172 531556 423224
rect 496820 423104 496872 423156
rect 545672 423104 545724 423156
rect 498200 423036 498252 423088
rect 548248 423036 548300 423088
rect 499580 422968 499632 423020
rect 550824 422968 550876 423020
rect 501052 422900 501104 422952
rect 553400 422900 553452 422952
rect 483112 421540 483164 421592
rect 521200 421540 521252 421592
rect 494060 420180 494112 420232
rect 541808 420180 541860 420232
rect 362408 418752 362460 418804
rect 440884 418752 440936 418804
rect 420368 418140 420420 418192
rect 426440 418072 426492 418124
rect 425980 417732 426032 417784
rect 507860 417732 507912 417784
rect 421472 417664 421524 417716
rect 503720 417664 503772 417716
rect 424692 417596 424744 417648
rect 506480 417596 506532 417648
rect 424048 417528 424100 417580
rect 506572 417528 506624 417580
rect 425336 417460 425388 417512
rect 507952 417460 508004 417512
rect 422116 417392 422168 417444
rect 503996 417392 504048 417444
rect 362316 416032 362368 416084
rect 436744 416032 436796 416084
rect 426440 415624 426492 415676
rect 429844 415624 429896 415676
rect 361580 413992 361632 414044
rect 439504 413992 439556 414044
rect 429844 410184 429896 410236
rect 431224 410184 431276 410236
rect 361580 402976 361632 403028
rect 442264 402976 442316 403028
rect 502616 402228 502668 402280
rect 557540 402228 557592 402280
rect 497464 400868 497516 400920
rect 546500 400868 546552 400920
rect 494152 399440 494204 399492
rect 539600 399440 539652 399492
rect 431224 398760 431276 398812
rect 432604 398760 432656 398812
rect 492680 398080 492732 398132
rect 538220 398080 538272 398132
rect 492772 396720 492824 396772
rect 536840 396720 536892 396772
rect 461400 395292 461452 395344
rect 490012 395292 490064 395344
rect 491576 395292 491628 395344
rect 535460 395292 535512 395344
rect 458456 393932 458508 393984
rect 478144 393932 478196 393984
rect 491392 393932 491444 393984
rect 534172 393932 534224 393984
rect 458180 392640 458232 392692
rect 476120 392640 476172 392692
rect 461124 392572 461176 392624
rect 486424 392572 486476 392624
rect 490564 392572 490616 392624
rect 534080 392572 534132 392624
rect 361580 391960 361632 392012
rect 440976 392028 441028 392080
rect 432604 391960 432656 392012
rect 433984 391960 434036 392012
rect 460388 391348 460440 391400
rect 482284 391348 482336 391400
rect 450452 391280 450504 391332
rect 491300 391280 491352 391332
rect 496452 391280 496504 391332
rect 543740 391280 543792 391332
rect 422392 391212 422444 391264
rect 506020 391212 506072 391264
rect 461676 389852 461728 389904
rect 481640 389852 481692 389904
rect 495716 389852 495768 389904
rect 542360 389852 542412 389904
rect 422300 389784 422352 389836
rect 505284 389784 505336 389836
rect 450084 389240 450136 389292
rect 450728 389240 450780 389292
rect 454040 389240 454092 389292
rect 454868 389240 454920 389292
rect 465080 389240 465132 389292
rect 465908 389240 465960 389292
rect 483020 389240 483072 389292
rect 483572 389240 483624 389292
rect 492680 389240 492732 389292
rect 493140 389240 493192 389292
rect 494060 389240 494112 389292
rect 494612 389240 494664 389292
rect 506480 389240 506532 389292
rect 507124 389240 507176 389292
rect 507860 389240 507912 389292
rect 508596 389240 508648 389292
rect 453764 389104 453816 389156
rect 454684 389104 454736 389156
rect 469956 388900 470008 388952
rect 477316 388900 477368 388952
rect 484676 388900 484728 388952
rect 502984 388900 503036 388952
rect 468484 388832 468536 388884
rect 475844 388832 475896 388884
rect 500868 388832 500920 388884
rect 523684 388832 523736 388884
rect 468576 388764 468628 388816
rect 481732 388764 481784 388816
rect 499396 388764 499448 388816
rect 522304 388764 522356 388816
rect 469864 388696 469916 388748
rect 478052 388696 478104 388748
rect 502340 388696 502392 388748
rect 526444 388696 526496 388748
rect 467104 388628 467156 388680
rect 482468 388628 482520 388680
rect 485412 388628 485464 388680
rect 524420 388628 524472 388680
rect 463056 388560 463108 388612
rect 480996 388560 481048 388612
rect 486884 388560 486936 388612
rect 527180 388560 527232 388612
rect 461584 388492 461636 388544
rect 478788 388492 478840 388544
rect 489828 388492 489880 388544
rect 530584 388492 530636 388544
rect 456708 388424 456760 388476
rect 457444 388424 457496 388476
rect 461768 388424 461820 388476
rect 480260 388424 480312 388476
rect 488356 388424 488408 388476
rect 529204 388424 529256 388476
rect 464344 388016 464396 388068
rect 469220 388016 469272 388068
rect 465724 387948 465776 388000
rect 469956 387948 470008 388000
rect 459652 387812 459704 387864
rect 461676 387812 461728 387864
rect 447692 387404 447744 387456
rect 452016 387404 452068 387456
rect 447784 387200 447836 387252
rect 462964 387200 463016 387252
rect 448980 387132 449032 387184
rect 491116 387132 491168 387184
rect 449072 387064 449124 387116
rect 513380 387064 513432 387116
rect 445576 386588 445628 386640
rect 553952 386588 554004 386640
rect 371884 386520 371936 386572
rect 512276 386520 512328 386572
rect 364984 386452 365036 386504
rect 512184 386452 512236 386504
rect 360844 386384 360896 386436
rect 512092 386384 512144 386436
rect 448428 385976 448480 386028
rect 451924 385976 451976 386028
rect 450360 385092 450412 385144
rect 563428 385092 563480 385144
rect 366364 385024 366416 385076
rect 512000 385024 512052 385076
rect 365076 384956 365128 385008
rect 447140 384956 447192 385008
rect 512736 383732 512788 383784
rect 530584 383732 530636 383784
rect 513288 383664 513340 383716
rect 547144 383664 547196 383716
rect 381544 383596 381596 383648
rect 447140 383596 447192 383648
rect 406384 383528 406436 383580
rect 447232 383528 447284 383580
rect 512000 383528 512052 383580
rect 512552 383528 512604 383580
rect 512828 382984 512880 383036
rect 518164 382984 518216 383036
rect 512460 382440 512512 382492
rect 515588 382440 515640 382492
rect 513012 382372 513064 382424
rect 519636 382372 519688 382424
rect 378784 382168 378836 382220
rect 447140 382168 447192 382220
rect 407764 382100 407816 382152
rect 447232 382100 447284 382152
rect 361580 380876 361632 380928
rect 442356 380876 442408 380928
rect 513288 380876 513340 380928
rect 549904 380876 549956 380928
rect 376024 380808 376076 380860
rect 447140 380808 447192 380860
rect 410524 380740 410576 380792
rect 447232 380740 447284 380792
rect 512092 379856 512144 379908
rect 514116 379856 514168 379908
rect 513288 379516 513340 379568
rect 544384 379516 544436 379568
rect 371976 379448 372028 379500
rect 447232 379448 447284 379500
rect 374644 379380 374696 379432
rect 447140 379380 447192 379432
rect 512184 378292 512236 378344
rect 522304 378292 522356 378344
rect 513288 378224 513340 378276
rect 548524 378224 548576 378276
rect 514024 378156 514076 378208
rect 579804 378156 579856 378208
rect 367744 378088 367796 378140
rect 447232 378088 447284 378140
rect 370504 378020 370556 378072
rect 447140 378020 447192 378072
rect 512828 377408 512880 377460
rect 549996 377408 550048 377460
rect 513288 376796 513340 376848
rect 517520 376796 517572 376848
rect 363696 376660 363748 376712
rect 447232 376660 447284 376712
rect 363604 376592 363656 376644
rect 447140 376592 447192 376644
rect 512368 375980 512420 376032
rect 547236 375980 547288 376032
rect 512460 375504 512512 375556
rect 520280 375504 520332 375556
rect 512736 375368 512788 375420
rect 516140 375368 516192 375420
rect 363788 375300 363840 375352
rect 447140 375300 447192 375352
rect 411904 375232 411956 375284
rect 447232 375232 447284 375284
rect 513288 374008 513340 374060
rect 518900 374008 518952 374060
rect 414664 373940 414716 373992
rect 447140 373940 447192 373992
rect 416320 373872 416372 373924
rect 447232 373872 447284 373924
rect 512644 373328 512696 373380
rect 517704 373328 517756 373380
rect 513288 372648 513340 372700
rect 518992 372648 519044 372700
rect 512644 372580 512696 372632
rect 523040 372580 523092 372632
rect 362224 372512 362276 372564
rect 447140 372512 447192 372564
rect 418712 372444 418764 372496
rect 447232 372444 447284 372496
rect 433984 371492 434036 371544
rect 435364 371492 435416 371544
rect 512092 371356 512144 371408
rect 514852 371356 514904 371408
rect 382924 371152 382976 371204
rect 447232 371152 447284 371204
rect 417424 371084 417476 371136
rect 447140 371084 447192 371136
rect 512092 370948 512144 371000
rect 514760 370948 514812 371000
rect 361580 369860 361632 369912
rect 429200 369860 429252 369912
rect 418620 369792 418672 369844
rect 447232 369792 447284 369844
rect 436744 369724 436796 369776
rect 447140 369724 447192 369776
rect 512276 368840 512328 368892
rect 514944 368840 514996 368892
rect 512736 368500 512788 368552
rect 516232 368500 516284 368552
rect 439504 368432 439556 368484
rect 447232 368432 447284 368484
rect 440884 368364 440936 368416
rect 447140 368364 447192 368416
rect 513288 367344 513340 367396
rect 520372 367344 520424 367396
rect 512000 367140 512052 367192
rect 514208 367140 514260 367192
rect 440976 367004 441028 367056
rect 447140 367004 447192 367056
rect 442264 366936 442316 366988
rect 447232 366936 447284 366988
rect 513288 365848 513340 365900
rect 517796 365848 517848 365900
rect 513012 365712 513064 365764
rect 516784 365712 516836 365764
rect 429200 365644 429252 365696
rect 447140 365644 447192 365696
rect 442356 365576 442408 365628
rect 447232 365576 447284 365628
rect 569500 364352 569552 364404
rect 580172 364352 580224 364404
rect 512000 363332 512052 363384
rect 513748 363332 513800 363384
rect 513288 363264 513340 363316
rect 517612 363264 517664 363316
rect 436928 362992 436980 363044
rect 447140 362992 447192 363044
rect 432604 362924 432656 362976
rect 447232 362924 447284 362976
rect 442264 361632 442316 361684
rect 447232 361632 447284 361684
rect 439688 361564 439740 361616
rect 447140 361564 447192 361616
rect 512000 361224 512052 361276
rect 513656 361224 513708 361276
rect 435548 360272 435600 360324
rect 435364 360204 435416 360256
rect 438124 360204 438176 360256
rect 441068 360272 441120 360324
rect 447140 360272 447192 360324
rect 447232 360204 447284 360256
rect 513288 360204 513340 360256
rect 520464 360204 520516 360256
rect 548524 360136 548576 360188
rect 552020 360136 552072 360188
rect 549904 359116 549956 359168
rect 558184 359116 558236 359168
rect 544384 359048 544436 359100
rect 553768 359048 553820 359100
rect 547144 358980 547196 359032
rect 565544 358980 565596 359032
rect 522304 358912 522356 358964
rect 550824 358912 550876 358964
rect 442356 358844 442408 358896
rect 447232 358844 447284 358896
rect 512644 358844 512696 358896
rect 516416 358844 516468 358896
rect 530584 358844 530636 358896
rect 567016 358844 567068 358896
rect 436836 358776 436888 358828
rect 447140 358776 447192 358828
rect 514116 358776 514168 358828
rect 555240 358776 555292 358828
rect 549996 358708 550048 358760
rect 556712 358708 556764 358760
rect 518164 358640 518216 358692
rect 562600 358640 562652 358692
rect 519636 358572 519688 358624
rect 564072 358572 564124 358624
rect 547236 358504 547288 358556
rect 559656 358504 559708 358556
rect 515588 358436 515640 358488
rect 561128 358436 561180 358488
rect 513196 357688 513248 357740
rect 517888 357688 517940 357740
rect 513288 356328 513340 356380
rect 519084 356328 519136 356380
rect 512276 355376 512328 355428
rect 515128 355376 515180 355428
rect 513288 354968 513340 355020
rect 520556 354968 520608 355020
rect 513288 354696 513340 354748
rect 517980 354696 518032 354748
rect 512828 353472 512880 353524
rect 516324 353472 516376 353524
rect 512460 353336 512512 353388
rect 515220 353336 515272 353388
rect 513012 352656 513064 352708
rect 516600 352656 516652 352708
rect 512460 351976 512512 352028
rect 515036 351976 515088 352028
rect 394700 351908 394752 351960
rect 447140 351908 447192 351960
rect 513288 350888 513340 350940
rect 518072 350888 518124 350940
rect 512460 350752 512512 350804
rect 513932 350752 513984 350804
rect 405740 350548 405792 350600
rect 447140 350548 447192 350600
rect 512828 349800 512880 349852
rect 516508 349800 516560 349852
rect 512460 349256 512512 349308
rect 513840 349256 513892 349308
rect 512552 349188 512604 349240
rect 515312 349188 515364 349240
rect 446956 349052 447008 349104
rect 447784 349052 447836 349104
rect 412640 348372 412692 348424
rect 435640 348372 435692 348424
rect 513288 347896 513340 347948
rect 519176 347896 519228 347948
rect 361764 347760 361816 347812
rect 389824 347760 389876 347812
rect 513104 347760 513156 347812
rect 516692 347760 516744 347812
rect 362316 347692 362368 347744
rect 447140 347692 447192 347744
rect 513288 345176 513340 345228
rect 520648 345176 520700 345228
rect 432696 344292 432748 344344
rect 442264 344292 442316 344344
rect 513288 344224 513340 344276
rect 518164 344224 518216 344276
rect 513288 343816 513340 343868
rect 520740 343816 520792 343868
rect 445576 343068 445628 343120
rect 449716 343068 449768 343120
rect 401600 342864 401652 342916
rect 445576 342864 445628 342916
rect 512460 342524 512512 342576
rect 515588 342524 515640 342576
rect 513288 342252 513340 342304
rect 521660 342252 521712 342304
rect 513288 341232 513340 341284
rect 519268 341232 519320 341284
rect 513104 341096 513156 341148
rect 516876 341096 516928 341148
rect 442908 340960 442960 341012
rect 447232 340960 447284 341012
rect 361764 340892 361816 340944
rect 447140 340892 447192 340944
rect 513288 339600 513340 339652
rect 520832 339600 520884 339652
rect 443736 339532 443788 339584
rect 447232 339532 447284 339584
rect 399484 339464 399536 339516
rect 447140 339464 447192 339516
rect 513288 339464 513340 339516
rect 518256 339464 518308 339516
rect 513288 338240 513340 338292
rect 519728 338240 519780 338292
rect 431224 338172 431276 338224
rect 447140 338172 447192 338224
rect 385960 338104 386012 338156
rect 447232 338104 447284 338156
rect 513012 338104 513064 338156
rect 521752 338104 521804 338156
rect 513012 337152 513064 337204
rect 516968 337152 517020 337204
rect 416780 336880 416832 336932
rect 429936 336880 429988 336932
rect 513288 336880 513340 336932
rect 520924 336880 520976 336932
rect 424140 336812 424192 336864
rect 431408 336812 431460 336864
rect 440976 336812 441028 336864
rect 447140 336812 447192 336864
rect 420460 336744 420512 336796
rect 435732 336744 435784 336796
rect 439596 336744 439648 336796
rect 447232 336744 447284 336796
rect 513104 336744 513156 336796
rect 523132 336744 523184 336796
rect 416228 336336 416280 336388
rect 438216 336336 438268 336388
rect 419448 336268 419500 336320
rect 443828 336268 443880 336320
rect 416044 336200 416096 336252
rect 441160 336200 441212 336252
rect 419356 336132 419408 336184
rect 446956 336132 447008 336184
rect 397460 336064 397512 336116
rect 449072 336064 449124 336116
rect 513288 336064 513340 336116
rect 518348 336064 518400 336116
rect 362224 335996 362276 336048
rect 442908 335996 442960 336048
rect 442264 335452 442316 335504
rect 447324 335452 447376 335504
rect 409420 335384 409472 335436
rect 431316 335384 431368 335436
rect 435456 335384 435508 335436
rect 447232 335384 447284 335436
rect 413100 335316 413152 335368
rect 439780 335316 439832 335368
rect 513288 335316 513340 335368
rect 521844 335316 521896 335368
rect 420184 335044 420236 335096
rect 442540 335044 442592 335096
rect 418804 334976 418856 335028
rect 443920 334976 443972 335028
rect 416136 334908 416188 334960
rect 444012 334908 444064 334960
rect 418896 334840 418948 334892
rect 447048 334840 447100 334892
rect 419264 334772 419316 334824
rect 448980 334772 449032 334824
rect 419080 334704 419132 334756
rect 449532 334704 449584 334756
rect 418988 334636 419040 334688
rect 449440 334636 449492 334688
rect 419172 334568 419224 334620
rect 450728 334568 450780 334620
rect 512460 334500 512512 334552
rect 514116 334500 514168 334552
rect 428096 334364 428148 334416
rect 438124 334228 438176 334280
rect 440240 334228 440292 334280
rect 512828 334160 512880 334212
rect 519452 334160 519504 334212
rect 448244 334092 448296 334144
rect 443644 334024 443696 334076
rect 447324 334024 447376 334076
rect 364064 333956 364116 334008
rect 447232 333956 447284 334008
rect 509240 333956 509292 334008
rect 509700 333956 509752 334008
rect 511356 333208 511408 333260
rect 580264 333208 580316 333260
rect 439504 332664 439556 332716
rect 447324 332664 447376 332716
rect 513288 332664 513340 332716
rect 519636 332664 519688 332716
rect 429844 332596 429896 332648
rect 447232 332596 447284 332648
rect 440240 332528 440292 332580
rect 442632 332528 442684 332580
rect 512828 331440 512880 331492
rect 519360 331440 519412 331492
rect 432880 331304 432932 331356
rect 439688 331304 439740 331356
rect 440884 331304 440936 331356
rect 447232 331304 447284 331356
rect 436744 331236 436796 331288
rect 447600 331236 447652 331288
rect 444196 330556 444248 330608
rect 445760 330556 445812 330608
rect 447232 330556 447284 330608
rect 432604 330488 432656 330540
rect 442356 330488 442408 330540
rect 442908 330080 442960 330132
rect 445852 330080 445904 330132
rect 447232 330080 447284 330132
rect 438768 329740 438820 329792
rect 444104 329740 444156 329792
rect 447232 329740 447284 329792
rect 432420 329672 432472 329724
rect 436928 329672 436980 329724
rect 435364 329060 435416 329112
rect 447232 329060 447284 329112
rect 432788 328856 432840 328908
rect 435548 328856 435600 328908
rect 431868 327700 431920 327752
rect 447232 327700 447284 327752
rect 435732 327020 435784 327072
rect 447232 327020 447284 327072
rect 447876 327020 447928 327072
rect 431408 326340 431460 326392
rect 441620 326340 441672 326392
rect 448152 326340 448204 326392
rect 429936 325592 429988 325644
rect 447784 325592 447836 325644
rect 448060 325592 448112 325644
rect 439780 325524 439832 325576
rect 447968 325524 448020 325576
rect 431316 323552 431368 323604
rect 447324 323552 447376 323604
rect 512920 322940 512972 322992
rect 519544 322940 519596 322992
rect 442632 322872 442684 322924
rect 449900 322872 449952 322924
rect 514024 322464 514076 322516
rect 514300 322464 514352 322516
rect 510528 322396 510580 322448
rect 580632 322396 580684 322448
rect 510068 322328 510120 322380
rect 580540 322328 580592 322380
rect 514024 322260 514076 322312
rect 580356 322260 580408 322312
rect 509148 322192 509200 322244
rect 580172 322192 580224 322244
rect 507216 321852 507268 321904
rect 509240 321852 509292 321904
rect 444012 321784 444064 321836
rect 462136 321784 462188 321836
rect 507584 321784 507636 321836
rect 509884 321784 509936 321836
rect 450728 321716 450780 321768
rect 482560 321716 482612 321768
rect 507952 321716 508004 321768
rect 510068 321716 510120 321768
rect 448980 321648 449032 321700
rect 472348 321648 472400 321700
rect 507860 321648 507912 321700
rect 514024 321648 514076 321700
rect 442540 321580 442592 321632
rect 482284 321580 482336 321632
rect 456616 321512 456668 321564
rect 580908 321512 580960 321564
rect 456340 321444 456392 321496
rect 580080 321444 580132 321496
rect 457996 321376 458048 321428
rect 580448 321376 580500 321428
rect 449164 321308 449216 321360
rect 459376 321308 459428 321360
rect 466828 321308 466880 321360
rect 569500 321308 569552 321360
rect 445024 321240 445076 321292
rect 459100 321240 459152 321292
rect 468208 321240 468260 321292
rect 567844 321240 567896 321292
rect 445116 321172 445168 321224
rect 458824 321172 458876 321224
rect 477592 321172 477644 321224
rect 569408 321172 569460 321224
rect 449256 321104 449308 321156
rect 460480 321104 460532 321156
rect 467656 321104 467708 321156
rect 515404 321104 515456 321156
rect 445208 321036 445260 321088
rect 460204 321036 460256 321088
rect 467380 321036 467432 321088
rect 511264 321036 511316 321088
rect 449072 320968 449124 321020
rect 479800 320968 479852 321020
rect 445668 320900 445720 320952
rect 469036 320900 469088 320952
rect 507400 320900 507452 320952
rect 513380 320900 513432 320952
rect 449900 320832 449952 320884
rect 469220 320832 469272 320884
rect 506940 320832 506992 320884
rect 516784 320832 516836 320884
rect 446496 320764 446548 320816
rect 480076 320764 480128 320816
rect 447048 320696 447100 320748
rect 482836 320696 482888 320748
rect 446404 320628 446456 320680
rect 469864 320628 469916 320680
rect 507032 320492 507084 320544
rect 509976 320492 510028 320544
rect 444288 320084 444340 320136
rect 458548 320084 458600 320136
rect 469220 320084 469272 320136
rect 472624 320084 472676 320136
rect 477040 320084 477092 320136
rect 509148 320084 509200 320136
rect 445392 320016 445444 320068
rect 461032 320016 461084 320068
rect 467104 320016 467156 320068
rect 580816 320016 580868 320068
rect 449532 319948 449584 320000
rect 461860 319948 461912 320000
rect 477868 319948 477920 320000
rect 569316 319948 569368 320000
rect 443920 319880 443972 319932
rect 461584 319880 461636 319932
rect 478696 319880 478748 319932
rect 569224 319880 569276 319932
rect 442448 319812 442500 319864
rect 471796 319812 471848 319864
rect 478420 319812 478472 319864
rect 567936 319812 567988 319864
rect 468760 319744 468812 319796
rect 515496 319744 515548 319796
rect 467932 319676 467984 319728
rect 507952 319676 508004 319728
rect 468484 319608 468536 319660
rect 507860 319608 507912 319660
rect 446680 319540 446732 319592
rect 469588 319540 469640 319592
rect 477316 319540 477368 319592
rect 514300 319540 514352 319592
rect 435640 319472 435692 319524
rect 469128 319472 469180 319524
rect 469220 319472 469272 319524
rect 472900 319472 472952 319524
rect 478972 319472 479024 319524
rect 511356 319472 511408 319524
rect 460204 319404 460256 319456
rect 474556 319404 474608 319456
rect 480812 319404 480864 319456
rect 483112 319404 483164 319456
rect 502156 319404 502208 319456
rect 543740 319404 543792 319456
rect 445300 319336 445352 319388
rect 471520 319336 471572 319388
rect 478144 319336 478196 319388
rect 510528 319336 510580 319388
rect 457168 319268 457220 319320
rect 580724 319268 580776 319320
rect 446864 319200 446916 319252
rect 480352 319200 480404 319252
rect 450544 319132 450596 319184
rect 482008 319132 482060 319184
rect 450636 319064 450688 319116
rect 479524 319064 479576 319116
rect 446588 318996 446640 319048
rect 470140 318996 470192 319048
rect 454316 318928 454368 318980
rect 454684 318928 454736 318980
rect 456892 318724 456944 318776
rect 578884 318724 578936 318776
rect 457444 318656 457496 318708
rect 577504 318656 577556 318708
rect 457720 318588 457772 318640
rect 571984 318588 572036 318640
rect 438216 318520 438268 318572
rect 470692 318520 470744 318572
rect 441160 318452 441212 318504
rect 470416 318452 470468 318504
rect 449440 318384 449492 318436
rect 472072 318384 472124 318436
rect 458824 318112 458876 318164
rect 486976 318112 487028 318164
rect 457444 318044 457496 318096
rect 489184 318044 489236 318096
rect 494428 318044 494480 318096
rect 540980 318044 541032 318096
rect 443828 317364 443880 317416
rect 481732 317364 481784 317416
rect 446956 317296 447008 317348
rect 481180 317296 481232 317348
rect 480260 317228 480312 317280
rect 483388 317228 483440 317280
rect 467104 317160 467156 317212
rect 469220 317160 469272 317212
rect 473452 317160 473504 317212
rect 473912 317160 473964 317212
rect 501604 317024 501656 317076
rect 539140 317024 539192 317076
rect 499672 316956 499724 317008
rect 542452 316956 542504 317008
rect 472624 316888 472676 316940
rect 480812 316888 480864 316940
rect 497188 316888 497240 316940
rect 541072 316888 541124 316940
rect 459008 316820 459060 316872
rect 492220 316820 492272 316872
rect 496084 316820 496136 316872
rect 543188 316820 543240 316872
rect 454776 316752 454828 316804
rect 502432 316752 502484 316804
rect 456064 316684 456116 316736
rect 461584 316684 461636 316736
rect 454684 316616 454736 316668
rect 502984 316684 503036 316736
rect 361764 315936 361816 315988
rect 399484 315936 399536 315988
rect 447784 315528 447836 315580
rect 456892 315528 456944 315580
rect 501052 315528 501104 315580
rect 542728 315528 542780 315580
rect 453396 315460 453448 315512
rect 494152 315460 494204 315512
rect 498292 315460 498344 315512
rect 541164 315460 541216 315512
rect 450636 315392 450688 315444
rect 504088 315392 504140 315444
rect 450544 315324 450596 315376
rect 503812 315324 503864 315376
rect 455512 315256 455564 315308
rect 570604 315256 570656 315308
rect 457628 314644 457680 314696
rect 462412 314644 462464 314696
rect 433248 314508 433300 314560
rect 441068 314508 441120 314560
rect 451924 313964 451976 314016
rect 487252 313964 487304 314016
rect 496636 313964 496688 314016
rect 539600 313964 539652 314016
rect 485596 313896 485648 313948
rect 529940 313896 529992 313948
rect 466552 313216 466604 313268
rect 580172 313216 580224 313268
rect 465172 312536 465224 312588
rect 551284 312536 551336 312588
rect 478144 312400 478196 312452
rect 480260 312400 480312 312452
rect 452108 311176 452160 311228
rect 492772 311176 492824 311228
rect 475384 311108 475436 311160
rect 544384 311108 544436 311160
rect 453304 309816 453356 309868
rect 488356 309816 488408 309868
rect 475108 309748 475160 309800
rect 563704 309748 563756 309800
rect 458916 308456 458968 308508
rect 488632 308456 488684 308508
rect 464620 308388 464672 308440
rect 562324 308388 562376 308440
rect 432236 307708 432288 307760
rect 436836 307708 436888 307760
rect 381636 306280 381688 306332
rect 463516 306280 463568 306332
rect 385868 306212 385920 306264
rect 474280 306212 474332 306264
rect 384580 306144 384632 306196
rect 474004 306144 474056 306196
rect 381728 306076 381780 306128
rect 473728 306076 473780 306128
rect 384764 306008 384816 306060
rect 484768 306008 484820 306060
rect 384856 305940 384908 305992
rect 484492 305940 484544 305992
rect 381544 305872 381596 305924
rect 484216 305872 484268 305924
rect 374644 305804 374696 305856
rect 485320 305804 485372 305856
rect 426348 305736 426400 305788
rect 441620 305736 441672 305788
rect 454224 305736 454276 305788
rect 565084 305736 565136 305788
rect 360936 305668 360988 305720
rect 512184 305668 512236 305720
rect 359464 305600 359516 305652
rect 512552 305600 512604 305652
rect 384396 305532 384448 305584
rect 464068 305532 464120 305584
rect 385776 305464 385828 305516
rect 463792 305464 463844 305516
rect 457536 305396 457588 305448
rect 490012 305396 490064 305448
rect 3424 304988 3476 305040
rect 4804 304988 4856 305040
rect 361764 304920 361816 304972
rect 443736 304920 443788 304972
rect 455788 304444 455840 304496
rect 573364 304444 573416 304496
rect 385684 304376 385736 304428
rect 519728 304376 519780 304428
rect 361028 304308 361080 304360
rect 512828 304308 512880 304360
rect 359556 304240 359608 304292
rect 512368 304240 512420 304292
rect 378692 303560 378744 303612
rect 483940 303560 483992 303612
rect 485872 303560 485924 303612
rect 530032 303560 530084 303612
rect 382004 303492 382056 303544
rect 511448 303492 511500 303544
rect 379060 303424 379112 303476
rect 509516 303424 509568 303476
rect 376024 303356 376076 303408
rect 506940 303356 506992 303408
rect 379244 303288 379296 303340
rect 511080 303288 511132 303340
rect 382096 303220 382148 303272
rect 515312 303220 515364 303272
rect 376208 303152 376260 303204
rect 509424 303152 509476 303204
rect 379336 303084 379388 303136
rect 513932 303084 513984 303136
rect 379152 303016 379204 303068
rect 515128 303016 515180 303068
rect 378968 302948 379020 303000
rect 515220 302948 515272 303000
rect 373264 302880 373316 302932
rect 513564 302880 513616 302932
rect 379428 302812 379480 302864
rect 473912 302812 473964 302864
rect 381452 302744 381504 302796
rect 463240 302744 463292 302796
rect 386144 302676 386196 302728
rect 462964 302676 463016 302728
rect 486424 301588 486476 301640
rect 529204 301588 529256 301640
rect 378784 301520 378836 301572
rect 464344 301520 464396 301572
rect 465724 301520 465776 301572
rect 537484 301520 537536 301572
rect 407120 301452 407172 301504
rect 502708 301452 502760 301504
rect 376300 300772 376352 300824
rect 510988 300772 511040 300824
rect 373632 300704 373684 300756
rect 511540 300704 511592 300756
rect 376392 300636 376444 300688
rect 513748 300636 513800 300688
rect 368296 300568 368348 300620
rect 507032 300568 507084 300620
rect 373540 300500 373592 300552
rect 513472 300500 513524 300552
rect 373448 300432 373500 300484
rect 514944 300432 514996 300484
rect 370872 300364 370924 300416
rect 514852 300364 514904 300416
rect 371056 300296 371108 300348
rect 516140 300296 516192 300348
rect 370964 300228 371016 300280
rect 517704 300228 517756 300280
rect 370780 300160 370832 300212
rect 517520 300160 517572 300212
rect 368112 300092 368164 300144
rect 518348 300092 518400 300144
rect 376484 300024 376536 300076
rect 509332 300024 509384 300076
rect 378600 299956 378652 300008
rect 483664 299956 483716 300008
rect 376668 299888 376720 299940
rect 473176 299888 473228 299940
rect 461584 299412 461636 299464
rect 580172 299412 580224 299464
rect 376576 298800 376628 298852
rect 485044 298800 485096 298852
rect 371976 298732 372028 298784
rect 513196 298732 513248 298784
rect 365168 298052 365220 298104
rect 507584 298052 507636 298104
rect 367836 297984 367888 298036
rect 514116 297984 514168 298036
rect 363604 297916 363656 297968
rect 512276 297916 512328 297968
rect 367928 297848 367980 297900
rect 516968 297848 517020 297900
rect 365076 297780 365128 297832
rect 515588 297780 515640 297832
rect 361212 297712 361264 297764
rect 512092 297712 512144 297764
rect 365536 297644 365588 297696
rect 516876 297644 516928 297696
rect 365260 297576 365312 297628
rect 516692 297576 516744 297628
rect 362316 297508 362368 297560
rect 513840 297508 513892 297560
rect 365444 297440 365496 297492
rect 518256 297440 518308 297492
rect 362224 297372 362276 297424
rect 518072 297372 518124 297424
rect 365352 297304 365404 297356
rect 507768 297304 507820 297356
rect 382924 297236 382976 297288
rect 518164 297236 518216 297288
rect 464344 297168 464396 297220
rect 467104 297168 467156 297220
rect 476212 297168 476264 297220
rect 548524 297168 548576 297220
rect 454408 295944 454460 295996
rect 578884 295944 578936 295996
rect 369216 295264 369268 295316
rect 514760 295264 514812 295316
rect 366640 295196 366692 295248
rect 514208 295196 514260 295248
rect 369124 295128 369176 295180
rect 516232 295128 516284 295180
rect 366456 295060 366508 295112
rect 513656 295060 513708 295112
rect 361304 294992 361356 295044
rect 510896 294992 510948 295044
rect 369308 294924 369360 294976
rect 518992 294924 519044 294976
rect 366732 294856 366784 294908
rect 517796 294856 517848 294908
rect 363972 294788 364024 294840
rect 516416 294788 516468 294840
rect 363880 294720 363932 294772
rect 517888 294720 517940 294772
rect 362408 294652 362460 294704
rect 516600 294652 516652 294704
rect 362500 294584 362552 294636
rect 517980 294584 518032 294636
rect 366548 294516 366600 294568
rect 510712 294516 510764 294568
rect 368204 294448 368256 294500
rect 509792 294448 509844 294500
rect 454316 294380 454368 294432
rect 576124 294380 576176 294432
rect 361764 293904 361816 293956
rect 385960 293904 386012 293956
rect 459100 293292 459152 293344
rect 488908 293292 488960 293344
rect 475936 293224 475988 293276
rect 536104 293224 536156 293276
rect 3516 292748 3568 292800
rect 4896 292748 4948 292800
rect 375104 292476 375156 292528
rect 507400 292476 507452 292528
rect 381820 292408 381872 292460
rect 519176 292408 519228 292460
rect 380164 292340 380216 292392
rect 520648 292340 520700 292392
rect 380256 292272 380308 292324
rect 520740 292272 520792 292324
rect 377588 292204 377640 292256
rect 519268 292204 519320 292256
rect 377404 292136 377456 292188
rect 520832 292136 520884 292188
rect 375012 292068 375064 292120
rect 519452 292068 519504 292120
rect 374736 292000 374788 292052
rect 519636 292000 519688 292052
rect 374920 291932 374972 291984
rect 520924 291932 520976 291984
rect 372252 291864 372304 291916
rect 518900 291864 518952 291916
rect 372344 291796 372396 291848
rect 520280 291796 520332 291848
rect 377680 291728 377732 291780
rect 507676 291728 507728 291780
rect 454960 291660 455012 291712
rect 574744 291660 574796 291712
rect 455236 290436 455288 290488
rect 533344 290436 533396 290488
rect 383200 289756 383252 289808
rect 516324 289756 516376 289808
rect 386236 289688 386288 289740
rect 520464 289688 520516 289740
rect 380440 289620 380492 289672
rect 515036 289620 515088 289672
rect 383292 289552 383344 289604
rect 519084 289552 519136 289604
rect 380348 289484 380400 289536
rect 516508 289484 516560 289536
rect 383016 289416 383068 289468
rect 519360 289416 519412 289468
rect 383108 289348 383160 289400
rect 520556 289348 520608 289400
rect 378876 289280 378928 289332
rect 517612 289280 517664 289332
rect 363788 289212 363840 289264
rect 507308 289212 507360 289264
rect 373356 289144 373408 289196
rect 520372 289144 520424 289196
rect 370596 289076 370648 289128
rect 523040 289076 523092 289128
rect 385960 289008 386012 289060
rect 507492 289008 507544 289060
rect 386052 288940 386104 288992
rect 507216 288940 507268 288992
rect 446588 288872 446640 288924
rect 464344 288872 464396 288924
rect 474004 288804 474056 288856
rect 478144 288804 478196 288856
rect 466000 287648 466052 287700
rect 569224 287648 569276 287700
rect 452016 286764 452068 286816
rect 487528 286764 487580 286816
rect 456800 286696 456852 286748
rect 504916 286696 504968 286748
rect 439688 286628 439740 286680
rect 446588 286628 446640 286680
rect 475660 286628 475712 286680
rect 571984 286628 572036 286680
rect 377496 286560 377548 286612
rect 507124 286560 507176 286612
rect 384948 286492 385000 286544
rect 521844 286492 521896 286544
rect 374828 286424 374880 286476
rect 521660 286424 521712 286476
rect 372068 286356 372120 286408
rect 521752 286356 521804 286408
rect 369400 286288 369452 286340
rect 523132 286288 523184 286340
rect 460388 285676 460440 285728
rect 462688 285676 462740 285728
rect 453580 285064 453632 285116
rect 493876 285064 493928 285116
rect 464896 284996 464948 285048
rect 547144 284996 547196 285048
rect 363696 284928 363748 284980
rect 474832 284928 474884 284980
rect 486148 284928 486200 284980
rect 531320 284928 531372 284980
rect 452292 283704 452344 283756
rect 493048 283704 493100 283756
rect 501880 283704 501932 283756
rect 539232 283704 539284 283756
rect 449900 283636 449952 283688
rect 504640 283636 504692 283688
rect 446404 283568 446456 283620
rect 457628 283568 457680 283620
rect 476488 283568 476540 283620
rect 566464 283568 566516 283620
rect 361764 282820 361816 282872
rect 431224 282820 431276 282872
rect 471244 282208 471296 282260
rect 474004 282208 474056 282260
rect 456248 282140 456300 282192
rect 492496 282140 492548 282192
rect 459284 280780 459336 280832
rect 491392 280780 491444 280832
rect 459192 279420 459244 279472
rect 490564 279420 490616 279472
rect 452384 277992 452436 278044
rect 493324 277992 493376 278044
rect 498844 277992 498896 278044
rect 541532 277992 541584 278044
rect 460296 276768 460348 276820
rect 489460 276768 489512 276820
rect 498016 276768 498068 276820
rect 539876 276768 539928 276820
rect 457720 276700 457772 276752
rect 491668 276700 491720 276752
rect 496912 276700 496964 276752
rect 539784 276700 539836 276752
rect 359648 276632 359700 276684
rect 512000 276632 512052 276684
rect 497740 275408 497792 275460
rect 541440 275408 541492 275460
rect 457628 275340 457680 275392
rect 490840 275340 490892 275392
rect 495256 275340 495308 275392
rect 541256 275340 541308 275392
rect 453488 275272 453540 275324
rect 488080 275272 488132 275324
rect 495808 275272 495860 275324
rect 542820 275272 542872 275324
rect 456984 274660 457036 274712
rect 460388 274660 460440 274712
rect 499120 274048 499172 274100
rect 540060 274048 540112 274100
rect 456156 273980 456208 274032
rect 490380 273980 490432 274032
rect 497464 273980 497516 274032
rect 541348 273980 541400 274032
rect 453672 273912 453724 273964
rect 493600 273912 493652 273964
rect 495532 273912 495584 273964
rect 542636 273912 542688 273964
rect 476764 273164 476816 273216
rect 580172 273164 580224 273216
rect 456064 272552 456116 272604
rect 489736 272552 489788 272604
rect 498568 272552 498620 272604
rect 539968 272552 540020 272604
rect 454960 272484 455012 272536
rect 491944 272484 491996 272536
rect 496360 272484 496412 272536
rect 542912 272484 542964 272536
rect 361764 271804 361816 271856
rect 439596 271804 439648 271856
rect 501328 271396 501380 271448
rect 540336 271396 540388 271448
rect 456340 271328 456392 271380
rect 491116 271328 491168 271380
rect 494980 271328 495032 271380
rect 539692 271328 539744 271380
rect 436836 271260 436888 271312
rect 439688 271260 439740 271312
rect 454868 271260 454920 271312
rect 504364 271260 504416 271312
rect 450728 271192 450780 271244
rect 503536 271192 503588 271244
rect 466276 271124 466328 271176
rect 580264 271124 580316 271176
rect 500500 270036 500552 270088
rect 540244 270036 540296 270088
rect 455052 269968 455104 270020
rect 486700 269968 486752 270020
rect 499948 269968 500000 270020
rect 543096 269968 543148 270020
rect 450820 269900 450872 269952
rect 503260 269900 503312 269952
rect 465448 269832 465500 269884
rect 554044 269832 554096 269884
rect 445668 269764 445720 269816
rect 510620 269764 510672 269816
rect 443000 269288 443052 269340
rect 446404 269288 446456 269340
rect 447784 268540 447836 268592
rect 456984 268540 457036 268592
rect 453764 268472 453816 268524
rect 472624 268472 472676 268524
rect 500224 268472 500276 268524
rect 540152 268472 540204 268524
rect 450084 268404 450136 268456
rect 471244 268404 471296 268456
rect 499396 268404 499448 268456
rect 543004 268404 543056 268456
rect 452200 268336 452252 268388
rect 487804 268336 487856 268388
rect 494704 268336 494756 268388
rect 542544 268336 542596 268388
rect 449624 263508 449676 263560
rect 456984 263508 457036 263560
rect 440240 262760 440292 262812
rect 443000 262760 443052 262812
rect 445024 262760 445076 262812
rect 450084 262760 450136 262812
rect 361764 260788 361816 260840
rect 440976 260788 441028 260840
rect 431960 260312 432012 260364
rect 440240 260312 440292 260364
rect 429936 254872 429988 254924
rect 431960 254872 432012 254924
rect 3792 253920 3844 253972
rect 4988 253920 5040 253972
rect 442448 252424 442500 252476
rect 447784 252424 447836 252476
rect 361764 249704 361816 249756
rect 435456 249704 435508 249756
rect 442356 249704 442408 249756
rect 445024 249704 445076 249756
rect 449716 249024 449768 249076
rect 458088 249024 458140 249076
rect 573364 245556 573416 245608
rect 580172 245556 580224 245608
rect 439596 244944 439648 244996
rect 442448 244944 442500 244996
rect 3884 241408 3936 241460
rect 5080 241408 5132 241460
rect 361764 238688 361816 238740
rect 442264 238688 442316 238740
rect 419448 233860 419500 233912
rect 456708 233860 456760 233912
rect 566464 233180 566516 233232
rect 579988 233180 580040 233232
rect 448244 232568 448296 232620
rect 454040 232568 454092 232620
rect 428464 232500 428516 232552
rect 453764 232500 453816 232552
rect 433984 230936 434036 230988
rect 439596 230936 439648 230988
rect 424324 227740 424376 227792
rect 429936 227740 429988 227792
rect 361764 227672 361816 227724
rect 443644 227672 443696 227724
rect 416044 221416 416096 221468
rect 454040 221416 454092 221468
rect 457904 221416 457956 221468
rect 569224 219376 569276 219428
rect 580172 219376 580224 219428
rect 427820 217540 427872 217592
rect 433984 217540 434036 217592
rect 423036 216656 423088 216708
rect 428464 216656 428516 216708
rect 361672 216316 361724 216368
rect 364064 216316 364116 216368
rect 3976 214752 4028 214804
rect 5172 214752 5224 214804
rect 422944 213120 422996 213172
rect 427820 213120 427872 213172
rect 434260 212984 434312 213036
rect 436836 212984 436888 213036
rect 406384 211760 406436 211812
rect 423036 211760 423088 211812
rect 420184 209788 420236 209840
rect 424324 209788 424376 209840
rect 428464 209788 428516 209840
rect 434260 209788 434312 209840
rect 570604 206932 570656 206984
rect 579804 206932 579856 206984
rect 411260 206252 411312 206304
rect 448336 206252 448388 206304
rect 456708 206252 456760 206304
rect 361764 205572 361816 205624
rect 439504 205572 439556 205624
rect 433248 203532 433300 203584
rect 442356 203532 442408 203584
rect 419540 201492 419592 201544
rect 422944 201492 422996 201544
rect 417424 200744 417476 200796
rect 433248 200744 433300 200796
rect 459468 200744 459520 200796
rect 485780 200744 485832 200796
rect 458088 200132 458140 200184
rect 462964 200132 463016 200184
rect 459376 199384 459428 199436
rect 481640 199384 481692 199436
rect 398104 196664 398156 196716
rect 419540 196664 419592 196716
rect 367744 196596 367796 196648
rect 406384 196596 406436 196648
rect 448428 196596 448480 196648
rect 461584 196596 461636 196648
rect 449992 195236 450044 195288
rect 528560 195236 528612 195288
rect 416136 194692 416188 194744
rect 420184 194692 420236 194744
rect 361764 194488 361816 194540
rect 429844 194488 429896 194540
rect 392584 193808 392636 193860
rect 398104 193808 398156 193860
rect 548524 193128 548576 193180
rect 580172 193128 580224 193180
rect 405004 189728 405056 189780
rect 416136 189728 416188 189780
rect 361764 183472 361816 183524
rect 436744 183472 436796 183524
rect 389916 182112 389968 182164
rect 392584 182112 392636 182164
rect 361580 180072 361632 180124
rect 417424 180072 417476 180124
rect 537484 179324 537536 179376
rect 580172 179324 580224 179376
rect 401600 172524 401652 172576
rect 405004 172524 405056 172576
rect 361764 171776 361816 171828
rect 440884 171776 440936 171828
rect 524420 171776 524472 171828
rect 397460 169736 397512 169788
rect 401600 169736 401652 169788
rect 362684 167628 362736 167680
rect 389916 167628 389968 167680
rect 533344 166948 533396 167000
rect 580172 166948 580224 167000
rect 390560 164840 390612 164892
rect 397460 164840 397512 164892
rect 414756 163888 414808 163940
rect 416044 163888 416096 163940
rect 434904 162800 434956 162852
rect 435364 162800 435416 162852
rect 365720 162188 365772 162240
rect 390560 162188 390612 162240
rect 389824 162120 389876 162172
rect 444932 162120 444984 162172
rect 425060 161848 425112 161900
rect 426348 161848 426400 161900
rect 496820 161848 496872 161900
rect 428648 161780 428700 161832
rect 500960 161780 501012 161832
rect 421748 161712 421800 161764
rect 494060 161712 494112 161764
rect 410524 161644 410576 161696
rect 425060 161644 425112 161696
rect 431868 161644 431920 161696
rect 505100 161644 505152 161696
rect 407764 161576 407816 161628
rect 434904 161576 434956 161628
rect 438768 161576 438820 161628
rect 513380 161576 513432 161628
rect 403624 161508 403676 161560
rect 442908 161508 442960 161560
rect 517520 161508 517572 161560
rect 362592 161440 362644 161492
rect 441620 161440 441672 161492
rect 444932 161440 444984 161492
rect 445668 161440 445720 161492
rect 532700 161440 532752 161492
rect 361764 161372 361816 161424
rect 444196 161372 444248 161424
rect 359832 160692 359884 160744
rect 367744 160692 367796 160744
rect 420920 160692 420972 160744
rect 428464 160692 428516 160744
rect 444196 160692 444248 160744
rect 521660 160692 521712 160744
rect 410616 160352 410668 160404
rect 428004 160352 428056 160404
rect 406384 160284 406436 160336
rect 431316 160284 431368 160336
rect 386328 160216 386380 160268
rect 414756 160216 414808 160268
rect 381360 160148 381412 160200
rect 421380 160148 421432 160200
rect 421748 160148 421800 160200
rect 434904 160148 434956 160200
rect 435272 160148 435324 160200
rect 450912 160148 450964 160200
rect 359740 160080 359792 160132
rect 362684 160080 362736 160132
rect 383384 160080 383436 160132
rect 418390 160080 418442 160132
rect 419448 160080 419500 160132
rect 461676 160080 461728 160132
rect 407396 159400 407448 159452
rect 420920 159468 420972 159520
rect 449808 159332 449860 159384
rect 536840 159332 536892 159384
rect 452568 158380 452620 158432
rect 455052 158380 455104 158432
rect 452384 157292 452436 157344
rect 453396 157292 453448 157344
rect 405648 156068 405700 156120
rect 407396 156068 407448 156120
rect 359924 155864 359976 155916
rect 365720 155864 365772 155916
rect 452384 155796 452436 155848
rect 453580 155796 453632 155848
rect 452384 154300 452436 154352
rect 453672 154300 453724 154352
rect 402336 153212 402388 153264
rect 405648 153212 405700 153264
rect 536104 153144 536156 153196
rect 580172 153144 580224 153196
rect 452568 148996 452620 149048
rect 456248 148996 456300 149048
rect 399484 147636 399536 147688
rect 402336 147636 402388 147688
rect 452568 147500 452620 147552
rect 459008 147500 459060 147552
rect 452568 146140 452620 146192
rect 454960 146140 455012 146192
rect 452568 144780 452620 144832
rect 457720 144780 457772 144832
rect 452568 143420 452620 143472
rect 459284 143420 459336 143472
rect 461676 142876 461728 142928
rect 489920 142876 489972 142928
rect 450912 142808 450964 142860
rect 509608 142808 509660 142860
rect 452568 142060 452620 142112
rect 456340 142060 456392 142112
rect 464344 140768 464396 140820
rect 481640 140768 481692 140820
rect 452568 140700 452620 140752
rect 457628 140700 457680 140752
rect 388444 140020 388496 140072
rect 399484 140020 399536 140072
rect 361764 139340 361816 139392
rect 403624 139340 403676 139392
rect 452568 139340 452620 139392
rect 459192 139340 459244 139392
rect 554044 139340 554096 139392
rect 580172 139340 580224 139392
rect 452568 137844 452620 137896
rect 456156 137844 456208 137896
rect 451556 136484 451608 136536
rect 457536 136484 457588 136536
rect 452568 135124 452620 135176
rect 456064 135124 456116 135176
rect 452568 133764 452620 133816
rect 460296 133764 460348 133816
rect 452568 132404 452620 132456
rect 457444 132404 457496 132456
rect 452568 131044 452620 131096
rect 459100 131044 459152 131096
rect 452568 129684 452620 129736
rect 458916 129684 458968 129736
rect 361764 128256 361816 128308
rect 407764 128256 407816 128308
rect 452292 128256 452344 128308
rect 453304 128256 453356 128308
rect 452384 126896 452436 126948
rect 453488 126896 453540 126948
rect 574744 126896 574796 126948
rect 580172 126896 580224 126948
rect 362592 124856 362644 124908
rect 388444 124856 388496 124908
rect 451924 122136 451976 122188
rect 458824 122136 458876 122188
rect 361764 117240 361816 117292
rect 406384 117240 406436 117292
rect 571984 113092 572036 113144
rect 579804 113092 579856 113144
rect 445300 107312 445352 107364
rect 454868 107312 454920 107364
rect 439136 107244 439188 107296
rect 450636 107244 450688 107296
rect 432972 107176 433024 107228
rect 450544 107176 450596 107228
rect 426808 107108 426860 107160
rect 450728 107108 450780 107160
rect 420644 107040 420696 107092
rect 450820 107040 450872 107092
rect 414480 106972 414532 107024
rect 454684 106972 454736 107024
rect 402152 106904 402204 106956
rect 454776 106904 454828 106956
rect 367744 106292 367796 106344
rect 389824 106292 389876 106344
rect 361764 106224 361816 106276
rect 410616 106224 410668 106276
rect 362684 105544 362736 105596
rect 410524 105544 410576 105596
rect 551284 100648 551336 100700
rect 580172 100648 580224 100700
rect 3700 98608 3752 98660
rect 19984 98608 20036 98660
rect 4896 97996 4948 98048
rect 8944 97928 8996 97980
rect 576124 86912 576176 86964
rect 580172 86912 580224 86964
rect 3148 84192 3200 84244
rect 20904 84192 20956 84244
rect 361764 84124 361816 84176
rect 381360 84124 381412 84176
rect 361764 73108 361816 73160
rect 383384 73108 383436 73160
rect 544384 73108 544436 73160
rect 580172 73108 580224 73160
rect 4988 71204 5040 71256
rect 6184 71204 6236 71256
rect 3148 70388 3200 70440
rect 20076 70388 20128 70440
rect 8944 67532 8996 67584
rect 10968 67532 11020 67584
rect 462504 67532 462556 67584
rect 464344 67532 464396 67584
rect 4804 66852 4856 66904
rect 7288 66852 7340 66904
rect 7288 63656 7340 63708
rect 9680 63656 9732 63708
rect 361764 62024 361816 62076
rect 386328 62024 386380 62076
rect 5080 60664 5132 60716
rect 6000 60664 6052 60716
rect 547144 60664 547196 60716
rect 580172 60664 580224 60716
rect 11060 59372 11112 59424
rect 13820 59304 13872 59356
rect 6000 58624 6052 58676
rect 11704 58624 11756 58676
rect 5172 57196 5224 57248
rect 8208 57196 8260 57248
rect 13820 56516 13872 56568
rect 16488 56516 16540 56568
rect 9680 55224 9732 55276
rect 13728 55156 13780 55208
rect 6184 53796 6236 53848
rect 8392 53728 8444 53780
rect 11704 53388 11756 53440
rect 13728 53388 13780 53440
rect 8208 52436 8260 52488
rect 11060 52368 11112 52420
rect 8392 51688 8444 51740
rect 19248 51688 19300 51740
rect 13728 51076 13780 51128
rect 361764 51076 361816 51128
rect 384212 51076 384264 51128
rect 540612 51076 540664 51128
rect 543740 51076 543792 51128
rect 17868 51008 17920 51060
rect 13820 50940 13872 50992
rect 18604 50940 18656 50992
rect 16580 50124 16632 50176
rect 19340 50124 19392 50176
rect 11060 49716 11112 49768
rect 18236 49648 18288 49700
rect 18604 48288 18656 48340
rect 20904 48220 20956 48272
rect 17868 48152 17920 48204
rect 20720 48152 20772 48204
rect 18236 47880 18288 47932
rect 20812 47880 20864 47932
rect 19340 46996 19392 47048
rect 21272 46996 21324 47048
rect 3516 46860 3568 46912
rect 386144 46860 386196 46912
rect 3700 46792 3752 46844
rect 385868 46792 385920 46844
rect 3240 46724 3292 46776
rect 384580 46724 384632 46776
rect 3332 46656 3384 46708
rect 381636 46656 381688 46708
rect 3976 46588 4028 46640
rect 381728 46588 381780 46640
rect 3884 46520 3936 46572
rect 381452 46520 381504 46572
rect 3608 46452 3660 46504
rect 379428 46452 379480 46504
rect 3792 46384 3844 46436
rect 378692 46384 378744 46436
rect 20076 46316 20128 46368
rect 384396 46316 384448 46368
rect 19984 46248 20036 46300
rect 376668 46248 376720 46300
rect 20812 46180 20864 46232
rect 359924 46180 359976 46232
rect 20720 46112 20772 46164
rect 359832 46112 359884 46164
rect 21272 46044 21324 46096
rect 359740 46044 359792 46096
rect 358176 45772 358228 45824
rect 362592 45772 362644 45824
rect 4068 45568 4120 45620
rect 381544 45500 381596 45552
rect 3516 45432 3568 45484
rect 376576 45432 376628 45484
rect 20904 45364 20956 45416
rect 358176 45364 358228 45416
rect 71780 45296 71832 45348
rect 378968 45296 379020 45348
rect 69020 45228 69072 45280
rect 379244 45228 379296 45280
rect 64880 45160 64932 45212
rect 379336 45160 379388 45212
rect 60740 45092 60792 45144
rect 382096 45092 382148 45144
rect 57980 45024 58032 45076
rect 382004 45024 382056 45076
rect 53840 44956 53892 45008
rect 381912 44956 381964 45008
rect 51080 44888 51132 44940
rect 382188 44888 382240 44940
rect 6920 44820 6972 44872
rect 384672 44820 384724 44872
rect 75920 44752 75972 44804
rect 379152 44752 379204 44804
rect 78680 44684 78732 44736
rect 379060 44684 379112 44736
rect 85580 44616 85632 44668
rect 376484 44616 376536 44668
rect 114560 42712 114612 42764
rect 370964 42712 371016 42764
rect 110420 42644 110472 42696
rect 370872 42644 370924 42696
rect 107660 42576 107712 42628
rect 373264 42576 373316 42628
rect 103520 42508 103572 42560
rect 373448 42508 373500 42560
rect 100760 42440 100812 42492
rect 373540 42440 373592 42492
rect 96620 42372 96672 42424
rect 373632 42372 373684 42424
rect 93860 42304 93912 42356
rect 376392 42304 376444 42356
rect 89720 42236 89772 42288
rect 376300 42236 376352 42288
rect 82820 42168 82872 42220
rect 376208 42168 376260 42220
rect 20720 42100 20772 42152
rect 368296 42100 368348 42152
rect 11060 42032 11112 42084
rect 376116 42032 376168 42084
rect 118700 41964 118752 42016
rect 371056 41964 371108 42016
rect 121460 41896 121512 41948
rect 370780 41896 370832 41948
rect 461584 41352 461636 41404
rect 536840 41352 536892 41404
rect 77300 39992 77352 40044
rect 361304 39992 361356 40044
rect 73160 39924 73212 39976
rect 362500 39924 362552 39976
rect 69112 39856 69164 39908
rect 362408 39856 362460 39908
rect 66260 39788 66312 39840
rect 362224 39788 362276 39840
rect 62120 39720 62172 39772
rect 362316 39720 362368 39772
rect 59360 39652 59412 39704
rect 365260 39652 365312 39704
rect 44180 39584 44232 39636
rect 365536 39584 365588 39636
rect 40040 39516 40092 39568
rect 365444 39516 365496 39568
rect 33140 39448 33192 39500
rect 368112 39448 368164 39500
rect 26240 39380 26292 39432
rect 368020 39380 368072 39432
rect 2780 39312 2832 39364
rect 365352 39312 365404 39364
rect 80060 39244 80112 39296
rect 363880 39244 363932 39296
rect 84200 39176 84252 39228
rect 363972 39176 364024 39228
rect 115940 37204 115992 37256
rect 372252 37204 372304 37256
rect 111800 37136 111852 37188
rect 369308 37136 369360 37188
rect 109040 37068 109092 37120
rect 369216 37068 369268 37120
rect 104900 37000 104952 37052
rect 369124 37000 369176 37052
rect 102140 36932 102192 36984
rect 366640 36932 366692 36984
rect 98000 36864 98052 36916
rect 366732 36864 366784 36916
rect 93952 36796 94004 36848
rect 366548 36796 366600 36848
rect 91100 36728 91152 36780
rect 368204 36728 368256 36780
rect 86960 36660 87012 36712
rect 366456 36660 366508 36712
rect 22100 36592 22152 36644
rect 375104 36592 375156 36644
rect 17960 36524 18012 36576
rect 372160 36524 372212 36576
rect 118792 36456 118844 36508
rect 372344 36456 372396 36508
rect 122840 36388 122892 36440
rect 371884 36388 371936 36440
rect 74540 34416 74592 34468
rect 383108 34416 383160 34468
rect 462964 34416 463016 34468
rect 536840 34416 536892 34468
rect 67640 34348 67692 34400
rect 380440 34348 380492 34400
rect 70400 34280 70452 34332
rect 383200 34280 383252 34332
rect 63500 34212 63552 34264
rect 380348 34212 380400 34264
rect 60832 34144 60884 34196
rect 381820 34144 381872 34196
rect 52460 34076 52512 34128
rect 380164 34076 380216 34128
rect 49700 34008 49752 34060
rect 380256 34008 380308 34060
rect 44272 33940 44324 33992
rect 377588 33940 377640 33992
rect 34520 33872 34572 33924
rect 374920 33872 374972 33924
rect 30380 33804 30432 33856
rect 375012 33804 375064 33856
rect 9680 33736 9732 33788
rect 377680 33736 377732 33788
rect 77392 33668 77444 33720
rect 383292 33668 383344 33720
rect 85672 33600 85724 33652
rect 386236 33600 386288 33652
rect 3516 33056 3568 33108
rect 378784 33056 378836 33108
rect 563704 33056 563756 33108
rect 580172 33056 580224 33108
rect 3424 31696 3476 31748
rect 460204 31696 460256 31748
rect 120080 31628 120132 31680
rect 364984 31628 365036 31680
rect 384212 31628 384264 31680
rect 462320 31628 462372 31680
rect 113180 31560 113232 31612
rect 370596 31560 370648 31612
rect 102232 31492 102284 31544
rect 373356 31492 373408 31544
rect 111064 31424 111116 31476
rect 386052 31424 386104 31476
rect 99380 31356 99432 31408
rect 376024 31356 376076 31408
rect 92480 31288 92532 31340
rect 378876 31288 378928 31340
rect 35900 31220 35952 31272
rect 369400 31220 369452 31272
rect 19340 31152 19392 31204
rect 363788 31152 363840 31204
rect 31760 31084 31812 31136
rect 384948 31084 385000 31136
rect 13820 31016 13872 31068
rect 385960 31016 386012 31068
rect 117320 30948 117372 31000
rect 360844 30948 360896 31000
rect 124220 30880 124272 30932
rect 366364 30880 366416 30932
rect 106924 28364 106976 28416
rect 377496 28364 377548 28416
rect 45560 28296 45612 28348
rect 374828 28296 374880 28348
rect 38660 28228 38712 28280
rect 372068 28228 372120 28280
rect 3424 20612 3476 20664
rect 363696 20612 363748 20664
rect 562324 20612 562376 20664
rect 579988 20612 580040 20664
rect 572 7556 624 7608
rect 367744 7556 367796 7608
rect 3424 6808 3476 6860
rect 374644 6808 374696 6860
rect 565084 6808 565136 6860
rect 580172 6808 580224 6860
rect 89168 4088 89220 4140
rect 363604 4088 363656 4140
rect 82084 4020 82136 4072
rect 359648 4020 359700 4072
rect 56048 3952 56100 4004
rect 359464 3952 359516 4004
rect 57244 3884 57296 3936
rect 371976 3884 372028 3936
rect 48964 3816 49016 3868
rect 365076 3816 365128 3868
rect 43076 3748 43128 3800
rect 361120 3748 361172 3800
rect 52552 3680 52604 3732
rect 382924 3680 382976 3732
rect 37188 3612 37240 3664
rect 367928 3612 367980 3664
rect 41880 3544 41932 3596
rect 377404 3544 377456 3596
rect 27712 3476 27764 3528
rect 374736 3476 374788 3528
rect 38384 3408 38436 3460
rect 385684 3408 385736 3460
rect 60740 3340 60792 3392
rect 61660 3340 61712 3392
rect 85580 3340 85632 3392
rect 86500 3340 86552 3392
rect 96252 3340 96304 3392
rect 359556 3340 359608 3392
rect 110420 3272 110472 3324
rect 111616 3272 111668 3324
rect 6460 3204 6512 3256
rect 106832 3204 106884 3256
rect 28908 3136 28960 3188
rect 106924 3136 106976 3188
rect 361212 3272 361264 3324
rect 111064 3068 111116 3120
rect 110512 3000 110564 3052
rect 360936 3204 360988 3256
rect 30104 2116 30156 2168
rect 367836 2116 367888 2168
rect 2872 2048 2924 2100
rect 384304 2048 384356 2100
<< metal2 >>
rect 6932 703582 7972 703610
rect 3976 684752 4028 684758
rect 3976 684694 4028 684700
rect 3608 684684 3660 684690
rect 3608 684626 3660 684632
rect 3424 684616 3476 684622
rect 3424 684558 3476 684564
rect 3332 684548 3384 684554
rect 3332 684490 3384 684496
rect 3238 684312 3294 684321
rect 3238 684247 3294 684256
rect 3252 683194 3280 684247
rect 3240 683188 3292 683194
rect 3240 683130 3292 683136
rect 3054 682816 3110 682825
rect 3054 682751 3110 682760
rect 3068 673454 3096 682751
rect 3148 682712 3200 682718
rect 3148 682654 3200 682660
rect 3160 678042 3188 682654
rect 3344 678994 3372 684490
rect 3436 679130 3464 684558
rect 3516 683392 3568 683398
rect 3516 683334 3568 683340
rect 3528 679250 3556 683334
rect 3620 679266 3648 684626
rect 3884 683460 3936 683466
rect 3884 683402 3936 683408
rect 3792 683256 3844 683262
rect 3792 683198 3844 683204
rect 3516 679244 3568 679250
rect 3620 679238 3740 679266
rect 3516 679186 3568 679192
rect 3436 679102 3648 679130
rect 3516 679040 3568 679046
rect 3344 678966 3464 678994
rect 3516 678982 3568 678988
rect 3160 678014 3372 678042
rect 3068 673426 3280 673454
rect 3148 658232 3200 658238
rect 3146 658200 3148 658209
rect 3200 658200 3202 658209
rect 3146 658135 3202 658144
rect 3252 580009 3280 673426
rect 3238 580000 3294 580009
rect 3238 579935 3294 579944
rect 3344 566953 3372 678014
rect 3330 566944 3386 566953
rect 3330 566879 3386 566888
rect 3436 449585 3464 678966
rect 3528 462641 3556 678982
rect 3620 475697 3648 679102
rect 3712 678570 3740 679238
rect 3700 678564 3752 678570
rect 3700 678506 3752 678512
rect 3804 678450 3832 683198
rect 3712 678422 3832 678450
rect 3712 632097 3740 678422
rect 3896 678314 3924 683402
rect 3804 678286 3924 678314
rect 3698 632088 3754 632097
rect 3698 632023 3754 632032
rect 3700 631372 3752 631378
rect 3700 631314 3752 631320
rect 3606 475688 3662 475697
rect 3606 475623 3662 475632
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3422 449576 3478 449585
rect 3422 449511 3478 449520
rect 3712 423609 3740 631314
rect 3804 501809 3832 678286
rect 3884 678224 3936 678230
rect 3884 678166 3936 678172
rect 3896 514865 3924 678166
rect 3988 527921 4016 684694
rect 6932 683777 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 19984 684820 20036 684826
rect 19984 684762 20036 684768
rect 6918 683768 6974 683777
rect 6918 683703 6974 683712
rect 4068 683324 4120 683330
rect 4068 683266 4120 683272
rect 4080 553897 4108 683266
rect 17684 670744 17736 670750
rect 17684 670686 17736 670692
rect 17696 667418 17724 670686
rect 13820 667412 13872 667418
rect 13820 667354 13872 667360
rect 17684 667412 17736 667418
rect 17684 667354 17736 667360
rect 13832 665242 13860 667354
rect 13820 665236 13872 665242
rect 13820 665178 13872 665184
rect 11796 665168 11848 665174
rect 11796 665110 11848 665116
rect 11808 659734 11836 665110
rect 11796 659728 11848 659734
rect 11796 659670 11848 659676
rect 7564 659660 7616 659666
rect 7564 659602 7616 659608
rect 7576 655586 7604 659602
rect 19996 658238 20024 684762
rect 23492 683913 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 40512 700330 40540 703520
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 40500 700324 40552 700330
rect 40500 700266 40552 700272
rect 71792 685166 71820 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 88352 685234 88380 702406
rect 105464 700398 105492 703520
rect 105452 700392 105504 700398
rect 137848 700369 137876 703520
rect 154132 700466 154160 703520
rect 170324 700505 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 170310 700496 170366 700505
rect 154120 700460 154172 700466
rect 170310 700431 170366 700440
rect 154120 700402 154172 700408
rect 105452 700334 105504 700340
rect 137834 700360 137890 700369
rect 137834 700295 137890 700304
rect 88340 685228 88392 685234
rect 88340 685170 88392 685176
rect 71780 685160 71832 685166
rect 71780 685102 71832 685108
rect 201512 684049 201540 702986
rect 218072 685302 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 235184 700641 235212 703520
rect 235170 700632 235226 700641
rect 235170 700567 235226 700576
rect 267660 697610 267688 703520
rect 283852 700534 283880 703520
rect 300136 700602 300164 703520
rect 332520 700670 332548 703520
rect 348804 702434 348832 703520
rect 347792 702406 348832 702434
rect 332508 700664 332560 700670
rect 332508 700606 332560 700612
rect 300124 700596 300176 700602
rect 300124 700538 300176 700544
rect 283840 700528 283892 700534
rect 283840 700470 283892 700476
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 218060 685296 218112 685302
rect 218060 685238 218112 685244
rect 201498 684040 201554 684049
rect 201498 683975 201554 683984
rect 23478 683904 23534 683913
rect 23478 683839 23534 683848
rect 266372 683806 266400 697546
rect 347792 685370 347820 702406
rect 364996 700738 365024 703520
rect 364984 700732 365036 700738
rect 364984 700674 365036 700680
rect 347780 685364 347832 685370
rect 347780 685306 347832 685312
rect 266360 683800 266412 683806
rect 266360 683742 266412 683748
rect 20812 683596 20864 683602
rect 20812 683538 20864 683544
rect 359464 683596 359516 683602
rect 359464 683538 359516 683544
rect 20824 681766 20852 683538
rect 21364 683528 21416 683534
rect 21364 683470 21416 683476
rect 20076 681760 20128 681766
rect 20076 681702 20128 681708
rect 20812 681760 20864 681766
rect 20812 681702 20864 681708
rect 20088 670750 20116 681702
rect 20076 670744 20128 670750
rect 20076 670686 20128 670692
rect 19984 658232 20036 658238
rect 19984 658174 20036 658180
rect 6184 655580 6236 655586
rect 6184 655522 6236 655528
rect 7564 655580 7616 655586
rect 7564 655522 7616 655528
rect 6196 652798 6224 655522
rect 4804 652792 4856 652798
rect 4804 652734 4856 652740
rect 6184 652792 6236 652798
rect 6184 652734 6236 652740
rect 4066 553888 4122 553897
rect 4066 553823 4122 553832
rect 3974 527912 4030 527921
rect 3974 527847 4030 527856
rect 3882 514856 3938 514865
rect 4816 514826 4844 652734
rect 21376 634814 21404 683470
rect 20916 634786 21404 634814
rect 20916 631378 20944 634786
rect 20904 631372 20956 631378
rect 20904 631314 20956 631320
rect 359476 616826 359504 683538
rect 361764 679040 361816 679046
rect 361762 679008 361764 679017
rect 365076 679040 365128 679046
rect 361816 679008 361818 679017
rect 365076 678982 365128 678988
rect 361762 678943 361818 678952
rect 361762 667992 361818 668001
rect 361762 667927 361764 667936
rect 361816 667927 361818 667936
rect 361764 667898 361816 667904
rect 361762 656976 361818 656985
rect 361762 656911 361764 656920
rect 361816 656911 361818 656920
rect 361764 656882 361816 656888
rect 361762 645960 361818 645969
rect 361762 645895 361764 645904
rect 361816 645895 361818 645904
rect 361764 645866 361816 645872
rect 361578 634944 361634 634953
rect 361578 634879 361634 634888
rect 361592 634846 361620 634879
rect 361580 634840 361632 634846
rect 361580 634782 361632 634788
rect 361578 623928 361634 623937
rect 361578 623863 361634 623872
rect 361592 623830 361620 623863
rect 361580 623824 361632 623830
rect 361580 623766 361632 623772
rect 359464 616820 359516 616826
rect 359464 616762 359516 616768
rect 360936 616820 360988 616826
rect 360936 616762 360988 616768
rect 360948 611250 360976 616762
rect 361578 612912 361634 612921
rect 361578 612847 361634 612856
rect 361592 612814 361620 612847
rect 361580 612808 361632 612814
rect 361580 612750 361632 612756
rect 360936 611244 360988 611250
rect 360936 611186 360988 611192
rect 362224 611244 362276 611250
rect 362224 611186 362276 611192
rect 361762 601896 361818 601905
rect 361762 601831 361818 601840
rect 361776 601730 361804 601831
rect 361764 601724 361816 601730
rect 361764 601666 361816 601672
rect 362236 600302 362264 611186
rect 362224 600296 362276 600302
rect 362224 600238 362276 600244
rect 362960 600296 363012 600302
rect 362960 600238 363012 600244
rect 362972 596834 363000 600238
rect 362960 596828 363012 596834
rect 362960 596770 363012 596776
rect 361762 590880 361818 590889
rect 361762 590815 361818 590824
rect 361776 590714 361804 590815
rect 361764 590708 361816 590714
rect 361764 590650 361816 590656
rect 361762 579864 361818 579873
rect 361762 579799 361818 579808
rect 361776 579698 361804 579799
rect 361764 579692 361816 579698
rect 361764 579634 361816 579640
rect 361762 568848 361818 568857
rect 361762 568783 361818 568792
rect 361776 568614 361804 568783
rect 361764 568608 361816 568614
rect 361764 568550 361816 568556
rect 361578 557832 361634 557841
rect 361578 557767 361580 557776
rect 361632 557767 361634 557776
rect 363604 557796 363656 557802
rect 361580 557738 361632 557744
rect 363604 557738 363656 557744
rect 361578 546816 361634 546825
rect 361578 546751 361634 546760
rect 361592 546650 361620 546751
rect 361580 546644 361632 546650
rect 361580 546586 361632 546592
rect 361578 535800 361634 535809
rect 361578 535735 361580 535744
rect 361632 535735 361634 535744
rect 361580 535706 361632 535712
rect 361762 524784 361818 524793
rect 361762 524719 361818 524728
rect 361776 524482 361804 524719
rect 361764 524476 361816 524482
rect 361764 524418 361816 524424
rect 3882 514791 3938 514800
rect 3976 514820 4028 514826
rect 3976 514762 4028 514768
rect 4804 514820 4856 514826
rect 4804 514762 4856 514768
rect 3790 501800 3846 501809
rect 3790 501735 3846 501744
rect 3698 423600 3754 423609
rect 3698 423535 3754 423544
rect 3988 410553 4016 514762
rect 361762 513768 361818 513777
rect 361762 513703 361818 513712
rect 361776 513398 361804 513703
rect 361764 513392 361816 513398
rect 361764 513334 361816 513340
rect 361762 502752 361818 502761
rect 361762 502687 361818 502696
rect 361776 502382 361804 502687
rect 361764 502376 361816 502382
rect 361764 502318 361816 502324
rect 362222 491736 362278 491745
rect 362222 491671 362278 491680
rect 361762 480720 361818 480729
rect 361762 480655 361818 480664
rect 361776 480282 361804 480655
rect 361764 480276 361816 480282
rect 361764 480218 361816 480224
rect 361762 469704 361818 469713
rect 361762 469639 361818 469648
rect 361776 469266 361804 469639
rect 361764 469260 361816 469266
rect 361764 469202 361816 469208
rect 361762 458688 361818 458697
rect 361762 458623 361818 458632
rect 361776 458250 361804 458623
rect 361764 458244 361816 458250
rect 361764 458186 361816 458192
rect 361762 436656 361818 436665
rect 361762 436591 361818 436600
rect 361776 436150 361804 436591
rect 361764 436144 361816 436150
rect 361764 436086 361816 436092
rect 361578 414624 361634 414633
rect 361578 414559 361634 414568
rect 361592 414050 361620 414559
rect 361580 414044 361632 414050
rect 361580 413986 361632 413992
rect 3974 410544 4030 410553
rect 3974 410479 4030 410488
rect 361578 403608 361634 403617
rect 361578 403543 361634 403552
rect 361592 403034 361620 403543
rect 361580 403028 361632 403034
rect 361580 402970 361632 402976
rect 3882 397488 3938 397497
rect 3882 397423 3938 397432
rect 3422 358456 3478 358465
rect 3422 358391 3478 358400
rect 3436 305046 3464 358391
rect 3514 345400 3570 345409
rect 3514 345335 3570 345344
rect 3424 305040 3476 305046
rect 3424 304982 3476 304988
rect 3422 293176 3478 293185
rect 3422 293111 3478 293120
rect 3330 162888 3386 162897
rect 3330 162823 3386 162832
rect 3238 149832 3294 149841
rect 3238 149767 3294 149776
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3160 84250 3188 84623
rect 3148 84244 3200 84250
rect 3148 84186 3200 84192
rect 3146 71632 3202 71641
rect 3146 71567 3202 71576
rect 3160 70446 3188 71567
rect 3148 70440 3200 70446
rect 3148 70382 3200 70388
rect 3252 46782 3280 149767
rect 3240 46776 3292 46782
rect 3240 46718 3292 46724
rect 3344 46714 3372 162823
rect 3436 59945 3464 293111
rect 3528 292806 3556 345335
rect 3790 319288 3846 319297
rect 3790 319223 3846 319232
rect 3698 306232 3754 306241
rect 3698 306167 3754 306176
rect 3516 292800 3568 292806
rect 3516 292742 3568 292748
rect 3514 267200 3570 267209
rect 3514 267135 3570 267144
rect 3422 59936 3478 59945
rect 3422 59871 3478 59880
rect 3422 58576 3478 58585
rect 3422 58511 3478 58520
rect 3332 46708 3384 46714
rect 3332 46650 3384 46656
rect 2780 39364 2832 39370
rect 2780 39306 2832 39312
rect 2792 16574 2820 39306
rect 3436 31754 3464 58511
rect 3528 46918 3556 267135
rect 3606 254144 3662 254153
rect 3606 254079 3662 254088
rect 3516 46912 3568 46918
rect 3516 46854 3568 46860
rect 3620 46510 3648 254079
rect 3712 98666 3740 306167
rect 3804 253978 3832 319223
rect 3792 253972 3844 253978
rect 3792 253914 3844 253920
rect 3896 241466 3924 397423
rect 361578 392592 361634 392601
rect 361578 392527 361634 392536
rect 361592 392018 361620 392527
rect 361580 392012 361632 392018
rect 361580 391954 361632 391960
rect 360844 386436 360896 386442
rect 360844 386378 360896 386384
rect 3974 371376 4030 371385
rect 3974 371311 4030 371320
rect 3884 241460 3936 241466
rect 3884 241402 3936 241408
rect 3790 241088 3846 241097
rect 3790 241023 3846 241032
rect 3700 98660 3752 98666
rect 3700 98602 3752 98608
rect 3698 97608 3754 97617
rect 3698 97543 3754 97552
rect 3712 46850 3740 97543
rect 3700 46844 3752 46850
rect 3700 46786 3752 46792
rect 3608 46504 3660 46510
rect 3608 46446 3660 46452
rect 3804 46442 3832 241023
rect 3882 214976 3938 214985
rect 3882 214911 3938 214920
rect 3896 46578 3924 214911
rect 3988 214810 4016 371311
rect 359464 305652 359516 305658
rect 359464 305594 359516 305600
rect 4804 305040 4856 305046
rect 4804 304982 4856 304988
rect 3976 214804 4028 214810
rect 3976 214746 4028 214752
rect 3974 201920 4030 201929
rect 3974 201855 4030 201864
rect 3988 46646 4016 201855
rect 4066 188864 4122 188873
rect 4066 188799 4122 188808
rect 3976 46640 4028 46646
rect 3976 46582 4028 46588
rect 3884 46572 3936 46578
rect 3884 46514 3936 46520
rect 3792 46436 3844 46442
rect 3792 46378 3844 46384
rect 4080 45626 4108 188799
rect 4816 66910 4844 304982
rect 4896 292800 4948 292806
rect 4896 292742 4948 292748
rect 4908 98054 4936 292742
rect 4988 253972 5040 253978
rect 4988 253914 5040 253920
rect 4896 98048 4948 98054
rect 4896 97990 4948 97996
rect 5000 71262 5028 253914
rect 5080 241460 5132 241466
rect 5080 241402 5132 241408
rect 4988 71256 5040 71262
rect 4988 71198 5040 71204
rect 4804 66904 4856 66910
rect 4804 66846 4856 66852
rect 5092 60722 5120 241402
rect 5172 214804 5224 214810
rect 5172 214746 5224 214752
rect 5080 60716 5132 60722
rect 5080 60658 5132 60664
rect 5184 57254 5212 214746
rect 19984 98660 20036 98666
rect 19984 98602 20036 98608
rect 8944 97980 8996 97986
rect 8944 97922 8996 97928
rect 6184 71256 6236 71262
rect 6184 71198 6236 71204
rect 6000 60716 6052 60722
rect 6000 60658 6052 60664
rect 6012 58682 6040 60658
rect 6000 58676 6052 58682
rect 6000 58618 6052 58624
rect 5172 57248 5224 57254
rect 5172 57190 5224 57196
rect 6196 53854 6224 71198
rect 8956 67590 8984 97922
rect 8944 67584 8996 67590
rect 8944 67526 8996 67532
rect 10968 67584 11020 67590
rect 10968 67526 11020 67532
rect 7288 66904 7340 66910
rect 7288 66846 7340 66852
rect 7300 63714 7328 66846
rect 10980 64874 11008 67526
rect 10980 64846 11100 64874
rect 7288 63708 7340 63714
rect 7288 63650 7340 63656
rect 9680 63708 9732 63714
rect 9680 63650 9732 63656
rect 8208 57248 8260 57254
rect 8208 57190 8260 57196
rect 6184 53848 6236 53854
rect 6184 53790 6236 53796
rect 8220 52494 8248 57190
rect 9692 55282 9720 63650
rect 11072 59430 11100 64846
rect 11060 59424 11112 59430
rect 11060 59366 11112 59372
rect 13820 59356 13872 59362
rect 13820 59298 13872 59304
rect 11704 58676 11756 58682
rect 11704 58618 11756 58624
rect 9680 55276 9732 55282
rect 9680 55218 9732 55224
rect 8392 53780 8444 53786
rect 8392 53722 8444 53728
rect 8208 52488 8260 52494
rect 8208 52430 8260 52436
rect 8404 51746 8432 53722
rect 11716 53446 11744 58618
rect 13832 56574 13860 59298
rect 13820 56568 13872 56574
rect 13820 56510 13872 56516
rect 16488 56568 16540 56574
rect 16488 56510 16540 56516
rect 13728 55208 13780 55214
rect 13728 55150 13780 55156
rect 13740 53802 13768 55150
rect 16500 53802 16528 56510
rect 13740 53774 13860 53802
rect 16500 53774 16620 53802
rect 11704 53440 11756 53446
rect 11704 53382 11756 53388
rect 13728 53440 13780 53446
rect 13728 53382 13780 53388
rect 11060 52420 11112 52426
rect 11060 52362 11112 52368
rect 8392 51740 8444 51746
rect 8392 51682 8444 51688
rect 11072 49774 11100 52362
rect 13740 51134 13768 53382
rect 13728 51128 13780 51134
rect 13728 51070 13780 51076
rect 13832 50998 13860 53774
rect 13820 50992 13872 50998
rect 13820 50934 13872 50940
rect 16592 50182 16620 53774
rect 19248 51740 19300 51746
rect 19248 51682 19300 51688
rect 17868 51060 17920 51066
rect 17868 51002 17920 51008
rect 16580 50176 16632 50182
rect 16580 50118 16632 50124
rect 11060 49768 11112 49774
rect 11060 49710 11112 49716
rect 17880 48210 17908 51002
rect 18604 50992 18656 50998
rect 18604 50934 18656 50940
rect 18236 49700 18288 49706
rect 18236 49642 18288 49648
rect 17868 48204 17920 48210
rect 17868 48146 17920 48152
rect 18248 47938 18276 49642
rect 18616 48346 18644 50934
rect 19260 49450 19288 51682
rect 19340 50176 19392 50182
rect 19340 50118 19392 50124
rect 19352 49609 19380 50118
rect 19338 49600 19394 49609
rect 19338 49535 19394 49544
rect 19260 49422 19380 49450
rect 18604 48340 18656 48346
rect 18604 48282 18656 48288
rect 18236 47932 18288 47938
rect 18236 47874 18288 47880
rect 19352 47054 19380 49422
rect 19340 47048 19392 47054
rect 19340 46990 19392 46996
rect 19996 46306 20024 98602
rect 20904 84244 20956 84250
rect 20956 84192 21404 84194
rect 20904 84186 21404 84192
rect 20916 84166 21404 84186
rect 20076 70440 20128 70446
rect 20076 70382 20128 70388
rect 20088 46374 20116 70382
rect 20904 48272 20956 48278
rect 20904 48214 20956 48220
rect 20720 48204 20772 48210
rect 20720 48146 20772 48152
rect 20076 46368 20128 46374
rect 20076 46310 20128 46316
rect 19984 46300 20036 46306
rect 19984 46242 20036 46248
rect 20732 46170 20760 48146
rect 20812 47932 20864 47938
rect 20812 47874 20864 47880
rect 20824 46238 20852 47874
rect 20812 46232 20864 46238
rect 20812 46174 20864 46180
rect 20720 46164 20772 46170
rect 20720 46106 20772 46112
rect 4068 45620 4120 45626
rect 4068 45562 4120 45568
rect 3514 45520 3570 45529
rect 3514 45455 3516 45464
rect 3568 45455 3570 45464
rect 3516 45426 3568 45432
rect 20916 45422 20944 48214
rect 21272 47048 21324 47054
rect 21272 46990 21324 46996
rect 21284 46102 21312 46990
rect 21376 46753 21404 84166
rect 21362 46744 21418 46753
rect 21362 46679 21418 46688
rect 21272 46096 21324 46102
rect 21272 46038 21324 46044
rect 358176 45824 358228 45830
rect 358176 45766 358228 45772
rect 358188 45422 358216 45766
rect 20904 45416 20956 45422
rect 20904 45358 20956 45364
rect 358176 45416 358228 45422
rect 358176 45358 358228 45364
rect 71780 45348 71832 45354
rect 71780 45290 71832 45296
rect 69020 45280 69072 45286
rect 69020 45222 69072 45228
rect 64880 45212 64932 45218
rect 64880 45154 64932 45160
rect 60740 45144 60792 45150
rect 60740 45086 60792 45092
rect 57980 45076 58032 45082
rect 57980 45018 58032 45024
rect 53840 45008 53892 45014
rect 53840 44950 53892 44956
rect 51080 44940 51132 44946
rect 51080 44882 51132 44888
rect 6920 44872 6972 44878
rect 6920 44814 6972 44820
rect 46938 44840 46994 44849
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3424 31748 3476 31754
rect 3424 31690 3476 31696
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 6932 16574 6960 44814
rect 46938 44775 46994 44784
rect 20720 42152 20772 42158
rect 20720 42094 20772 42100
rect 11060 42084 11112 42090
rect 11060 42026 11112 42032
rect 9680 33788 9732 33794
rect 9680 33730 9732 33736
rect 2792 16546 3648 16574
rect 6932 16546 7696 16574
rect 572 7608 624 7614
rect 572 7550 624 7556
rect 584 480 612 7550
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 1674 3360 1730 3369
rect 1674 3295 1730 3304
rect 1688 480 1716 3295
rect 2872 2100 2924 2106
rect 2872 2042 2924 2048
rect 2884 480 2912 2042
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3620 354 3648 16546
rect 5262 3904 5318 3913
rect 5262 3839 5318 3848
rect 5276 480 5304 3839
rect 6460 3256 6512 3262
rect 6460 3198 6512 3204
rect 6472 480 6500 3198
rect 7668 480 7696 16546
rect 8758 3768 8814 3777
rect 8758 3703 8814 3712
rect 8772 480 8800 3703
rect 4038 354 4150 480
rect 3620 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 33730
rect 11072 16574 11100 42026
rect 17960 36576 18012 36582
rect 17960 36518 18012 36524
rect 13820 31068 13872 31074
rect 13820 31010 13872 31016
rect 13832 16574 13860 31010
rect 11072 16546 11928 16574
rect 13832 16546 14320 16574
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 11900 354 11928 16546
rect 13542 3632 13598 3641
rect 13542 3567 13598 3576
rect 13556 480 13584 3567
rect 12318 354 12430 480
rect 11900 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 17038 4040 17094 4049
rect 17038 3975 17094 3984
rect 17052 480 17080 3975
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 36518
rect 19340 31204 19392 31210
rect 19340 31146 19392 31152
rect 19352 16574 19380 31146
rect 20732 16574 20760 42094
rect 44180 39636 44232 39642
rect 44180 39578 44232 39584
rect 40040 39568 40092 39574
rect 40040 39510 40092 39516
rect 33140 39500 33192 39506
rect 33140 39442 33192 39448
rect 26240 39432 26292 39438
rect 26240 39374 26292 39380
rect 22100 36644 22152 36650
rect 22100 36586 22152 36592
rect 22112 16574 22140 36586
rect 19352 16546 19472 16574
rect 20732 16546 21864 16574
rect 22112 16546 22600 16574
rect 19444 480 19472 16546
rect 21836 480 21864 16546
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 24214 3496 24270 3505
rect 24214 3431 24270 3440
rect 24228 480 24256 3431
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 39374
rect 30380 33856 30432 33862
rect 30380 33798 30432 33804
rect 30392 16574 30420 33798
rect 31760 31136 31812 31142
rect 31760 31078 31812 31084
rect 31772 16574 31800 31078
rect 33152 16574 33180 39442
rect 34520 33924 34572 33930
rect 34520 33866 34572 33872
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 33152 16546 33640 16574
rect 27712 3528 27764 3534
rect 27712 3470 27764 3476
rect 27724 480 27752 3470
rect 28908 3188 28960 3194
rect 28908 3130 28960 3136
rect 28920 480 28948 3130
rect 30104 2168 30156 2174
rect 30104 2110 30156 2116
rect 30116 480 30144 2110
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 33612 480 33640 16546
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 33866
rect 35900 31272 35952 31278
rect 35900 31214 35952 31220
rect 35912 16574 35940 31214
rect 38660 28280 38712 28286
rect 38660 28222 38712 28228
rect 38672 16574 38700 28222
rect 40052 16574 40080 39510
rect 35912 16546 36032 16574
rect 38672 16546 39160 16574
rect 40052 16546 40264 16574
rect 36004 480 36032 16546
rect 37188 3664 37240 3670
rect 37188 3606 37240 3612
rect 37200 480 37228 3606
rect 38384 3460 38436 3466
rect 38384 3402 38436 3408
rect 38396 480 38424 3402
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 44192 6914 44220 39578
rect 44272 33992 44324 33998
rect 44272 33934 44324 33940
rect 44284 16574 44312 33934
rect 45560 28348 45612 28354
rect 45560 28290 45612 28296
rect 45572 16574 45600 28290
rect 46952 16574 46980 44775
rect 49700 34060 49752 34066
rect 49700 34002 49752 34008
rect 49712 16574 49740 34002
rect 44284 16546 45048 16574
rect 45572 16546 46704 16574
rect 46952 16546 47440 16574
rect 49712 16546 50200 16574
rect 44192 6886 44312 6914
rect 43076 3800 43128 3806
rect 43076 3742 43128 3748
rect 41880 3596 41932 3602
rect 41880 3538 41932 3544
rect 41892 480 41920 3538
rect 43088 480 43116 3742
rect 44284 480 44312 6886
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45020 354 45048 16546
rect 46676 480 46704 16546
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 48964 3868 49016 3874
rect 48964 3810 49016 3816
rect 48976 480 49004 3810
rect 50172 480 50200 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 47830 -960 47942 326
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51092 354 51120 44882
rect 52460 34128 52512 34134
rect 52460 34070 52512 34076
rect 52472 16574 52500 34070
rect 53852 16574 53880 44950
rect 57992 16574 58020 45018
rect 59360 39704 59412 39710
rect 59360 39646 59412 39652
rect 52472 16546 53328 16574
rect 53852 16546 54984 16574
rect 57992 16546 58480 16574
rect 52552 3732 52604 3738
rect 52552 3674 52604 3680
rect 52564 480 52592 3674
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53300 354 53328 16546
rect 54956 480 54984 16546
rect 56048 4004 56100 4010
rect 56048 3946 56100 3952
rect 56060 480 56088 3946
rect 57244 3936 57296 3942
rect 57244 3878 57296 3884
rect 57256 480 57284 3878
rect 58452 480 58480 16546
rect 53718 354 53830 480
rect 53300 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59372 354 59400 39646
rect 60752 3398 60780 45086
rect 62120 39772 62172 39778
rect 62120 39714 62172 39720
rect 60832 34196 60884 34202
rect 60832 34138 60884 34144
rect 60740 3392 60792 3398
rect 60740 3334 60792 3340
rect 60844 480 60872 34138
rect 62132 16574 62160 39714
rect 63500 34264 63552 34270
rect 63500 34206 63552 34212
rect 63512 16574 63540 34206
rect 64892 16574 64920 45154
rect 66260 39840 66312 39846
rect 66260 39782 66312 39788
rect 66272 16574 66300 39782
rect 67640 34400 67692 34406
rect 67640 34342 67692 34348
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 64892 16546 65104 16574
rect 66272 16546 66760 16574
rect 61660 3392 61712 3398
rect 61660 3334 61712 3340
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61672 354 61700 3334
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 61998 354 62110 480
rect 61672 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66732 480 66760 16546
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 34342
rect 69032 6914 69060 45222
rect 69112 39908 69164 39914
rect 69112 39850 69164 39856
rect 69124 16574 69152 39850
rect 70400 34332 70452 34338
rect 70400 34274 70452 34280
rect 70412 16574 70440 34274
rect 71792 16574 71820 45290
rect 75920 44804 75972 44810
rect 75920 44746 75972 44752
rect 73160 39976 73212 39982
rect 73160 39918 73212 39924
rect 73172 16574 73200 39918
rect 74540 34468 74592 34474
rect 74540 34410 74592 34416
rect 74552 16574 74580 34410
rect 69124 16546 69888 16574
rect 70412 16546 71544 16574
rect 71792 16546 72648 16574
rect 73172 16546 73384 16574
rect 74552 16546 75040 16574
rect 69032 6886 69152 6914
rect 69124 480 69152 6886
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 16546
rect 71516 480 71544 16546
rect 72620 480 72648 16546
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 75012 480 75040 16546
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 44746
rect 78680 44736 78732 44742
rect 78680 44678 78732 44684
rect 77300 40044 77352 40050
rect 77300 39986 77352 39992
rect 77312 6914 77340 39986
rect 77392 33720 77444 33726
rect 77392 33662 77444 33668
rect 77404 16574 77432 33662
rect 78692 16574 78720 44678
rect 85580 44668 85632 44674
rect 85580 44610 85632 44616
rect 82820 42220 82872 42226
rect 82820 42162 82872 42168
rect 80060 39296 80112 39302
rect 80060 39238 80112 39244
rect 80072 16574 80100 39238
rect 82832 16574 82860 42162
rect 84200 39228 84252 39234
rect 84200 39170 84252 39176
rect 77404 16546 78168 16574
rect 78692 16546 79272 16574
rect 80072 16546 80928 16574
rect 82832 16546 83320 16574
rect 77312 6886 77432 6914
rect 77404 480 77432 6886
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78140 354 78168 16546
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 79244 354 79272 16546
rect 80900 480 80928 16546
rect 82084 4072 82136 4078
rect 82084 4014 82136 4020
rect 82096 480 82124 4014
rect 83292 480 83320 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84212 354 84240 39170
rect 85592 3398 85620 44610
rect 114560 42764 114612 42770
rect 114560 42706 114612 42712
rect 110420 42696 110472 42702
rect 110420 42638 110472 42644
rect 107660 42628 107712 42634
rect 107660 42570 107712 42576
rect 103520 42560 103572 42566
rect 103520 42502 103572 42508
rect 100760 42492 100812 42498
rect 100760 42434 100812 42440
rect 96620 42424 96672 42430
rect 96620 42366 96672 42372
rect 93860 42356 93912 42362
rect 93860 42298 93912 42304
rect 89720 42288 89772 42294
rect 89720 42230 89772 42236
rect 86960 36712 87012 36718
rect 86960 36654 87012 36660
rect 85672 33652 85724 33658
rect 85672 33594 85724 33600
rect 85580 3392 85632 3398
rect 85580 3334 85632 3340
rect 85684 480 85712 33594
rect 86972 16574 87000 36654
rect 89732 16574 89760 42230
rect 91100 36780 91152 36786
rect 91100 36722 91152 36728
rect 91112 16574 91140 36722
rect 92480 31340 92532 31346
rect 92480 31282 92532 31288
rect 86972 16546 87552 16574
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 86500 3392 86552 3398
rect 86500 3334 86552 3340
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86512 354 86540 3334
rect 86838 354 86950 480
rect 86512 326 86950 354
rect 87524 354 87552 16546
rect 89168 4140 89220 4146
rect 89168 4082 89220 4088
rect 89180 480 89208 4082
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 31282
rect 93872 6914 93900 42298
rect 93952 36848 94004 36854
rect 93952 36790 94004 36796
rect 93964 16574 93992 36790
rect 96632 16574 96660 42366
rect 98000 36916 98052 36922
rect 98000 36858 98052 36864
rect 98012 16574 98040 36858
rect 99380 31408 99432 31414
rect 99380 31350 99432 31356
rect 99392 16574 99420 31350
rect 93964 16546 94728 16574
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 93872 6886 93992 6914
rect 93964 480 93992 6886
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94700 354 94728 16546
rect 96252 3392 96304 3398
rect 96252 3334 96304 3340
rect 96264 480 96292 3334
rect 97460 480 97488 16546
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95118 -960 95230 326
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 42434
rect 102140 36984 102192 36990
rect 102140 36926 102192 36932
rect 102152 6914 102180 36926
rect 102232 31544 102284 31550
rect 102232 31486 102284 31492
rect 102244 16574 102272 31486
rect 103532 16574 103560 42502
rect 104900 37052 104952 37058
rect 104900 36994 104952 37000
rect 104912 16574 104940 36994
rect 106924 28416 106976 28422
rect 106924 28358 106976 28364
rect 102244 16546 103376 16574
rect 103532 16546 104112 16574
rect 104912 16546 105768 16574
rect 102152 6886 102272 6914
rect 102244 480 102272 6886
rect 103348 480 103376 16546
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105740 480 105768 16546
rect 106936 6914 106964 28358
rect 107672 16574 107700 42570
rect 109040 37120 109092 37126
rect 109040 37062 109092 37068
rect 107672 16546 108160 16574
rect 106844 6886 106964 6914
rect 106844 3262 106872 6886
rect 106832 3256 106884 3262
rect 106832 3198 106884 3204
rect 106924 3188 106976 3194
rect 106924 3130 106976 3136
rect 106936 480 106964 3130
rect 108132 480 108160 16546
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109052 354 109080 37062
rect 110432 3330 110460 42638
rect 111800 37188 111852 37194
rect 111800 37130 111852 37136
rect 111064 31476 111116 31482
rect 111064 31418 111116 31424
rect 110420 3324 110472 3330
rect 110420 3266 110472 3272
rect 111076 3126 111104 31418
rect 111812 16574 111840 37130
rect 113180 31612 113232 31618
rect 113180 31554 113232 31560
rect 113192 16574 113220 31554
rect 114572 16574 114600 42706
rect 118700 42016 118752 42022
rect 118700 41958 118752 41964
rect 115940 37256 115992 37262
rect 115940 37198 115992 37204
rect 115952 16574 115980 37198
rect 117320 31000 117372 31006
rect 117320 30942 117372 30948
rect 111812 16546 112392 16574
rect 113192 16546 114048 16574
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 111616 3324 111668 3330
rect 111616 3266 111668 3272
rect 111064 3120 111116 3126
rect 111064 3062 111116 3068
rect 110512 3052 110564 3058
rect 110512 2994 110564 3000
rect 110524 480 110552 2994
rect 111628 480 111656 3266
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114020 480 114048 16546
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 30942
rect 118712 6914 118740 41958
rect 121460 41948 121512 41954
rect 121460 41890 121512 41896
rect 118792 36508 118844 36514
rect 118792 36450 118844 36456
rect 118804 16574 118832 36450
rect 120080 31680 120132 31686
rect 120080 31622 120132 31628
rect 120092 16574 120120 31622
rect 121472 16574 121500 41890
rect 122840 36440 122892 36446
rect 122840 36382 122892 36388
rect 122852 16574 122880 36382
rect 124220 30932 124272 30938
rect 124220 30874 124272 30880
rect 124232 16574 124260 30874
rect 118804 16546 119936 16574
rect 120092 16546 120672 16574
rect 121472 16546 122328 16574
rect 122852 16546 123064 16574
rect 124232 16546 124720 16574
rect 118712 6886 118832 6914
rect 118804 480 118832 6886
rect 119908 480 119936 16546
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 122300 480 122328 16546
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124692 480 124720 16546
rect 359476 4010 359504 305594
rect 359556 304292 359608 304298
rect 359556 304234 359608 304240
rect 359464 4004 359516 4010
rect 359464 3946 359516 3952
rect 359568 3398 359596 304234
rect 359648 276684 359700 276690
rect 359648 276626 359700 276632
rect 359660 4078 359688 276626
rect 359832 160744 359884 160750
rect 359832 160686 359884 160692
rect 359740 160132 359792 160138
rect 359740 160074 359792 160080
rect 359752 46102 359780 160074
rect 359844 46170 359872 160686
rect 359924 155916 359976 155922
rect 359924 155858 359976 155864
rect 359936 46238 359964 155858
rect 359924 46232 359976 46238
rect 359924 46174 359976 46180
rect 359832 46164 359884 46170
rect 359832 46106 359884 46112
rect 359740 46096 359792 46102
rect 359740 46038 359792 46044
rect 360856 31006 360884 386378
rect 361578 381576 361634 381585
rect 361578 381511 361634 381520
rect 361592 380934 361620 381511
rect 361580 380928 361632 380934
rect 361580 380870 361632 380876
rect 362236 372570 362264 491671
rect 362314 447672 362370 447681
rect 362314 447607 362370 447616
rect 362328 416090 362356 447607
rect 362406 425640 362462 425649
rect 362406 425575 362462 425584
rect 362420 418810 362448 425575
rect 362408 418804 362460 418810
rect 362408 418746 362460 418752
rect 362316 416084 362368 416090
rect 362316 416026 362368 416032
rect 363616 376650 363644 557738
rect 363696 546644 363748 546650
rect 363696 546586 363748 546592
rect 363708 376718 363736 546586
rect 363788 535764 363840 535770
rect 363788 535706 363840 535712
rect 363696 376712 363748 376718
rect 363696 376654 363748 376660
rect 363604 376644 363656 376650
rect 363604 376586 363656 376592
rect 363800 375358 363828 535706
rect 364984 386504 365036 386510
rect 364984 386446 365036 386452
rect 363788 375352 363840 375358
rect 363788 375294 363840 375300
rect 362224 372564 362276 372570
rect 362224 372506 362276 372512
rect 361578 370560 361634 370569
rect 361578 370495 361634 370504
rect 361592 369918 361620 370495
rect 361580 369912 361632 369918
rect 361580 369854 361632 369860
rect 362314 359544 362370 359553
rect 362314 359479 362370 359488
rect 361762 348528 361818 348537
rect 361762 348463 361818 348472
rect 361776 347818 361804 348463
rect 361764 347812 361816 347818
rect 361764 347754 361816 347760
rect 362328 347750 362356 359479
rect 362316 347744 362368 347750
rect 362316 347686 362368 347692
rect 361764 340944 361816 340950
rect 361764 340886 361816 340892
rect 361776 337521 361804 340886
rect 361762 337512 361818 337521
rect 361762 337447 361818 337456
rect 362224 336048 362276 336054
rect 362224 335990 362276 335996
rect 362236 326505 362264 335990
rect 364064 334008 364116 334014
rect 364064 333950 364116 333956
rect 362222 326496 362278 326505
rect 362222 326431 362278 326440
rect 361764 315988 361816 315994
rect 361764 315930 361816 315936
rect 361776 315489 361804 315930
rect 361762 315480 361818 315489
rect 361762 315415 361818 315424
rect 360936 305720 360988 305726
rect 360936 305662 360988 305668
rect 360844 31000 360896 31006
rect 360844 30942 360896 30948
rect 359648 4072 359700 4078
rect 359648 4014 359700 4020
rect 359556 3392 359608 3398
rect 359556 3334 359608 3340
rect 360948 3262 360976 305662
rect 361764 304972 361816 304978
rect 361764 304914 361816 304920
rect 361776 304473 361804 304914
rect 361762 304464 361818 304473
rect 361762 304399 361818 304408
rect 361028 304360 361080 304366
rect 361028 304302 361080 304308
rect 361040 3913 361068 304302
rect 361118 302832 361174 302841
rect 361118 302767 361174 302776
rect 361026 3904 361082 3913
rect 361026 3839 361082 3848
rect 361132 3806 361160 302767
rect 363604 297968 363656 297974
rect 363604 297910 363656 297916
rect 361212 297764 361264 297770
rect 361212 297706 361264 297712
rect 361120 3800 361172 3806
rect 361120 3742 361172 3748
rect 361224 3330 361252 297706
rect 362316 297560 362368 297566
rect 362316 297502 362368 297508
rect 362224 297424 362276 297430
rect 362224 297366 362276 297372
rect 361304 295044 361356 295050
rect 361304 294986 361356 294992
rect 361316 40050 361344 294986
rect 361764 293956 361816 293962
rect 361764 293898 361816 293904
rect 361776 293457 361804 293898
rect 361762 293448 361818 293457
rect 361762 293383 361818 293392
rect 361764 282872 361816 282878
rect 361764 282814 361816 282820
rect 361776 282441 361804 282814
rect 361762 282432 361818 282441
rect 361762 282367 361818 282376
rect 361764 271856 361816 271862
rect 361764 271798 361816 271804
rect 361776 271425 361804 271798
rect 361762 271416 361818 271425
rect 361762 271351 361818 271360
rect 361764 260840 361816 260846
rect 361764 260782 361816 260788
rect 361776 260409 361804 260782
rect 361762 260400 361818 260409
rect 361762 260335 361818 260344
rect 361764 249756 361816 249762
rect 361764 249698 361816 249704
rect 361776 249393 361804 249698
rect 361762 249384 361818 249393
rect 361762 249319 361818 249328
rect 361764 238740 361816 238746
rect 361764 238682 361816 238688
rect 361776 238377 361804 238682
rect 361762 238368 361818 238377
rect 361762 238303 361818 238312
rect 361764 227724 361816 227730
rect 361764 227666 361816 227672
rect 361776 227361 361804 227666
rect 361762 227352 361818 227361
rect 361762 227287 361818 227296
rect 361672 216368 361724 216374
rect 361670 216336 361672 216345
rect 361724 216336 361726 216345
rect 361670 216271 361726 216280
rect 361764 205624 361816 205630
rect 361764 205566 361816 205572
rect 361776 205329 361804 205566
rect 361762 205320 361818 205329
rect 361762 205255 361818 205264
rect 361764 194540 361816 194546
rect 361764 194482 361816 194488
rect 361776 194313 361804 194482
rect 361762 194304 361818 194313
rect 361762 194239 361818 194248
rect 361764 183524 361816 183530
rect 361764 183466 361816 183472
rect 361776 183297 361804 183466
rect 361762 183288 361818 183297
rect 361762 183223 361818 183232
rect 361580 180124 361632 180130
rect 361580 180066 361632 180072
rect 361592 173890 361620 180066
rect 361408 173862 361620 173890
rect 361408 46481 361436 173862
rect 361762 172272 361818 172281
rect 361762 172207 361818 172216
rect 361776 171834 361804 172207
rect 361764 171828 361816 171834
rect 361764 171770 361816 171776
rect 361764 161424 361816 161430
rect 361764 161366 361816 161372
rect 361776 161265 361804 161366
rect 361762 161256 361818 161265
rect 361762 161191 361818 161200
rect 361764 139392 361816 139398
rect 361764 139334 361816 139340
rect 361776 139233 361804 139334
rect 361762 139224 361818 139233
rect 361762 139159 361818 139168
rect 361764 128308 361816 128314
rect 361764 128250 361816 128256
rect 361776 128217 361804 128250
rect 361762 128208 361818 128217
rect 361762 128143 361818 128152
rect 361764 117292 361816 117298
rect 361764 117234 361816 117240
rect 361776 117201 361804 117234
rect 361762 117192 361818 117201
rect 361762 117127 361818 117136
rect 361764 106276 361816 106282
rect 361764 106218 361816 106224
rect 361776 106185 361804 106218
rect 361762 106176 361818 106185
rect 361762 106111 361818 106120
rect 361764 84176 361816 84182
rect 361762 84144 361764 84153
rect 361816 84144 361818 84153
rect 361762 84079 361818 84088
rect 361764 73160 361816 73166
rect 361762 73128 361764 73137
rect 361816 73128 361818 73137
rect 361762 73063 361818 73072
rect 361762 62112 361818 62121
rect 361762 62047 361764 62056
rect 361816 62047 361818 62056
rect 361764 62018 361816 62024
rect 361764 51128 361816 51134
rect 361762 51096 361764 51105
rect 361816 51096 361818 51105
rect 361762 51031 361818 51040
rect 361394 46472 361450 46481
rect 361394 46407 361450 46416
rect 361304 40044 361356 40050
rect 361304 39986 361356 39992
rect 362236 39846 362264 297366
rect 362224 39840 362276 39846
rect 362224 39782 362276 39788
rect 362328 39778 362356 297502
rect 362408 294704 362460 294710
rect 362408 294646 362460 294652
rect 362420 39914 362448 294646
rect 362500 294636 362552 294642
rect 362500 294578 362552 294584
rect 362512 39982 362540 294578
rect 362684 167680 362736 167686
rect 362684 167622 362736 167628
rect 362592 161492 362644 161498
rect 362592 161434 362644 161440
rect 362604 150249 362632 161434
rect 362696 160138 362724 167622
rect 362684 160132 362736 160138
rect 362684 160074 362736 160080
rect 362590 150240 362646 150249
rect 362590 150175 362646 150184
rect 362592 124908 362644 124914
rect 362592 124850 362644 124856
rect 362604 45830 362632 124850
rect 362684 105596 362736 105602
rect 362684 105538 362736 105544
rect 362696 95169 362724 105538
rect 362682 95160 362738 95169
rect 362682 95095 362738 95104
rect 362592 45824 362644 45830
rect 362592 45766 362644 45772
rect 362500 39976 362552 39982
rect 362500 39918 362552 39924
rect 362408 39908 362460 39914
rect 362408 39850 362460 39856
rect 362316 39772 362368 39778
rect 362316 39714 362368 39720
rect 363616 4146 363644 297910
rect 363972 294840 364024 294846
rect 363972 294782 364024 294788
rect 363880 294772 363932 294778
rect 363880 294714 363932 294720
rect 363788 289264 363840 289270
rect 363788 289206 363840 289212
rect 363696 284980 363748 284986
rect 363696 284922 363748 284928
rect 363708 20670 363736 284922
rect 363800 31210 363828 289206
rect 363892 39302 363920 294714
rect 363880 39296 363932 39302
rect 363880 39238 363932 39244
rect 363984 39234 364012 294782
rect 364076 216374 364104 333950
rect 364064 216368 364116 216374
rect 364064 216310 364116 216316
rect 363972 39228 364024 39234
rect 363972 39170 364024 39176
rect 364996 31686 365024 386446
rect 365088 385014 365116 678982
rect 381544 667956 381596 667962
rect 381544 667898 381596 667904
rect 378784 645924 378836 645930
rect 378784 645866 378836 645872
rect 376024 623824 376076 623830
rect 376024 623766 376076 623772
rect 374644 601724 374696 601730
rect 374644 601666 374696 601672
rect 368388 596828 368440 596834
rect 368388 596770 368440 596776
rect 368400 596174 368428 596770
rect 368400 596146 368520 596174
rect 368492 589354 368520 596146
rect 371976 590708 372028 590714
rect 371976 590650 372028 590656
rect 368480 589348 368532 589354
rect 368480 589290 368532 589296
rect 370504 579692 370556 579698
rect 370504 579634 370556 579640
rect 367744 568608 367796 568614
rect 367744 568550 367796 568556
rect 366364 385076 366416 385082
rect 366364 385018 366416 385024
rect 365076 385008 365128 385014
rect 365076 384950 365128 384956
rect 365168 298104 365220 298110
rect 365168 298046 365220 298052
rect 365076 297832 365128 297838
rect 365076 297774 365128 297780
rect 364984 31680 365036 31686
rect 364984 31622 365036 31628
rect 363788 31204 363840 31210
rect 363788 31146 363840 31152
rect 363696 20664 363748 20670
rect 363696 20606 363748 20612
rect 363604 4140 363656 4146
rect 363604 4082 363656 4088
rect 365088 3874 365116 297774
rect 365076 3868 365128 3874
rect 365076 3810 365128 3816
rect 365180 3777 365208 298046
rect 365536 297696 365588 297702
rect 365536 297638 365588 297644
rect 365260 297628 365312 297634
rect 365260 297570 365312 297576
rect 365272 39710 365300 297570
rect 365444 297492 365496 297498
rect 365444 297434 365496 297440
rect 365352 297356 365404 297362
rect 365352 297298 365404 297304
rect 365260 39704 365312 39710
rect 365260 39646 365312 39652
rect 365364 39370 365392 297298
rect 365456 39574 365484 297434
rect 365548 39642 365576 297638
rect 365720 162240 365772 162246
rect 365720 162182 365772 162188
rect 365732 155922 365760 162182
rect 365720 155916 365772 155922
rect 365720 155858 365772 155864
rect 365536 39636 365588 39642
rect 365536 39578 365588 39584
rect 365444 39568 365496 39574
rect 365444 39510 365496 39516
rect 365352 39364 365404 39370
rect 365352 39306 365404 39312
rect 366376 30938 366404 385018
rect 367756 378146 367784 568550
rect 367744 378140 367796 378146
rect 367744 378082 367796 378088
rect 370516 378078 370544 579634
rect 371884 386572 371936 386578
rect 371884 386514 371936 386520
rect 370504 378072 370556 378078
rect 370504 378014 370556 378020
rect 370502 305688 370558 305697
rect 370502 305623 370558 305632
rect 368296 300620 368348 300626
rect 368296 300562 368348 300568
rect 368112 300144 368164 300150
rect 368018 300112 368074 300121
rect 368112 300086 368164 300092
rect 368018 300047 368074 300056
rect 367836 298036 367888 298042
rect 367836 297978 367888 297984
rect 366640 295248 366692 295254
rect 366640 295190 366692 295196
rect 366456 295112 366508 295118
rect 366456 295054 366508 295060
rect 366468 36718 366496 295054
rect 366548 294568 366600 294574
rect 366548 294510 366600 294516
rect 366560 36854 366588 294510
rect 366652 36990 366680 295190
rect 366732 294908 366784 294914
rect 366732 294850 366784 294856
rect 366640 36984 366692 36990
rect 366640 36926 366692 36932
rect 366744 36922 366772 294850
rect 367744 196648 367796 196654
rect 367744 196590 367796 196596
rect 367756 160750 367784 196590
rect 367744 160744 367796 160750
rect 367744 160686 367796 160692
rect 367744 106344 367796 106350
rect 367744 106286 367796 106292
rect 366732 36916 366784 36922
rect 366732 36858 366784 36864
rect 366548 36848 366600 36854
rect 366548 36790 366600 36796
rect 366456 36712 366508 36718
rect 366456 36654 366508 36660
rect 366364 30932 366416 30938
rect 366364 30874 366416 30880
rect 367756 7614 367784 106286
rect 367744 7608 367796 7614
rect 367744 7550 367796 7556
rect 365166 3768 365222 3777
rect 365166 3703 365222 3712
rect 361212 3324 361264 3330
rect 361212 3266 361264 3272
rect 360936 3256 360988 3262
rect 360936 3198 360988 3204
rect 367848 2174 367876 297978
rect 367928 297900 367980 297906
rect 367928 297842 367980 297848
rect 367940 3670 367968 297842
rect 368032 39438 368060 300047
rect 368124 39506 368152 300086
rect 368204 294500 368256 294506
rect 368204 294442 368256 294448
rect 368112 39500 368164 39506
rect 368112 39442 368164 39448
rect 368020 39432 368072 39438
rect 368020 39374 368072 39380
rect 368216 36786 368244 294442
rect 368308 42158 368336 300562
rect 369216 295316 369268 295322
rect 369216 295258 369268 295264
rect 369124 295180 369176 295186
rect 369124 295122 369176 295128
rect 368296 42152 368348 42158
rect 368296 42094 368348 42100
rect 369136 37058 369164 295122
rect 369228 37126 369256 295258
rect 369308 294976 369360 294982
rect 369308 294918 369360 294924
rect 369320 37194 369348 294918
rect 369400 286340 369452 286346
rect 369400 286282 369452 286288
rect 369308 37188 369360 37194
rect 369308 37130 369360 37136
rect 369216 37120 369268 37126
rect 369216 37062 369268 37068
rect 369124 37052 369176 37058
rect 369124 36994 369176 37000
rect 368204 36780 368256 36786
rect 368204 36722 368256 36728
rect 369412 31278 369440 286282
rect 369400 31272 369452 31278
rect 369400 31214 369452 31220
rect 367928 3664 367980 3670
rect 370516 3641 370544 305623
rect 370872 300416 370924 300422
rect 370872 300358 370924 300364
rect 370686 300248 370742 300257
rect 370686 300183 370742 300192
rect 370780 300212 370832 300218
rect 370596 289128 370648 289134
rect 370596 289070 370648 289076
rect 370608 31618 370636 289070
rect 370596 31612 370648 31618
rect 370596 31554 370648 31560
rect 370700 4049 370728 300183
rect 370780 300154 370832 300160
rect 370792 41954 370820 300154
rect 370884 42702 370912 300358
rect 371056 300348 371108 300354
rect 371056 300290 371108 300296
rect 370964 300280 371016 300286
rect 370964 300222 371016 300228
rect 370976 42770 371004 300222
rect 370964 42764 371016 42770
rect 370964 42706 371016 42712
rect 370872 42696 370924 42702
rect 370872 42638 370924 42644
rect 371068 42022 371096 300290
rect 371056 42016 371108 42022
rect 371056 41958 371108 41964
rect 370780 41948 370832 41954
rect 370780 41890 370832 41896
rect 371896 36446 371924 386514
rect 371988 379506 372016 590650
rect 372804 589280 372856 589286
rect 372804 589222 372856 589228
rect 372816 584458 372844 589222
rect 372804 584452 372856 584458
rect 372804 584394 372856 584400
rect 371976 379500 372028 379506
rect 371976 379442 372028 379448
rect 374656 379438 374684 601666
rect 376036 380866 376064 623766
rect 378796 382226 378824 645866
rect 379520 584452 379572 584458
rect 379520 584394 379572 584400
rect 379532 582690 379560 584394
rect 379520 582684 379572 582690
rect 379520 582626 379572 582632
rect 381556 383654 381584 667898
rect 381636 582684 381688 582690
rect 381636 582626 381688 582632
rect 381648 559366 381676 582626
rect 381636 559360 381688 559366
rect 381636 559302 381688 559308
rect 383752 559360 383804 559366
rect 383752 559302 383804 559308
rect 383764 554198 383792 559302
rect 383752 554192 383804 554198
rect 383752 554134 383804 554140
rect 385684 554192 385736 554198
rect 385684 554134 385736 554140
rect 385696 550594 385724 554134
rect 385684 550588 385736 550594
rect 385684 550530 385736 550536
rect 387432 550588 387484 550594
rect 387432 550530 387484 550536
rect 387444 546514 387472 550530
rect 387432 546508 387484 546514
rect 387432 546450 387484 546456
rect 388444 546508 388496 546514
rect 388444 546450 388496 546456
rect 388456 535498 388484 546450
rect 388444 535492 388496 535498
rect 388444 535434 388496 535440
rect 389824 535492 389876 535498
rect 389824 535434 389876 535440
rect 389836 524550 389864 535434
rect 389824 524544 389876 524550
rect 389824 524486 389876 524492
rect 391204 524544 391256 524550
rect 391204 524486 391256 524492
rect 391216 517546 391244 524486
rect 391204 517540 391256 517546
rect 391204 517482 391256 517488
rect 394608 517472 394660 517478
rect 394608 517414 394660 517420
rect 394620 513346 394648 517414
rect 394620 513318 394740 513346
rect 394712 510678 394740 513318
rect 394700 510672 394752 510678
rect 394700 510614 394752 510620
rect 382924 458244 382976 458250
rect 382924 458186 382976 458192
rect 381544 383648 381596 383654
rect 381544 383590 381596 383596
rect 378784 382220 378836 382226
rect 378784 382162 378836 382168
rect 376024 380860 376076 380866
rect 376024 380802 376076 380808
rect 374644 379432 374696 379438
rect 374644 379374 374696 379380
rect 382936 371210 382964 458186
rect 382924 371204 382976 371210
rect 382924 371146 382976 371152
rect 394700 351960 394752 351966
rect 394700 351902 394752 351908
rect 389824 347812 389876 347818
rect 389824 347754 389876 347760
rect 385960 338156 386012 338162
rect 385960 338098 386012 338104
rect 381636 306332 381688 306338
rect 381636 306274 381688 306280
rect 381544 305924 381596 305930
rect 381544 305866 381596 305872
rect 374644 305856 374696 305862
rect 374644 305798 374696 305804
rect 373264 302932 373316 302938
rect 373264 302874 373316 302880
rect 371976 298784 372028 298790
rect 371976 298726 372028 298732
rect 371884 36440 371936 36446
rect 371884 36382 371936 36388
rect 370686 4040 370742 4049
rect 370686 3975 370742 3984
rect 371988 3942 372016 298726
rect 372252 291916 372304 291922
rect 372252 291858 372304 291864
rect 372158 291816 372214 291825
rect 372158 291751 372214 291760
rect 372068 286408 372120 286414
rect 372068 286350 372120 286356
rect 372080 28286 372108 286350
rect 372172 36582 372200 291751
rect 372264 37262 372292 291858
rect 372344 291848 372396 291854
rect 372344 291790 372396 291796
rect 372252 37256 372304 37262
rect 372252 37198 372304 37204
rect 372160 36576 372212 36582
rect 372160 36518 372212 36524
rect 372356 36514 372384 291790
rect 373276 42634 373304 302874
rect 373632 300756 373684 300762
rect 373632 300698 373684 300704
rect 373540 300552 373592 300558
rect 373540 300494 373592 300500
rect 373448 300484 373500 300490
rect 373448 300426 373500 300432
rect 373356 289196 373408 289202
rect 373356 289138 373408 289144
rect 373264 42628 373316 42634
rect 373264 42570 373316 42576
rect 372344 36508 372396 36514
rect 372344 36450 372396 36456
rect 373368 31550 373396 289138
rect 373460 42566 373488 300426
rect 373448 42560 373500 42566
rect 373448 42502 373500 42508
rect 373552 42498 373580 300494
rect 373540 42492 373592 42498
rect 373540 42434 373592 42440
rect 373644 42430 373672 300698
rect 373632 42424 373684 42430
rect 373632 42366 373684 42372
rect 373356 31544 373408 31550
rect 373356 31486 373408 31492
rect 372068 28280 372120 28286
rect 372068 28222 372120 28228
rect 374656 6866 374684 305798
rect 378692 303612 378744 303618
rect 378692 303554 378744 303560
rect 376024 303408 376076 303414
rect 376024 303350 376076 303356
rect 375104 292528 375156 292534
rect 375104 292470 375156 292476
rect 375012 292120 375064 292126
rect 375012 292062 375064 292068
rect 374736 292052 374788 292058
rect 374736 291994 374788 292000
rect 374644 6860 374696 6866
rect 374644 6802 374696 6808
rect 371976 3936 372028 3942
rect 371976 3878 372028 3884
rect 367928 3606 367980 3612
rect 370502 3632 370558 3641
rect 370502 3567 370558 3576
rect 374748 3534 374776 291994
rect 374920 291984 374972 291990
rect 374920 291926 374972 291932
rect 374828 286476 374880 286482
rect 374828 286418 374880 286424
rect 374840 28354 374868 286418
rect 374932 33930 374960 291926
rect 374920 33924 374972 33930
rect 374920 33866 374972 33872
rect 375024 33862 375052 292062
rect 375116 36650 375144 292470
rect 375104 36644 375156 36650
rect 375104 36586 375156 36592
rect 375012 33856 375064 33862
rect 375012 33798 375064 33804
rect 376036 31414 376064 303350
rect 376208 303204 376260 303210
rect 376208 303146 376260 303152
rect 376114 302968 376170 302977
rect 376114 302903 376170 302912
rect 376128 42090 376156 302903
rect 376220 42226 376248 303146
rect 376300 300824 376352 300830
rect 376300 300766 376352 300772
rect 376312 42294 376340 300766
rect 376392 300688 376444 300694
rect 376392 300630 376444 300636
rect 376404 42362 376432 300630
rect 376484 300076 376536 300082
rect 376484 300018 376536 300024
rect 376496 44674 376524 300018
rect 378600 300008 378652 300014
rect 378600 299950 378652 299956
rect 376668 299940 376720 299946
rect 376668 299882 376720 299888
rect 376576 298852 376628 298858
rect 376576 298794 376628 298800
rect 376588 45490 376616 298794
rect 376680 46306 376708 299882
rect 377588 292256 377640 292262
rect 377588 292198 377640 292204
rect 377404 292188 377456 292194
rect 377404 292130 377456 292136
rect 376668 46300 376720 46306
rect 376668 46242 376720 46248
rect 376576 45484 376628 45490
rect 376576 45426 376628 45432
rect 376484 44668 376536 44674
rect 376484 44610 376536 44616
rect 376392 42356 376444 42362
rect 376392 42298 376444 42304
rect 376300 42288 376352 42294
rect 376300 42230 376352 42236
rect 376208 42220 376260 42226
rect 376208 42162 376260 42168
rect 376116 42084 376168 42090
rect 376116 42026 376168 42032
rect 376024 31408 376076 31414
rect 376024 31350 376076 31356
rect 374828 28348 374880 28354
rect 374828 28290 374880 28296
rect 377416 3602 377444 292130
rect 377496 286612 377548 286618
rect 377496 286554 377548 286560
rect 377508 28422 377536 286554
rect 377600 33998 377628 292198
rect 377680 291780 377732 291786
rect 377680 291722 377732 291728
rect 377588 33992 377640 33998
rect 377588 33934 377640 33940
rect 377692 33794 377720 291722
rect 378612 46617 378640 299950
rect 378598 46608 378654 46617
rect 378598 46543 378654 46552
rect 378704 46442 378732 303554
rect 379060 303476 379112 303482
rect 379060 303418 379112 303424
rect 378968 303000 379020 303006
rect 378968 302942 379020 302948
rect 378784 301572 378836 301578
rect 378784 301514 378836 301520
rect 378692 46436 378744 46442
rect 378692 46378 378744 46384
rect 377680 33788 377732 33794
rect 377680 33730 377732 33736
rect 378796 33114 378824 301514
rect 378876 289332 378928 289338
rect 378876 289274 378928 289280
rect 378784 33108 378836 33114
rect 378784 33050 378836 33056
rect 378888 31346 378916 289274
rect 378980 45354 379008 302942
rect 378968 45348 379020 45354
rect 378968 45290 379020 45296
rect 379072 44742 379100 303418
rect 379244 303340 379296 303346
rect 379244 303282 379296 303288
rect 379152 303068 379204 303074
rect 379152 303010 379204 303016
rect 379164 44810 379192 303010
rect 379256 45286 379284 303282
rect 379336 303136 379388 303142
rect 379336 303078 379388 303084
rect 379244 45280 379296 45286
rect 379244 45222 379296 45228
rect 379348 45218 379376 303078
rect 379428 302864 379480 302870
rect 379428 302806 379480 302812
rect 379440 46510 379468 302806
rect 381452 302796 381504 302802
rect 381452 302738 381504 302744
rect 380164 292392 380216 292398
rect 380164 292334 380216 292340
rect 379428 46504 379480 46510
rect 379428 46446 379480 46452
rect 379336 45212 379388 45218
rect 379336 45154 379388 45160
rect 379152 44804 379204 44810
rect 379152 44746 379204 44752
rect 379060 44736 379112 44742
rect 379060 44678 379112 44684
rect 380176 34134 380204 292334
rect 380256 292324 380308 292330
rect 380256 292266 380308 292272
rect 380164 34128 380216 34134
rect 380164 34070 380216 34076
rect 380268 34066 380296 292266
rect 380440 289672 380492 289678
rect 380440 289614 380492 289620
rect 380348 289536 380400 289542
rect 380348 289478 380400 289484
rect 380360 34270 380388 289478
rect 380452 34406 380480 289614
rect 381360 160200 381412 160206
rect 381360 160142 381412 160148
rect 381372 84182 381400 160142
rect 381360 84176 381412 84182
rect 381360 84118 381412 84124
rect 381464 46578 381492 302738
rect 381452 46572 381504 46578
rect 381452 46514 381504 46520
rect 381556 45558 381584 305866
rect 381648 46714 381676 306274
rect 385868 306264 385920 306270
rect 384486 306232 384542 306241
rect 385868 306206 385920 306212
rect 384486 306167 384542 306176
rect 384580 306196 384632 306202
rect 381728 306128 381780 306134
rect 381728 306070 381780 306076
rect 384302 306096 384358 306105
rect 381636 46708 381688 46714
rect 381636 46650 381688 46656
rect 381740 46646 381768 306070
rect 384302 306031 384358 306040
rect 382004 303544 382056 303550
rect 382004 303486 382056 303492
rect 381910 303104 381966 303113
rect 381910 303039 381966 303048
rect 381820 292460 381872 292466
rect 381820 292402 381872 292408
rect 381728 46640 381780 46646
rect 381728 46582 381780 46588
rect 381544 45552 381596 45558
rect 381544 45494 381596 45500
rect 380440 34400 380492 34406
rect 380440 34342 380492 34348
rect 380348 34264 380400 34270
rect 380348 34206 380400 34212
rect 381832 34202 381860 292402
rect 381924 45014 381952 303039
rect 382016 45082 382044 303486
rect 382096 303272 382148 303278
rect 382096 303214 382148 303220
rect 382186 303240 382242 303249
rect 382108 45150 382136 303214
rect 382186 303175 382242 303184
rect 382096 45144 382148 45150
rect 382096 45086 382148 45092
rect 382004 45076 382056 45082
rect 382004 45018 382056 45024
rect 381912 45008 381964 45014
rect 381912 44950 381964 44956
rect 382200 44946 382228 303175
rect 382924 297288 382976 297294
rect 382924 297230 382976 297236
rect 382188 44940 382240 44946
rect 382188 44882 382240 44888
rect 381820 34196 381872 34202
rect 381820 34138 381872 34144
rect 380256 34060 380308 34066
rect 380256 34002 380308 34008
rect 378876 31340 378928 31346
rect 378876 31282 378928 31288
rect 377496 28416 377548 28422
rect 377496 28358 377548 28364
rect 382936 3738 382964 297230
rect 383200 289808 383252 289814
rect 383200 289750 383252 289756
rect 383016 289468 383068 289474
rect 383016 289410 383068 289416
rect 382924 3732 382976 3738
rect 382924 3674 382976 3680
rect 377404 3596 377456 3602
rect 377404 3538 377456 3544
rect 374736 3528 374788 3534
rect 383028 3505 383056 289410
rect 383108 289400 383160 289406
rect 383108 289342 383160 289348
rect 383120 34474 383148 289342
rect 383108 34468 383160 34474
rect 383108 34410 383160 34416
rect 383212 34338 383240 289750
rect 383292 289604 383344 289610
rect 383292 289546 383344 289552
rect 383200 34332 383252 34338
rect 383200 34274 383252 34280
rect 383304 33726 383332 289546
rect 383384 160132 383436 160138
rect 383384 160074 383436 160080
rect 383396 73166 383424 160074
rect 383384 73160 383436 73166
rect 383384 73102 383436 73108
rect 384212 51128 384264 51134
rect 384212 51070 384264 51076
rect 383292 33720 383344 33726
rect 383292 33662 383344 33668
rect 384224 31686 384252 51070
rect 384212 31680 384264 31686
rect 384212 31622 384264 31628
rect 374736 3470 374788 3476
rect 383014 3496 383070 3505
rect 383014 3431 383070 3440
rect 367836 2168 367888 2174
rect 367836 2110 367888 2116
rect 384316 2106 384344 306031
rect 384396 305584 384448 305590
rect 384396 305526 384448 305532
rect 384408 46374 384436 305526
rect 384396 46368 384448 46374
rect 384396 46310 384448 46316
rect 384500 3369 384528 306167
rect 384580 306138 384632 306144
rect 384592 46782 384620 306138
rect 384764 306060 384816 306066
rect 384764 306002 384816 306008
rect 384670 305960 384726 305969
rect 384670 305895 384726 305904
rect 384580 46776 384632 46782
rect 384580 46718 384632 46724
rect 384684 44878 384712 305895
rect 384776 46753 384804 306002
rect 384856 305992 384908 305998
rect 384856 305934 384908 305940
rect 384868 47025 384896 305934
rect 385776 305516 385828 305522
rect 385776 305458 385828 305464
rect 385684 304428 385736 304434
rect 385684 304370 385736 304376
rect 384948 286544 385000 286550
rect 384948 286486 385000 286492
rect 384854 47016 384910 47025
rect 384854 46951 384910 46960
rect 384762 46744 384818 46753
rect 384762 46679 384818 46688
rect 384672 44872 384724 44878
rect 384672 44814 384724 44820
rect 384960 31142 384988 286486
rect 384948 31136 385000 31142
rect 384948 31078 385000 31084
rect 385696 3466 385724 304370
rect 385788 46889 385816 305458
rect 385774 46880 385830 46889
rect 385880 46850 385908 306206
rect 385972 293962 386000 338098
rect 386144 302728 386196 302734
rect 386144 302670 386196 302676
rect 385960 293956 386012 293962
rect 385960 293898 386012 293904
rect 385960 289060 386012 289066
rect 385960 289002 386012 289008
rect 385774 46815 385830 46824
rect 385868 46844 385920 46850
rect 385868 46786 385920 46792
rect 385972 31074 386000 289002
rect 386052 288992 386104 288998
rect 386052 288934 386104 288940
rect 386064 31482 386092 288934
rect 386156 46918 386184 302670
rect 386236 289740 386288 289746
rect 386236 289682 386288 289688
rect 386144 46912 386196 46918
rect 386144 46854 386196 46860
rect 386248 33658 386276 289682
rect 389836 162178 389864 347754
rect 392584 193860 392636 193866
rect 392584 193802 392636 193808
rect 392596 182170 392624 193802
rect 389916 182164 389968 182170
rect 389916 182106 389968 182112
rect 392584 182164 392636 182170
rect 392584 182106 392636 182112
rect 389928 167686 389956 182106
rect 389916 167680 389968 167686
rect 389916 167622 389968 167628
rect 390560 164892 390612 164898
rect 390560 164834 390612 164840
rect 390572 162246 390600 164834
rect 390560 162240 390612 162246
rect 390560 162182 390612 162188
rect 389824 162172 389876 162178
rect 389824 162114 389876 162120
rect 386328 160268 386380 160274
rect 386328 160210 386380 160216
rect 386340 62082 386368 160210
rect 388444 140072 388496 140078
rect 388444 140014 388496 140020
rect 388456 124914 388484 140014
rect 388444 124908 388496 124914
rect 388444 124850 388496 124856
rect 389836 106350 389864 162114
rect 394712 113174 394740 351902
rect 397472 336122 397500 703520
rect 406384 656940 406436 656946
rect 406384 656882 406436 656888
rect 402244 510604 402296 510610
rect 402244 510546 402296 510552
rect 402256 469334 402284 510546
rect 402244 469328 402296 469334
rect 402244 469270 402296 469276
rect 405004 469328 405056 469334
rect 405004 469270 405056 469276
rect 405016 455394 405044 469270
rect 405004 455388 405056 455394
rect 405004 455330 405056 455336
rect 406396 383586 406424 656882
rect 407764 634840 407816 634846
rect 407764 634782 407816 634788
rect 406476 455388 406528 455394
rect 406476 455330 406528 455336
rect 406488 450974 406516 455330
rect 406476 450968 406528 450974
rect 406476 450910 406528 450916
rect 406384 383580 406436 383586
rect 406384 383522 406436 383528
rect 407776 382158 407804 634782
rect 410524 612808 410576 612814
rect 410524 612750 410576 612756
rect 408500 450968 408552 450974
rect 408500 450910 408552 450916
rect 408512 441658 408540 450910
rect 408500 441652 408552 441658
rect 408500 441594 408552 441600
rect 407764 382152 407816 382158
rect 407764 382094 407816 382100
rect 410536 380798 410564 612750
rect 411904 524476 411956 524482
rect 411904 524418 411956 524424
rect 410524 380792 410576 380798
rect 410524 380734 410576 380740
rect 411916 375290 411944 524418
rect 411904 375284 411956 375290
rect 411904 375226 411956 375232
rect 405740 350600 405792 350606
rect 405740 350542 405792 350548
rect 401600 342916 401652 342922
rect 401600 342858 401652 342864
rect 399484 339516 399536 339522
rect 399484 339458 399536 339464
rect 397460 336116 397512 336122
rect 397460 336058 397512 336064
rect 399496 315994 399524 339458
rect 401612 334914 401640 342858
rect 401612 334886 402086 334914
rect 405752 334900 405780 350542
rect 412652 348430 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 429856 700806 429884 703520
rect 429844 700800 429896 700806
rect 429844 700742 429896 700748
rect 445116 700800 445168 700806
rect 445116 700742 445168 700748
rect 445024 700732 445076 700738
rect 445024 700674 445076 700680
rect 416044 700460 416096 700466
rect 416044 700402 416096 700408
rect 444288 700460 444340 700466
rect 444288 700402 444340 700408
rect 414664 513392 414716 513398
rect 414664 513334 414716 513340
rect 413744 441584 413796 441590
rect 413744 441526 413796 441532
rect 413756 437578 413784 441526
rect 413744 437572 413796 437578
rect 413744 437514 413796 437520
rect 414676 373998 414704 513334
rect 414756 437572 414808 437578
rect 414756 437514 414808 437520
rect 414768 431390 414796 437514
rect 414756 431384 414808 431390
rect 414756 431326 414808 431332
rect 414664 373992 414716 373998
rect 414664 373934 414716 373940
rect 412640 348424 412692 348430
rect 412640 348366 412692 348372
rect 416056 336258 416084 700402
rect 416228 685228 416280 685234
rect 416228 685170 416280 685176
rect 416136 683528 416188 683534
rect 416136 683470 416188 683476
rect 416044 336252 416096 336258
rect 416044 336194 416096 336200
rect 409420 335436 409472 335442
rect 409420 335378 409472 335384
rect 409432 334900 409460 335378
rect 413100 335368 413152 335374
rect 413100 335310 413152 335316
rect 413112 334900 413140 335310
rect 416148 334966 416176 683470
rect 416240 336394 416268 685170
rect 419356 685160 419408 685166
rect 419356 685102 419408 685108
rect 418804 684752 418856 684758
rect 418804 684694 418856 684700
rect 416320 502376 416372 502382
rect 416320 502318 416372 502324
rect 416332 373930 416360 502318
rect 418712 480276 418764 480282
rect 418712 480218 418764 480224
rect 417424 469260 417476 469266
rect 417424 469202 417476 469208
rect 416688 431384 416740 431390
rect 416688 431326 416740 431332
rect 416700 429078 416728 431326
rect 416688 429072 416740 429078
rect 416688 429014 416740 429020
rect 416320 373924 416372 373930
rect 416320 373866 416372 373872
rect 417436 371142 417464 469202
rect 418620 436144 418672 436150
rect 418620 436086 418672 436092
rect 417424 371136 417476 371142
rect 417424 371078 417476 371084
rect 418632 369850 418660 436086
rect 418724 372502 418752 480218
rect 418712 372496 418764 372502
rect 418712 372438 418764 372444
rect 418620 369844 418672 369850
rect 418620 369786 418672 369792
rect 416780 336932 416832 336938
rect 416780 336874 416832 336880
rect 416228 336388 416280 336394
rect 416228 336330 416280 336336
rect 416136 334960 416188 334966
rect 416136 334902 416188 334908
rect 416792 334900 416820 336874
rect 418816 335034 418844 684694
rect 418988 684684 419040 684690
rect 418988 684626 419040 684632
rect 418896 684548 418948 684554
rect 418896 684490 418948 684496
rect 418804 335028 418856 335034
rect 418804 334970 418856 334976
rect 418908 334898 418936 684490
rect 418896 334892 418948 334898
rect 418896 334834 418948 334840
rect 419000 334694 419028 684626
rect 419080 684616 419132 684622
rect 419080 684558 419132 684564
rect 419092 334762 419120 684558
rect 419172 683460 419224 683466
rect 419172 683402 419224 683408
rect 419080 334756 419132 334762
rect 419080 334698 419132 334704
rect 418988 334688 419040 334694
rect 418988 334630 419040 334636
rect 419184 334626 419212 683402
rect 419264 683392 419316 683398
rect 419264 683334 419316 683340
rect 419276 334830 419304 683334
rect 419368 336190 419396 685102
rect 419448 684820 419500 684826
rect 419448 684762 419500 684768
rect 419460 336326 419488 684762
rect 420184 683324 420236 683330
rect 420184 683266 420236 683272
rect 419448 336320 419500 336326
rect 419448 336262 419500 336268
rect 419356 336184 419408 336190
rect 419356 336126 419408 336132
rect 420196 335102 420224 683266
rect 420274 682952 420330 682961
rect 420274 682887 420330 682896
rect 420184 335096 420236 335102
rect 420184 335038 420236 335044
rect 419264 334824 419316 334830
rect 419264 334766 419316 334772
rect 420090 334656 420146 334665
rect 419172 334620 419224 334626
rect 420288 334642 420316 682887
rect 420552 682712 420604 682718
rect 420552 682654 420604 682660
rect 420368 429072 420420 429078
rect 420368 429014 420420 429020
rect 420380 418198 420408 429014
rect 420368 418192 420420 418198
rect 420368 418134 420420 418140
rect 420564 345014 420592 682654
rect 436100 462460 436152 462466
rect 436100 462402 436152 462408
rect 433248 462392 433300 462398
rect 433248 462334 433300 462340
rect 422300 455456 422352 455462
rect 422300 455398 422352 455404
rect 422312 444394 422340 455398
rect 427452 447160 427504 447166
rect 427452 447102 427504 447108
rect 427464 444924 427492 447102
rect 433260 445806 433288 462334
rect 432420 445800 432472 445806
rect 432420 445742 432472 445748
rect 433248 445800 433300 445806
rect 433248 445742 433300 445748
rect 432432 444924 432460 445742
rect 436112 445738 436140 462402
rect 444104 445800 444156 445806
rect 444104 445742 444156 445748
rect 436100 445732 436152 445738
rect 436100 445674 436152 445680
rect 437388 445732 437440 445738
rect 437388 445674 437440 445680
rect 437400 444938 437428 445674
rect 437308 444924 437428 444938
rect 437308 444910 437414 444924
rect 437308 444582 437336 444910
rect 437296 444576 437348 444582
rect 437296 444518 437348 444524
rect 442382 444514 442672 444530
rect 442382 444508 442684 444514
rect 442382 444502 442632 444508
rect 442632 444450 442684 444456
rect 422760 444440 422812 444446
rect 422312 444388 422760 444394
rect 422312 444382 422812 444388
rect 422312 444366 422800 444382
rect 421484 417722 421512 420036
rect 421472 417716 421524 417722
rect 421472 417658 421524 417664
rect 422128 417450 422156 420036
rect 422312 420022 422786 420050
rect 422864 420022 423430 420050
rect 422116 417444 422168 417450
rect 422116 417386 422168 417392
rect 422312 389842 422340 420022
rect 422864 412634 422892 420022
rect 424060 417586 424088 420036
rect 424704 417654 424732 420036
rect 424692 417648 424744 417654
rect 424692 417590 424744 417596
rect 424048 417580 424100 417586
rect 424048 417522 424100 417528
rect 425348 417518 425376 420036
rect 425992 417790 426020 420036
rect 440884 418804 440936 418810
rect 440884 418746 440936 418752
rect 426440 418124 426492 418130
rect 426440 418066 426492 418072
rect 425980 417784 426032 417790
rect 425980 417726 426032 417732
rect 425336 417512 425388 417518
rect 425336 417454 425388 417460
rect 426452 415682 426480 418066
rect 436744 416084 436796 416090
rect 436744 416026 436796 416032
rect 426440 415676 426492 415682
rect 426440 415618 426492 415624
rect 429844 415676 429896 415682
rect 429844 415618 429896 415624
rect 422404 412606 422892 412634
rect 422404 391270 422432 412606
rect 429856 410242 429884 415618
rect 429844 410236 429896 410242
rect 429844 410178 429896 410184
rect 431224 410236 431276 410242
rect 431224 410178 431276 410184
rect 431236 398818 431264 410178
rect 431224 398812 431276 398818
rect 431224 398754 431276 398760
rect 432604 398812 432656 398818
rect 432604 398754 432656 398760
rect 432616 392018 432644 398754
rect 432604 392012 432656 392018
rect 432604 391954 432656 391960
rect 433984 392012 434036 392018
rect 433984 391954 434036 391960
rect 422392 391264 422444 391270
rect 422392 391206 422444 391212
rect 422300 389836 422352 389842
rect 422300 389778 422352 389784
rect 433996 371550 434024 391954
rect 433984 371544 434036 371550
rect 433984 371486 434036 371492
rect 435364 371544 435416 371550
rect 435364 371486 435416 371492
rect 429200 369912 429252 369918
rect 429200 369854 429252 369860
rect 429212 365702 429240 369854
rect 429200 365696 429252 365702
rect 429200 365638 429252 365644
rect 432604 362976 432656 362982
rect 432604 362918 432656 362924
rect 420564 344986 420776 345014
rect 420460 336796 420512 336802
rect 420460 336738 420512 336744
rect 420146 334614 420316 334642
rect 420472 334642 420500 336738
rect 420748 334801 420776 344986
rect 431224 338224 431276 338230
rect 431224 338166 431276 338172
rect 429936 336932 429988 336938
rect 429936 336874 429988 336880
rect 424140 336864 424192 336870
rect 424140 336806 424192 336812
rect 424152 334900 424180 336806
rect 420734 334792 420790 334801
rect 420734 334727 420790 334736
rect 420472 334628 420592 334642
rect 420486 334614 420592 334628
rect 420090 334591 420146 334600
rect 419172 334562 419224 334568
rect 420564 334506 420592 334614
rect 420734 334520 420790 334529
rect 420486 334478 420734 334506
rect 428094 334520 428150 334529
rect 427846 334478 428094 334506
rect 420734 334455 420790 334464
rect 428094 334455 428150 334464
rect 428108 334422 428136 334455
rect 428096 334416 428148 334422
rect 428096 334358 428148 334364
rect 429844 332648 429896 332654
rect 429844 332590 429896 332596
rect 399484 315988 399536 315994
rect 399484 315930 399536 315936
rect 426348 305788 426400 305794
rect 426348 305730 426400 305736
rect 407120 301504 407172 301510
rect 407120 301446 407172 301452
rect 406384 211812 406436 211818
rect 406384 211754 406436 211760
rect 398104 196716 398156 196722
rect 398104 196658 398156 196664
rect 398116 193866 398144 196658
rect 406396 196654 406424 211754
rect 406384 196648 406436 196654
rect 406384 196590 406436 196596
rect 398104 193860 398156 193866
rect 398104 193802 398156 193808
rect 405004 189780 405056 189786
rect 405004 189722 405056 189728
rect 405016 172582 405044 189722
rect 401600 172576 401652 172582
rect 401600 172518 401652 172524
rect 405004 172576 405056 172582
rect 405004 172518 405056 172524
rect 401612 169794 401640 172518
rect 397460 169788 397512 169794
rect 397460 169730 397512 169736
rect 401600 169788 401652 169794
rect 401600 169730 401652 169736
rect 397472 164898 397500 169730
rect 397460 164892 397512 164898
rect 397460 164834 397512 164840
rect 403624 161560 403676 161566
rect 403624 161502 403676 161508
rect 402336 153264 402388 153270
rect 402336 153206 402388 153212
rect 402348 147694 402376 153206
rect 399484 147688 399536 147694
rect 399484 147630 399536 147636
rect 402336 147688 402388 147694
rect 402336 147630 402388 147636
rect 399496 140078 399524 147630
rect 399484 140072 399536 140078
rect 399484 140014 399536 140020
rect 403636 139398 403664 161502
rect 406384 160336 406436 160342
rect 406384 160278 406436 160284
rect 405648 156120 405700 156126
rect 405648 156062 405700 156068
rect 405660 153270 405688 156062
rect 405648 153264 405700 153270
rect 405648 153206 405700 153212
rect 403624 139392 403676 139398
rect 403624 139334 403676 139340
rect 406396 117298 406424 160278
rect 406384 117292 406436 117298
rect 406384 117234 406436 117240
rect 407132 113174 407160 301446
rect 419448 233912 419500 233918
rect 419448 233854 419500 233860
rect 416044 221468 416096 221474
rect 416044 221410 416096 221416
rect 411260 206304 411312 206310
rect 411260 206246 411312 206252
rect 411272 171134 411300 206246
rect 411272 171106 411392 171134
rect 410524 161696 410576 161702
rect 410524 161638 410576 161644
rect 407764 161628 407816 161634
rect 407764 161570 407816 161576
rect 407396 159452 407448 159458
rect 407396 159394 407448 159400
rect 407408 156126 407436 159394
rect 407396 156120 407448 156126
rect 407396 156062 407448 156068
rect 407776 128314 407804 161570
rect 407764 128308 407816 128314
rect 407764 128250 407816 128256
rect 394712 113146 395292 113174
rect 407132 113146 407620 113174
rect 389824 106344 389876 106350
rect 389824 106286 389876 106292
rect 389836 104938 389864 106286
rect 389528 104910 389864 104938
rect 395264 104938 395292 113146
rect 402152 106956 402204 106962
rect 402152 106898 402204 106904
rect 402164 104938 402192 106898
rect 395264 104910 395692 104938
rect 401856 104910 402192 104938
rect 407592 104938 407620 113146
rect 410536 105602 410564 161638
rect 410616 160404 410668 160410
rect 410616 160346 410668 160352
rect 410628 106282 410656 160346
rect 411364 159882 411392 171106
rect 416056 163946 416084 221410
rect 417424 200796 417476 200802
rect 417424 200738 417476 200744
rect 416136 194744 416188 194750
rect 416136 194686 416188 194692
rect 416148 189786 416176 194686
rect 416136 189780 416188 189786
rect 416136 189722 416188 189728
rect 417436 180130 417464 200738
rect 417424 180124 417476 180130
rect 417424 180066 417476 180072
rect 414756 163940 414808 163946
rect 414756 163882 414808 163888
rect 416044 163940 416096 163946
rect 416044 163882 416096 163888
rect 414768 160274 414796 163882
rect 414756 160268 414808 160274
rect 414756 160210 414808 160216
rect 414768 159882 414796 160210
rect 419460 160138 419488 233854
rect 424324 227792 424376 227798
rect 424324 227734 424376 227740
rect 423036 216708 423088 216714
rect 423036 216650 423088 216656
rect 422944 213172 422996 213178
rect 422944 213114 422996 213120
rect 420184 209840 420236 209846
rect 420184 209782 420236 209788
rect 419540 201544 419592 201550
rect 419540 201486 419592 201492
rect 419552 196722 419580 201486
rect 419540 196716 419592 196722
rect 419540 196658 419592 196664
rect 420196 194750 420224 209782
rect 422956 201550 422984 213114
rect 423048 211818 423076 216650
rect 423036 211812 423088 211818
rect 423036 211754 423088 211760
rect 424336 209846 424364 227734
rect 424324 209840 424376 209846
rect 424324 209782 424376 209788
rect 422944 201544 422996 201550
rect 422944 201486 422996 201492
rect 420184 194744 420236 194750
rect 420184 194686 420236 194692
rect 421746 162752 421802 162761
rect 421746 162687 421802 162696
rect 421760 161770 421788 162687
rect 426360 161906 426388 305730
rect 428464 232552 428516 232558
rect 428464 232494 428516 232500
rect 427820 217592 427872 217598
rect 427820 217534 427872 217540
rect 427832 213178 427860 217534
rect 428476 216714 428504 232494
rect 428464 216708 428516 216714
rect 428464 216650 428516 216656
rect 427820 213172 427872 213178
rect 427820 213114 427872 213120
rect 428464 209840 428516 209846
rect 428464 209782 428516 209788
rect 425060 161900 425112 161906
rect 425060 161842 425112 161848
rect 426348 161900 426400 161906
rect 426348 161842 426400 161848
rect 421748 161764 421800 161770
rect 421748 161706 421800 161712
rect 420920 160744 420972 160750
rect 420920 160686 420972 160692
rect 418390 160132 418442 160138
rect 418390 160074 418442 160080
rect 419448 160132 419500 160138
rect 419448 160074 419500 160080
rect 411364 159854 411792 159882
rect 414768 159854 415104 159882
rect 418402 159868 418430 160074
rect 420932 159526 420960 160686
rect 421760 160206 421788 161706
rect 425072 161702 425100 161842
rect 425060 161696 425112 161702
rect 425060 161638 425112 161644
rect 421380 160200 421432 160206
rect 421380 160142 421432 160148
rect 421748 160200 421800 160206
rect 425072 160154 425100 161638
rect 428476 160750 428504 209782
rect 429856 194546 429884 332590
rect 429948 325650 429976 336874
rect 429936 325644 429988 325650
rect 429936 325586 429988 325592
rect 431236 282878 431264 338166
rect 431408 336864 431460 336870
rect 431408 336806 431460 336812
rect 431316 335436 431368 335442
rect 431316 335378 431368 335384
rect 431328 323610 431356 335378
rect 431420 326398 431448 336806
rect 432616 332897 432644 362918
rect 435376 360262 435404 371486
rect 436756 369782 436784 416026
rect 439504 414044 439556 414050
rect 439504 413986 439556 413992
rect 436744 369776 436796 369782
rect 436744 369718 436796 369724
rect 439516 368490 439544 413986
rect 439504 368484 439556 368490
rect 439504 368426 439556 368432
rect 440896 368422 440924 418746
rect 442264 403028 442316 403034
rect 442264 402970 442316 402976
rect 440976 392080 441028 392086
rect 440976 392022 441028 392028
rect 440884 368416 440936 368422
rect 440884 368358 440936 368364
rect 440988 367062 441016 392022
rect 440976 367056 441028 367062
rect 440976 366998 441028 367004
rect 442276 366994 442304 402970
rect 442356 380928 442408 380934
rect 442356 380870 442408 380876
rect 442264 366988 442316 366994
rect 442264 366930 442316 366936
rect 442368 365634 442396 380870
rect 442356 365628 442408 365634
rect 442356 365570 442408 365576
rect 436928 363044 436980 363050
rect 436928 362986 436980 362992
rect 435548 360324 435600 360330
rect 435548 360266 435600 360272
rect 435364 360256 435416 360262
rect 435364 360198 435416 360204
rect 432696 344344 432748 344350
rect 432696 344286 432748 344292
rect 432602 332888 432658 332897
rect 432602 332823 432658 332832
rect 432604 330540 432656 330546
rect 432604 330482 432656 330488
rect 432420 329724 432472 329730
rect 432420 329666 432472 329672
rect 432432 329225 432460 329666
rect 432418 329216 432474 329225
rect 432418 329151 432474 329160
rect 431868 327752 431920 327758
rect 431868 327694 431920 327700
rect 431408 326392 431460 326398
rect 431408 326334 431460 326340
rect 431316 323604 431368 323610
rect 431316 323546 431368 323552
rect 431224 282872 431276 282878
rect 431224 282814 431276 282820
rect 429936 254924 429988 254930
rect 429936 254866 429988 254872
rect 429948 227798 429976 254866
rect 429936 227792 429988 227798
rect 429936 227734 429988 227740
rect 429844 194540 429896 194546
rect 429844 194482 429896 194488
rect 428646 162752 428702 162761
rect 428646 162687 428702 162696
rect 428660 161838 428688 162687
rect 428648 161832 428700 161838
rect 428648 161774 428700 161780
rect 428464 160744 428516 160750
rect 428464 160686 428516 160692
rect 428004 160404 428056 160410
rect 428004 160346 428056 160352
rect 421748 160142 421800 160148
rect 421392 159610 421420 160142
rect 425026 160126 425100 160154
rect 425026 159868 425054 160126
rect 428016 159882 428044 160346
rect 428660 159882 428688 161774
rect 431880 161702 431908 327694
rect 432616 310865 432644 330482
rect 432708 325553 432736 344286
rect 435456 335436 435508 335442
rect 435456 335378 435508 335384
rect 432880 331356 432932 331362
rect 432880 331298 432932 331304
rect 432788 328908 432840 328914
rect 432788 328850 432840 328856
rect 432694 325544 432750 325553
rect 432694 325479 432750 325488
rect 432800 318209 432828 328850
rect 432892 321881 432920 331298
rect 435364 329112 435416 329118
rect 435364 329054 435416 329060
rect 432878 321872 432934 321881
rect 432878 321807 432934 321816
rect 432786 318200 432842 318209
rect 432786 318135 432842 318144
rect 433248 314560 433300 314566
rect 433246 314528 433248 314537
rect 433300 314528 433302 314537
rect 433246 314463 433302 314472
rect 432602 310856 432658 310865
rect 432602 310791 432658 310800
rect 432236 307760 432288 307766
rect 432236 307702 432288 307708
rect 432248 307193 432276 307702
rect 432234 307184 432290 307193
rect 432234 307119 432290 307128
rect 431960 260364 432012 260370
rect 431960 260306 432012 260312
rect 431972 254930 432000 260306
rect 431960 254924 432012 254930
rect 431960 254866 432012 254872
rect 433984 230988 434036 230994
rect 433984 230930 434036 230936
rect 433996 217598 434024 230930
rect 433984 217592 434036 217598
rect 433984 217534 434036 217540
rect 434260 213036 434312 213042
rect 434260 212978 434312 212984
rect 434272 209846 434300 212978
rect 434260 209840 434312 209846
rect 434260 209782 434312 209788
rect 433248 203584 433300 203590
rect 433248 203526 433300 203532
rect 433260 200802 433288 203526
rect 433248 200796 433300 200802
rect 433248 200738 433300 200744
rect 435376 162858 435404 329054
rect 435468 249762 435496 335378
rect 435560 328914 435588 360266
rect 436836 358828 436888 358834
rect 436836 358770 436888 358776
rect 435640 348424 435692 348430
rect 435640 348366 435692 348372
rect 435548 328908 435600 328914
rect 435548 328850 435600 328856
rect 435652 319530 435680 348366
rect 435732 336796 435784 336802
rect 435732 336738 435784 336744
rect 435744 327078 435772 336738
rect 436744 331288 436796 331294
rect 436744 331230 436796 331236
rect 435732 327072 435784 327078
rect 435732 327014 435784 327020
rect 435640 319524 435692 319530
rect 435640 319466 435692 319472
rect 435456 249756 435508 249762
rect 435456 249698 435508 249704
rect 436756 183530 436784 331230
rect 436848 307766 436876 358770
rect 436940 329730 436968 362986
rect 442264 361684 442316 361690
rect 442264 361626 442316 361632
rect 439688 361616 439740 361622
rect 439688 361558 439740 361564
rect 438124 360256 438176 360262
rect 438124 360198 438176 360204
rect 438136 334286 438164 360198
rect 439596 336796 439648 336802
rect 439596 336738 439648 336744
rect 438216 336388 438268 336394
rect 438216 336330 438268 336336
rect 438124 334280 438176 334286
rect 438124 334222 438176 334228
rect 436928 329724 436980 329730
rect 436928 329666 436980 329672
rect 438228 318578 438256 336330
rect 439504 332716 439556 332722
rect 439504 332658 439556 332664
rect 438768 329792 438820 329798
rect 438768 329734 438820 329740
rect 438216 318572 438268 318578
rect 438216 318514 438268 318520
rect 436836 307760 436888 307766
rect 436836 307702 436888 307708
rect 436836 271312 436888 271318
rect 436836 271254 436888 271260
rect 436848 213042 436876 271254
rect 436836 213036 436888 213042
rect 436836 212978 436888 212984
rect 436744 183524 436796 183530
rect 436744 183466 436796 183472
rect 434904 162852 434956 162858
rect 434904 162794 434956 162800
rect 435364 162852 435416 162858
rect 435364 162794 435416 162800
rect 431868 161696 431920 161702
rect 431868 161638 431920 161644
rect 431316 160336 431368 160342
rect 431316 160278 431368 160284
rect 428016 159854 428688 159882
rect 431328 159882 431356 160278
rect 431880 159882 431908 161638
rect 434916 161634 434944 162794
rect 438780 161634 438808 329734
rect 439516 205630 439544 332658
rect 439608 271862 439636 336738
rect 439700 331362 439728 361558
rect 441068 360324 441120 360330
rect 441068 360266 441120 360272
rect 440976 336864 441028 336870
rect 440976 336806 441028 336812
rect 439780 335368 439832 335374
rect 439780 335310 439832 335316
rect 439688 331356 439740 331362
rect 439688 331298 439740 331304
rect 439792 325582 439820 335310
rect 440240 334280 440292 334286
rect 440240 334222 440292 334228
rect 440252 332586 440280 334222
rect 440240 332580 440292 332586
rect 440240 332522 440292 332528
rect 440884 331356 440936 331362
rect 440884 331298 440936 331304
rect 439780 325576 439832 325582
rect 439780 325518 439832 325524
rect 439688 286680 439740 286686
rect 439688 286622 439740 286628
rect 439596 271856 439648 271862
rect 439596 271798 439648 271804
rect 439700 271318 439728 286622
rect 439688 271312 439740 271318
rect 439688 271254 439740 271260
rect 440240 262812 440292 262818
rect 440240 262754 440292 262760
rect 440252 260370 440280 262754
rect 440240 260364 440292 260370
rect 440240 260306 440292 260312
rect 439596 244996 439648 245002
rect 439596 244938 439648 244944
rect 439608 230994 439636 244938
rect 439596 230988 439648 230994
rect 439596 230930 439648 230936
rect 439504 205624 439556 205630
rect 439504 205566 439556 205572
rect 440896 171834 440924 331298
rect 440988 260846 441016 336806
rect 441080 314566 441108 360266
rect 442276 344350 442304 361626
rect 442356 358896 442408 358902
rect 442356 358838 442408 358844
rect 442264 344344 442316 344350
rect 442264 344286 442316 344292
rect 441160 336252 441212 336258
rect 441160 336194 441212 336200
rect 441172 318510 441200 336194
rect 442264 335504 442316 335510
rect 442264 335446 442316 335452
rect 441620 326392 441672 326398
rect 441620 326334 441672 326340
rect 441160 318504 441212 318510
rect 441160 318446 441212 318452
rect 441068 314560 441120 314566
rect 441068 314502 441120 314508
rect 441632 305794 441660 326334
rect 441620 305788 441672 305794
rect 441620 305730 441672 305736
rect 440976 260840 441028 260846
rect 440976 260782 441028 260788
rect 442276 238746 442304 335446
rect 442368 330546 442396 358838
rect 442908 341012 442960 341018
rect 442908 340954 442960 340960
rect 442920 336054 442948 340954
rect 443736 339584 443788 339590
rect 443736 339526 443788 339532
rect 442908 336048 442960 336054
rect 442908 335990 442960 335996
rect 442540 335096 442592 335102
rect 442540 335038 442592 335044
rect 442446 334792 442502 334801
rect 442446 334727 442502 334736
rect 442356 330540 442408 330546
rect 442356 330482 442408 330488
rect 442460 319870 442488 334727
rect 442552 321638 442580 335038
rect 443644 334076 443696 334082
rect 443644 334018 443696 334024
rect 442632 332580 442684 332586
rect 442632 332522 442684 332528
rect 442644 322930 442672 332522
rect 442908 330132 442960 330138
rect 442908 330074 442960 330080
rect 442632 322924 442684 322930
rect 442632 322866 442684 322872
rect 442540 321632 442592 321638
rect 442540 321574 442592 321580
rect 442448 319864 442500 319870
rect 442448 319806 442500 319812
rect 442448 252476 442500 252482
rect 442448 252418 442500 252424
rect 442356 249756 442408 249762
rect 442356 249698 442408 249704
rect 442264 238740 442316 238746
rect 442264 238682 442316 238688
rect 442368 203590 442396 249698
rect 442460 245002 442488 252418
rect 442448 244996 442500 245002
rect 442448 244938 442500 244944
rect 442356 203584 442408 203590
rect 442356 203526 442408 203532
rect 440884 171828 440936 171834
rect 440884 171770 440936 171776
rect 434904 161628 434956 161634
rect 434904 161570 434956 161576
rect 438768 161628 438820 161634
rect 438768 161570 438820 161576
rect 434916 160206 434944 161570
rect 438780 161474 438808 161570
rect 442920 161566 442948 330074
rect 443000 269340 443052 269346
rect 443000 269282 443052 269288
rect 443012 262818 443040 269282
rect 443000 262812 443052 262818
rect 443000 262754 443052 262760
rect 443656 227730 443684 334018
rect 443748 304978 443776 339526
rect 443828 336320 443880 336326
rect 443828 336262 443880 336268
rect 443840 317422 443868 336262
rect 443920 335028 443972 335034
rect 443920 334970 443972 334976
rect 443932 319938 443960 334970
rect 444012 334960 444064 334966
rect 444012 334902 444064 334908
rect 444024 321842 444052 334902
rect 444116 329798 444144 445742
rect 444196 330608 444248 330614
rect 444196 330550 444248 330556
rect 444104 329792 444156 329798
rect 444104 329734 444156 329740
rect 444012 321836 444064 321842
rect 444012 321778 444064 321784
rect 443920 319932 443972 319938
rect 443920 319874 443972 319880
rect 443828 317416 443880 317422
rect 443828 317358 443880 317364
rect 443736 304972 443788 304978
rect 443736 304914 443788 304920
rect 443644 227724 443696 227730
rect 443644 227666 443696 227672
rect 442908 161560 442960 161566
rect 442908 161502 442960 161508
rect 438596 161446 438808 161474
rect 441620 161492 441672 161498
rect 434904 160200 434956 160206
rect 434904 160142 434956 160148
rect 435272 160200 435324 160206
rect 435272 160142 435324 160148
rect 431328 159854 431908 159882
rect 435284 159610 435312 160142
rect 438596 159882 438624 161446
rect 441620 161434 441672 161440
rect 441632 160154 441660 161434
rect 444208 161430 444236 330550
rect 444300 320142 444328 700402
rect 445036 321298 445064 700674
rect 445024 321292 445076 321298
rect 445024 321234 445076 321240
rect 445128 321230 445156 700742
rect 446496 700664 446548 700670
rect 446496 700606 446548 700612
rect 446404 700528 446456 700534
rect 446404 700470 446456 700476
rect 445208 700392 445260 700398
rect 445208 700334 445260 700340
rect 445668 700392 445720 700398
rect 445668 700334 445720 700340
rect 445116 321224 445168 321230
rect 445116 321166 445168 321172
rect 445220 321094 445248 700334
rect 445298 683360 445354 683369
rect 445298 683295 445354 683304
rect 445208 321088 445260 321094
rect 445208 321030 445260 321036
rect 444288 320136 444340 320142
rect 444288 320078 444340 320084
rect 445312 319394 445340 683295
rect 445392 683256 445444 683262
rect 445392 683198 445444 683204
rect 445404 320074 445432 683198
rect 445484 683188 445536 683194
rect 445484 683130 445536 683136
rect 445496 321201 445524 683130
rect 445576 444440 445628 444446
rect 445576 444382 445628 444388
rect 445588 386646 445616 444382
rect 445576 386640 445628 386646
rect 445576 386582 445628 386588
rect 445588 343126 445616 386582
rect 445576 343120 445628 343126
rect 445576 343062 445628 343068
rect 445588 342922 445616 343062
rect 445576 342916 445628 342922
rect 445576 342858 445628 342864
rect 445482 321192 445538 321201
rect 445482 321127 445538 321136
rect 445680 320958 445708 700334
rect 445852 444576 445904 444582
rect 445852 444518 445904 444524
rect 445760 444508 445812 444514
rect 445760 444450 445812 444456
rect 445772 330614 445800 444450
rect 445760 330608 445812 330614
rect 445760 330550 445812 330556
rect 445864 330138 445892 444518
rect 445852 330132 445904 330138
rect 445852 330074 445904 330080
rect 445668 320952 445720 320958
rect 445668 320894 445720 320900
rect 446416 320686 446444 700470
rect 446508 320822 446536 700606
rect 449164 700596 449216 700602
rect 449164 700538 449216 700544
rect 446680 685364 446732 685370
rect 446680 685306 446732 685312
rect 446588 685296 446640 685302
rect 446588 685238 446640 685244
rect 446496 320816 446548 320822
rect 446496 320758 446548 320764
rect 446404 320680 446456 320686
rect 446404 320622 446456 320628
rect 445392 320068 445444 320074
rect 445392 320010 445444 320016
rect 445300 319388 445352 319394
rect 445300 319330 445352 319336
rect 446600 319054 446628 685238
rect 446692 319598 446720 685306
rect 446864 683800 446916 683806
rect 446864 683742 446916 683748
rect 446770 683224 446826 683233
rect 446770 683159 446826 683168
rect 446784 319705 446812 683159
rect 446770 319696 446826 319705
rect 446770 319631 446826 319640
rect 446680 319592 446732 319598
rect 446680 319534 446732 319540
rect 446876 319258 446904 683742
rect 448336 526448 448388 526454
rect 448336 526390 448388 526396
rect 448244 522300 448296 522306
rect 448244 522242 448296 522248
rect 448060 519580 448112 519586
rect 448060 519522 448112 519528
rect 447968 518220 448020 518226
rect 447968 518162 448020 518168
rect 447322 516216 447378 516225
rect 447322 516151 447378 516160
rect 447336 499594 447364 516151
rect 447690 507240 447746 507249
rect 447690 507175 447746 507184
rect 447704 501650 447732 507175
rect 447874 503432 447930 503441
rect 447874 503367 447930 503376
rect 447888 501786 447916 503367
rect 447980 501945 448008 518162
rect 448072 505209 448100 519522
rect 448256 512825 448284 522242
rect 448348 514321 448376 526390
rect 448428 520940 448480 520946
rect 448428 520882 448480 520888
rect 448440 516338 448468 520882
rect 448440 516310 448560 516338
rect 448532 516225 448560 516310
rect 448518 516216 448574 516225
rect 448428 516180 448480 516186
rect 448518 516151 448574 516160
rect 448428 516122 448480 516128
rect 448334 514312 448390 514321
rect 448334 514247 448390 514256
rect 448242 512816 448298 512825
rect 448242 512751 448298 512760
rect 448150 510504 448206 510513
rect 448150 510439 448206 510448
rect 448058 505200 448114 505209
rect 448058 505135 448114 505144
rect 447966 501936 448022 501945
rect 447966 501871 448022 501880
rect 447888 501758 448008 501786
rect 447704 501622 447916 501650
rect 447324 499588 447376 499594
rect 447324 499530 447376 499536
rect 446956 447160 447008 447166
rect 446956 447102 447008 447108
rect 446968 349110 446996 447102
rect 447140 385008 447192 385014
rect 447140 384950 447192 384956
rect 447152 383897 447180 384950
rect 447138 383888 447194 383897
rect 447138 383823 447194 383832
rect 447140 383648 447192 383654
rect 447140 383590 447192 383596
rect 447152 383217 447180 383590
rect 447232 383580 447284 383586
rect 447232 383522 447284 383528
rect 447138 383208 447194 383217
rect 447138 383143 447194 383152
rect 447244 382537 447272 383522
rect 447230 382528 447286 382537
rect 447230 382463 447286 382472
rect 447140 382220 447192 382226
rect 447140 382162 447192 382168
rect 447152 381857 447180 382162
rect 447232 382152 447284 382158
rect 447232 382094 447284 382100
rect 447138 381848 447194 381857
rect 447138 381783 447194 381792
rect 447244 381177 447272 382094
rect 447230 381168 447286 381177
rect 447230 381103 447286 381112
rect 447140 380860 447192 380866
rect 447140 380802 447192 380808
rect 447152 380497 447180 380802
rect 447232 380792 447284 380798
rect 447232 380734 447284 380740
rect 447138 380488 447194 380497
rect 447138 380423 447194 380432
rect 447244 379817 447272 380734
rect 447230 379808 447286 379817
rect 447230 379743 447286 379752
rect 447232 379500 447284 379506
rect 447232 379442 447284 379448
rect 447140 379432 447192 379438
rect 447140 379374 447192 379380
rect 447152 379137 447180 379374
rect 447138 379128 447194 379137
rect 447138 379063 447194 379072
rect 447244 378457 447272 379442
rect 447230 378448 447286 378457
rect 447230 378383 447286 378392
rect 447232 378140 447284 378146
rect 447232 378082 447284 378088
rect 447140 378072 447192 378078
rect 447140 378014 447192 378020
rect 447152 377777 447180 378014
rect 447138 377768 447194 377777
rect 447138 377703 447194 377712
rect 447244 377097 447272 378082
rect 447230 377088 447286 377097
rect 447230 377023 447286 377032
rect 447232 376712 447284 376718
rect 447232 376654 447284 376660
rect 447140 376644 447192 376650
rect 447140 376586 447192 376592
rect 447152 376417 447180 376586
rect 447138 376408 447194 376417
rect 447138 376343 447194 376352
rect 447244 375737 447272 376654
rect 447230 375728 447286 375737
rect 447230 375663 447286 375672
rect 447140 375352 447192 375358
rect 447140 375294 447192 375300
rect 447152 375057 447180 375294
rect 447232 375284 447284 375290
rect 447232 375226 447284 375232
rect 447138 375048 447194 375057
rect 447138 374983 447194 374992
rect 447244 374377 447272 375226
rect 447230 374368 447286 374377
rect 447230 374303 447286 374312
rect 447140 373992 447192 373998
rect 447140 373934 447192 373940
rect 447152 373697 447180 373934
rect 447232 373924 447284 373930
rect 447232 373866 447284 373872
rect 447138 373688 447194 373697
rect 447138 373623 447194 373632
rect 447244 373017 447272 373866
rect 447230 373008 447286 373017
rect 447230 372943 447286 372952
rect 447140 372564 447192 372570
rect 447140 372506 447192 372512
rect 447152 372337 447180 372506
rect 447232 372496 447284 372502
rect 447232 372438 447284 372444
rect 447138 372328 447194 372337
rect 447138 372263 447194 372272
rect 447244 371657 447272 372438
rect 447230 371648 447286 371657
rect 447230 371583 447286 371592
rect 447232 371204 447284 371210
rect 447232 371146 447284 371152
rect 447140 371136 447192 371142
rect 447140 371078 447192 371084
rect 447152 370977 447180 371078
rect 447138 370968 447194 370977
rect 447138 370903 447194 370912
rect 447244 370297 447272 371146
rect 447230 370288 447286 370297
rect 447230 370223 447286 370232
rect 447232 369844 447284 369850
rect 447232 369786 447284 369792
rect 447140 369776 447192 369782
rect 447140 369718 447192 369724
rect 447152 369617 447180 369718
rect 447138 369608 447194 369617
rect 447138 369543 447194 369552
rect 447244 368937 447272 369786
rect 447230 368928 447286 368937
rect 447230 368863 447286 368872
rect 447232 368484 447284 368490
rect 447232 368426 447284 368432
rect 447140 368416 447192 368422
rect 447140 368358 447192 368364
rect 447152 368257 447180 368358
rect 447138 368248 447194 368257
rect 447138 368183 447194 368192
rect 447244 367577 447272 368426
rect 447230 367568 447286 367577
rect 447230 367503 447286 367512
rect 447140 367056 447192 367062
rect 447140 366998 447192 367004
rect 447152 366217 447180 366998
rect 447232 366988 447284 366994
rect 447232 366930 447284 366936
rect 447244 366897 447272 366930
rect 447230 366888 447286 366897
rect 447230 366823 447286 366832
rect 447138 366208 447194 366217
rect 447138 366143 447194 366152
rect 447140 365696 447192 365702
rect 447140 365638 447192 365644
rect 447152 364857 447180 365638
rect 447232 365628 447284 365634
rect 447232 365570 447284 365576
rect 447244 365537 447272 365570
rect 447230 365528 447286 365537
rect 447230 365463 447286 365472
rect 447138 364848 447194 364857
rect 447138 364783 447194 364792
rect 447230 364168 447286 364177
rect 447230 364103 447286 364112
rect 447138 363488 447194 363497
rect 447138 363423 447194 363432
rect 447152 363050 447180 363423
rect 447140 363044 447192 363050
rect 447140 362986 447192 362992
rect 447244 362982 447272 364103
rect 447232 362976 447284 362982
rect 447232 362918 447284 362924
rect 447230 362808 447286 362817
rect 447230 362743 447286 362752
rect 447138 362128 447194 362137
rect 447138 362063 447194 362072
rect 447152 361622 447180 362063
rect 447244 361690 447272 362743
rect 447232 361684 447284 361690
rect 447232 361626 447284 361632
rect 447140 361616 447192 361622
rect 447140 361558 447192 361564
rect 447230 361448 447286 361457
rect 447230 361383 447286 361392
rect 447138 360768 447194 360777
rect 447138 360703 447194 360712
rect 447152 360330 447180 360703
rect 447140 360324 447192 360330
rect 447140 360266 447192 360272
rect 447244 360262 447272 361383
rect 447232 360256 447284 360262
rect 447232 360198 447284 360204
rect 447230 360088 447286 360097
rect 447230 360023 447286 360032
rect 447138 359408 447194 359417
rect 447138 359343 447194 359352
rect 447152 358834 447180 359343
rect 447244 358902 447272 360023
rect 447232 358896 447284 358902
rect 447232 358838 447284 358844
rect 447140 358828 447192 358834
rect 447140 358770 447192 358776
rect 447140 351960 447192 351966
rect 447138 351928 447140 351937
rect 447192 351928 447194 351937
rect 447138 351863 447194 351872
rect 447140 350600 447192 350606
rect 447138 350568 447140 350577
rect 447192 350568 447194 350577
rect 447138 350503 447194 350512
rect 446956 349104 447008 349110
rect 446956 349046 447008 349052
rect 447140 347744 447192 347750
rect 447140 347686 447192 347692
rect 447152 347177 447180 347686
rect 447138 347168 447194 347177
rect 447138 347103 447194 347112
rect 447336 345014 447364 499530
rect 447888 499526 447916 501622
rect 447876 499520 447928 499526
rect 447876 499462 447928 499468
rect 447692 387456 447744 387462
rect 447692 387398 447744 387404
rect 447704 353297 447732 387398
rect 447784 387252 447836 387258
rect 447784 387194 447836 387200
rect 447690 353288 447746 353297
rect 447690 353223 447746 353232
rect 447796 349217 447824 387194
rect 447782 349208 447838 349217
rect 447782 349143 447838 349152
rect 447784 349104 447836 349110
rect 447784 349046 447836 349052
rect 447336 344986 447456 345014
rect 447322 343768 447378 343777
rect 447322 343703 447378 343712
rect 447138 341728 447194 341737
rect 447138 341663 447194 341672
rect 447152 340950 447180 341663
rect 447230 341048 447286 341057
rect 447230 340983 447232 340992
rect 447284 340983 447286 340992
rect 447232 340954 447284 340960
rect 447140 340944 447192 340950
rect 447140 340886 447192 340892
rect 447138 340368 447194 340377
rect 447138 340303 447194 340312
rect 447152 339522 447180 340303
rect 447230 339688 447286 339697
rect 447230 339623 447286 339632
rect 447244 339590 447272 339623
rect 447232 339584 447284 339590
rect 447232 339526 447284 339532
rect 447140 339516 447192 339522
rect 447140 339458 447192 339464
rect 447230 339008 447286 339017
rect 447230 338943 447286 338952
rect 447138 338328 447194 338337
rect 447138 338263 447194 338272
rect 447152 338230 447180 338263
rect 447140 338224 447192 338230
rect 447140 338166 447192 338172
rect 447244 338162 447272 338943
rect 447232 338156 447284 338162
rect 447232 338098 447284 338104
rect 447230 337648 447286 337657
rect 447230 337583 447286 337592
rect 447138 336968 447194 336977
rect 447138 336903 447194 336912
rect 447152 336870 447180 336903
rect 447140 336864 447192 336870
rect 447140 336806 447192 336812
rect 447244 336802 447272 337583
rect 447232 336796 447284 336802
rect 447232 336738 447284 336744
rect 447336 336682 447364 343703
rect 447152 336654 447364 336682
rect 446956 336184 447008 336190
rect 446956 336126 447008 336132
rect 446864 319252 446916 319258
rect 446864 319194 446916 319200
rect 446588 319048 446640 319054
rect 446588 318990 446640 318996
rect 446968 317354 446996 336126
rect 447048 334892 447100 334898
rect 447048 334834 447100 334840
rect 447060 320754 447088 334834
rect 447048 320748 447100 320754
rect 447048 320690 447100 320696
rect 446956 317348 447008 317354
rect 446956 317290 447008 317296
rect 446588 288924 446640 288930
rect 446588 288866 446640 288872
rect 446600 286686 446628 288866
rect 446588 286680 446640 286686
rect 446588 286622 446640 286628
rect 446404 283620 446456 283626
rect 446404 283562 446456 283568
rect 445668 269816 445720 269822
rect 445668 269758 445720 269764
rect 445024 262812 445076 262818
rect 445024 262754 445076 262760
rect 445036 249762 445064 262754
rect 445024 249756 445076 249762
rect 445024 249698 445076 249704
rect 444932 162172 444984 162178
rect 444932 162114 444984 162120
rect 444944 161498 444972 162114
rect 445680 161498 445708 269758
rect 446416 269346 446444 283562
rect 446404 269340 446456 269346
rect 446404 269282 446456 269288
rect 447152 171134 447180 336654
rect 447230 336288 447286 336297
rect 447230 336223 447286 336232
rect 447244 335442 447272 336223
rect 447322 335608 447378 335617
rect 447322 335543 447378 335552
rect 447336 335510 447364 335543
rect 447324 335504 447376 335510
rect 447324 335446 447376 335452
rect 447232 335436 447284 335442
rect 447232 335378 447284 335384
rect 447322 334928 447378 334937
rect 447322 334863 447378 334872
rect 447230 334248 447286 334257
rect 447230 334183 447286 334192
rect 447244 334014 447272 334183
rect 447336 334082 447364 334863
rect 447324 334076 447376 334082
rect 447324 334018 447376 334024
rect 447232 334008 447284 334014
rect 447232 333950 447284 333956
rect 447322 333568 447378 333577
rect 447322 333503 447378 333512
rect 447230 332888 447286 332897
rect 447230 332823 447286 332832
rect 447244 332654 447272 332823
rect 447336 332722 447364 333503
rect 447324 332716 447376 332722
rect 447324 332658 447376 332664
rect 447232 332648 447284 332654
rect 447232 332590 447284 332596
rect 447230 331528 447286 331537
rect 447230 331463 447286 331472
rect 447244 331362 447272 331463
rect 447232 331356 447284 331362
rect 447232 331298 447284 331304
rect 447230 330848 447286 330857
rect 447230 330783 447286 330792
rect 447244 330614 447272 330783
rect 447232 330608 447284 330614
rect 447232 330550 447284 330556
rect 447230 330168 447286 330177
rect 447230 330103 447232 330112
rect 447284 330103 447286 330112
rect 447232 330074 447284 330080
rect 447232 329792 447284 329798
rect 447232 329734 447284 329740
rect 447244 329497 447272 329734
rect 447230 329488 447286 329497
rect 447230 329423 447286 329432
rect 447428 329338 447456 344986
rect 447796 344457 447824 349046
rect 447782 344448 447838 344457
rect 447782 344383 447838 344392
rect 447598 332208 447654 332217
rect 447598 332143 447654 332152
rect 447612 331294 447640 332143
rect 447600 331288 447652 331294
rect 447600 331230 447652 331236
rect 447244 329310 447456 329338
rect 447244 329118 447272 329310
rect 447232 329112 447284 329118
rect 447232 329054 447284 329060
rect 447244 328817 447272 329054
rect 447230 328808 447286 328817
rect 447230 328743 447286 328752
rect 447230 328128 447286 328137
rect 447230 328063 447286 328072
rect 447244 327758 447272 328063
rect 447232 327752 447284 327758
rect 447232 327694 447284 327700
rect 447888 327078 447916 499462
rect 447980 499458 448008 501758
rect 447968 499452 448020 499458
rect 447968 499394 448020 499400
rect 447232 327072 447284 327078
rect 447232 327014 447284 327020
rect 447876 327072 447928 327078
rect 447876 327014 447928 327020
rect 447244 326097 447272 327014
rect 447230 326088 447286 326097
rect 447230 326023 447286 326032
rect 447784 325644 447836 325650
rect 447784 325586 447836 325592
rect 447322 324048 447378 324057
rect 447322 323983 447378 323992
rect 447336 323610 447364 323983
rect 447324 323604 447376 323610
rect 447324 323546 447376 323552
rect 447796 315586 447824 325586
rect 447980 325582 448008 499394
rect 448072 325650 448100 505135
rect 448164 326777 448192 510439
rect 448256 498914 448284 512751
rect 448348 500290 448376 514247
rect 448440 510513 448468 516122
rect 448426 510504 448482 510513
rect 448426 510439 448482 510448
rect 448348 500274 448560 500290
rect 448348 500268 448572 500274
rect 448348 500262 448520 500268
rect 448244 498908 448296 498914
rect 448244 498850 448296 498856
rect 448256 334150 448284 498850
rect 448244 334144 448296 334150
rect 448244 334086 448296 334092
rect 448256 327457 448284 334086
rect 448348 328137 448376 500262
rect 448520 500210 448572 500216
rect 448980 387184 449032 387190
rect 448980 387126 449032 387132
rect 448428 386028 448480 386034
rect 448428 385970 448480 385976
rect 448440 357377 448468 385970
rect 448992 358057 449020 387126
rect 449072 387116 449124 387122
rect 449072 387058 449124 387064
rect 448978 358048 449034 358057
rect 448978 357983 449034 357992
rect 448426 357368 448482 357377
rect 448426 357303 448482 357312
rect 448426 351248 448482 351257
rect 448426 351183 448482 351192
rect 448334 328128 448390 328137
rect 448334 328063 448390 328072
rect 448242 327448 448298 327457
rect 448242 327383 448298 327392
rect 448150 326768 448206 326777
rect 448150 326703 448206 326712
rect 448164 326398 448192 326703
rect 448152 326392 448204 326398
rect 448152 326334 448204 326340
rect 448060 325644 448112 325650
rect 448060 325586 448112 325592
rect 447968 325576 448020 325582
rect 447968 325518 448020 325524
rect 447980 324737 448008 325518
rect 448072 325417 448100 325586
rect 448058 325408 448114 325417
rect 448058 325343 448114 325352
rect 447966 324728 448022 324737
rect 447966 324663 448022 324672
rect 448242 324728 448298 324737
rect 448242 324663 448298 324672
rect 447784 315580 447836 315586
rect 447784 315522 447836 315528
rect 447784 268592 447836 268598
rect 447784 268534 447836 268540
rect 447796 252482 447824 268534
rect 447784 252476 447836 252482
rect 447784 252418 447836 252424
rect 448256 232626 448284 324663
rect 448334 324048 448390 324057
rect 448334 323983 448390 323992
rect 448244 232620 448296 232626
rect 448244 232562 448296 232568
rect 448348 206310 448376 323983
rect 448336 206304 448388 206310
rect 448336 206246 448388 206252
rect 448440 196654 448468 351183
rect 449084 342417 449112 387058
rect 449070 342408 449126 342417
rect 449070 342343 449126 342352
rect 449072 336116 449124 336122
rect 449072 336058 449124 336064
rect 448980 334824 449032 334830
rect 448980 334766 449032 334772
rect 448992 321706 449020 334766
rect 448980 321700 449032 321706
rect 448980 321642 449032 321648
rect 449084 321026 449112 336058
rect 449176 321366 449204 700538
rect 449256 700324 449308 700330
rect 449256 700266 449308 700272
rect 449164 321360 449216 321366
rect 449164 321302 449216 321308
rect 449268 321162 449296 700266
rect 462332 670002 462360 703520
rect 478524 700398 478552 703520
rect 494808 700466 494836 703520
rect 494796 700460 494848 700466
rect 494796 700402 494848 700408
rect 478512 700392 478564 700398
rect 478512 700334 478564 700340
rect 527192 699825 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 527178 699816 527234 699825
rect 527178 699751 527234 699760
rect 450636 669996 450688 670002
rect 450636 669938 450688 669944
rect 462320 669996 462372 670002
rect 462320 669938 462372 669944
rect 449900 598324 449952 598330
rect 449900 598266 449952 598272
rect 449808 596828 449860 596834
rect 449808 596770 449860 596776
rect 449820 503441 449848 596770
rect 449806 503432 449862 503441
rect 449806 503367 449862 503376
rect 449716 499588 449768 499594
rect 449716 499530 449768 499536
rect 449728 498846 449756 499530
rect 449716 498840 449768 498846
rect 449716 498782 449768 498788
rect 449808 497548 449860 497554
rect 449808 497490 449860 497496
rect 449440 457496 449492 457502
rect 449440 457438 449492 457444
rect 449346 385656 449402 385665
rect 449346 385591 449402 385600
rect 449360 324057 449388 385591
rect 449452 356697 449480 457438
rect 449532 456068 449584 456074
rect 449532 456010 449584 456016
rect 449438 356688 449494 356697
rect 449438 356623 449494 356632
rect 449544 355337 449572 456010
rect 449716 454776 449768 454782
rect 449716 454718 449768 454724
rect 449624 454708 449676 454714
rect 449624 454650 449676 454656
rect 449530 355328 449586 355337
rect 449530 355263 449586 355272
rect 449636 354657 449664 454650
rect 449622 354648 449678 354657
rect 449622 354583 449678 354592
rect 449728 353977 449756 454718
rect 449820 356017 449848 497490
rect 449806 356008 449862 356017
rect 449806 355943 449862 355952
rect 449714 353968 449770 353977
rect 449714 353903 449770 353912
rect 449622 349888 449678 349897
rect 449622 349823 449678 349832
rect 449532 334756 449584 334762
rect 449532 334698 449584 334704
rect 449440 334688 449492 334694
rect 449440 334630 449492 334636
rect 449346 324048 449402 324057
rect 449346 323983 449402 323992
rect 449256 321156 449308 321162
rect 449256 321098 449308 321104
rect 449072 321020 449124 321026
rect 449072 320962 449124 320968
rect 449452 318442 449480 334630
rect 449544 320006 449572 334698
rect 449532 320000 449584 320006
rect 449532 319942 449584 319948
rect 449440 318436 449492 318442
rect 449440 318378 449492 318384
rect 449636 263566 449664 349823
rect 449912 346225 449940 598266
rect 450084 499860 450136 499866
rect 450084 499802 450136 499808
rect 449992 460964 450044 460970
rect 449992 460906 450044 460912
rect 450004 346905 450032 460906
rect 450096 389298 450124 499802
rect 450176 455524 450228 455530
rect 450176 455466 450228 455472
rect 450084 389292 450136 389298
rect 450084 389234 450136 389240
rect 450188 348945 450216 455466
rect 450268 454844 450320 454850
rect 450268 454786 450320 454792
rect 450280 353025 450308 454786
rect 450452 391332 450504 391338
rect 450452 391274 450504 391280
rect 450360 385144 450412 385150
rect 450360 385086 450412 385092
rect 450266 353016 450322 353025
rect 450266 352951 450322 352960
rect 450174 348936 450230 348945
rect 450174 348871 450230 348880
rect 450372 348265 450400 385086
rect 450464 358873 450492 391274
rect 450450 358864 450506 358873
rect 450450 358799 450506 358808
rect 450358 348256 450414 348265
rect 450358 348191 450414 348200
rect 449990 346896 450046 346905
rect 449990 346831 450046 346840
rect 449898 346216 449954 346225
rect 449898 346151 449954 346160
rect 449806 345128 449862 345137
rect 449806 345063 449862 345072
rect 449728 343126 449756 343157
rect 449716 343120 449768 343126
rect 449714 343088 449716 343097
rect 449768 343088 449770 343097
rect 449714 343023 449770 343032
rect 449624 263560 449676 263566
rect 449624 263502 449676 263508
rect 449728 249082 449756 343023
rect 449716 249076 449768 249082
rect 449716 249018 449768 249024
rect 448428 196648 448480 196654
rect 448428 196590 448480 196596
rect 447152 171106 447824 171134
rect 444932 161492 444984 161498
rect 444932 161434 444984 161440
rect 445668 161492 445720 161498
rect 445668 161434 445720 161440
rect 444196 161424 444248 161430
rect 444196 161366 444248 161372
rect 444208 160750 444236 161366
rect 444196 160744 444248 160750
rect 444196 160686 444248 160692
rect 444944 160154 444972 161434
rect 438288 159854 438624 159882
rect 441586 160126 441660 160154
rect 444898 160126 444972 160154
rect 441586 159868 441614 160126
rect 444898 159868 444926 160126
rect 447796 159882 447824 171106
rect 447796 159854 448224 159882
rect 421392 159582 421728 159610
rect 434976 159582 435312 159610
rect 420920 159520 420972 159526
rect 420920 159462 420972 159468
rect 449820 159390 449848 345063
rect 450542 334656 450598 334665
rect 450542 334591 450598 334600
rect 449990 331664 450046 331673
rect 449990 331599 450046 331608
rect 449900 322924 449952 322930
rect 449900 322866 449952 322872
rect 449912 320890 449940 322866
rect 449900 320884 449952 320890
rect 449900 320826 449952 320832
rect 449900 283688 449952 283694
rect 449900 283630 449952 283636
rect 449808 159384 449860 159390
rect 449808 159326 449860 159332
rect 449912 113174 449940 283630
rect 450004 195294 450032 331599
rect 450556 319190 450584 334591
rect 450544 319184 450596 319190
rect 450544 319126 450596 319132
rect 450648 319122 450676 669938
rect 459650 667992 459706 668001
rect 459650 667927 459706 667936
rect 458086 659968 458142 659977
rect 458086 659903 458142 659912
rect 457994 657520 458050 657529
rect 457994 657455 458050 657464
rect 457626 652896 457682 652905
rect 457626 652831 457682 652840
rect 457534 650176 457590 650185
rect 457534 650111 457590 650120
rect 457442 647728 457498 647737
rect 457442 647663 457498 647672
rect 457350 623928 457406 623937
rect 457350 623863 457406 623872
rect 457258 618352 457314 618361
rect 457258 618287 457314 618296
rect 457272 519654 457300 618287
rect 457364 596902 457392 623863
rect 457456 599622 457484 647663
rect 457548 599690 457576 650111
rect 457640 600302 457668 652831
rect 457902 643240 457958 643249
rect 457902 643175 457958 643184
rect 457718 621072 457774 621081
rect 457718 621007 457774 621016
rect 457628 600296 457680 600302
rect 457628 600238 457680 600244
rect 457536 599684 457588 599690
rect 457536 599626 457588 599632
rect 457444 599616 457496 599622
rect 457444 599558 457496 599564
rect 457352 596896 457404 596902
rect 457352 596838 457404 596844
rect 457732 543114 457760 621007
rect 457810 616040 457866 616049
rect 457810 615975 457866 615984
rect 457720 543108 457772 543114
rect 457720 543050 457772 543056
rect 457260 519648 457312 519654
rect 457260 519590 457312 519596
rect 457824 518430 457852 615975
rect 457916 598262 457944 643175
rect 457904 598256 457956 598262
rect 457904 598198 457956 598204
rect 457812 518424 457864 518430
rect 457812 518366 457864 518372
rect 458008 518022 458036 657455
rect 458100 520062 458128 659903
rect 459190 655752 459246 655761
rect 459190 655687 459246 655696
rect 459006 645960 459062 645969
rect 459006 645895 459062 645904
rect 458914 640384 458970 640393
rect 458914 640319 458970 640328
rect 458822 611416 458878 611425
rect 458822 611351 458878 611360
rect 458638 608696 458694 608705
rect 458638 608631 458694 608640
rect 458652 598398 458680 608631
rect 458732 603764 458784 603770
rect 458732 603706 458784 603712
rect 458640 598392 458692 598398
rect 458640 598334 458692 598340
rect 458744 598233 458772 603706
rect 458836 599758 458864 611351
rect 458824 599752 458876 599758
rect 458824 599694 458876 599700
rect 458928 599593 458956 640319
rect 459020 603770 459048 645895
rect 459098 628144 459154 628153
rect 459098 628079 459154 628088
rect 459008 603764 459060 603770
rect 459008 603706 459060 603712
rect 459006 603664 459062 603673
rect 459006 603599 459062 603608
rect 459020 599894 459048 603599
rect 459008 599888 459060 599894
rect 459008 599830 459060 599836
rect 458914 599584 458970 599593
rect 458914 599519 458970 599528
rect 458730 598224 458786 598233
rect 458730 598159 458786 598168
rect 458088 520056 458140 520062
rect 458088 519998 458140 520004
rect 459112 518294 459140 628079
rect 459204 543017 459232 655687
rect 459466 637936 459522 637945
rect 459466 637871 459522 637880
rect 459374 635488 459430 635497
rect 459374 635423 459430 635432
rect 459282 633448 459338 633457
rect 459282 633383 459338 633392
rect 459190 543008 459246 543017
rect 459190 542943 459246 542952
rect 459296 519625 459324 633383
rect 459282 519616 459338 519625
rect 459282 519551 459338 519560
rect 459388 519489 459416 635423
rect 459480 520985 459508 637871
rect 459558 626308 459614 626317
rect 459558 626243 459614 626252
rect 459466 520976 459522 520985
rect 459466 520911 459522 520920
rect 459374 519480 459430 519489
rect 459374 519415 459430 519424
rect 459572 518362 459600 626243
rect 459664 564398 459692 667927
rect 459834 614136 459890 614145
rect 459834 614071 459890 614080
rect 459742 601896 459798 601905
rect 459742 601831 459798 601840
rect 459652 564392 459704 564398
rect 459652 564334 459704 564340
rect 459756 518770 459784 601831
rect 459848 543046 459876 614071
rect 459926 606384 459982 606393
rect 459926 606319 459982 606328
rect 459940 598466 459968 606319
rect 461584 600296 461636 600302
rect 461584 600238 461636 600244
rect 459928 598460 459980 598466
rect 459928 598402 459980 598408
rect 459836 543040 459888 543046
rect 459836 542982 459888 542988
rect 459744 518764 459796 518770
rect 459744 518706 459796 518712
rect 459560 518356 459612 518362
rect 459560 518298 459612 518304
rect 459100 518288 459152 518294
rect 459100 518230 459152 518236
rect 457996 518016 458048 518022
rect 457996 517958 458048 517964
rect 450740 499866 450768 500140
rect 451292 500126 452226 500154
rect 450728 499860 450780 499866
rect 450728 499802 450780 499808
rect 450728 389292 450780 389298
rect 450728 389234 450780 389240
rect 450740 385914 450768 389234
rect 451292 385914 451320 500126
rect 452016 497616 452068 497622
rect 452016 497558 452068 497564
rect 451924 497480 451976 497486
rect 451924 497422 451976 497428
rect 451372 496868 451424 496874
rect 451372 496810 451424 496816
rect 451384 402974 451412 496810
rect 451384 402946 451872 402974
rect 451844 385914 451872 402946
rect 451936 386034 451964 497422
rect 452028 387462 452056 497558
rect 452844 496936 452896 496942
rect 452844 496878 452896 496884
rect 452016 387456 452068 387462
rect 452016 387398 452068 387404
rect 451924 386028 451976 386034
rect 451924 385970 451976 385976
rect 452856 385914 452884 496878
rect 453684 496874 453712 500140
rect 454040 497140 454092 497146
rect 454040 497082 454092 497088
rect 453672 496868 453724 496874
rect 453672 496810 453724 496816
rect 454052 389298 454080 497082
rect 454132 497072 454184 497078
rect 454132 497014 454184 497020
rect 454040 389292 454092 389298
rect 454040 389234 454092 389240
rect 453764 389156 453816 389162
rect 453764 389098 453816 389104
rect 450740 385886 450846 385914
rect 451292 385886 451582 385914
rect 451844 385886 452318 385914
rect 452856 385886 453054 385914
rect 453776 385900 453804 389098
rect 454144 385914 454172 497014
rect 455156 496942 455184 500140
rect 455420 497004 455472 497010
rect 455420 496946 455472 496952
rect 455144 496936 455196 496942
rect 455144 496878 455196 496884
rect 454684 496868 454736 496874
rect 454684 496810 454736 496816
rect 454696 389162 454724 496810
rect 455432 402974 455460 496946
rect 456628 496874 456656 500140
rect 458100 497078 458128 500140
rect 459572 497146 459600 500140
rect 459560 497140 459612 497146
rect 459560 497082 459612 497088
rect 458088 497072 458140 497078
rect 458088 497014 458140 497020
rect 461044 497010 461072 500140
rect 461032 497004 461084 497010
rect 461032 496946 461084 496952
rect 456616 496868 456668 496874
rect 456616 496810 456668 496816
rect 456892 429888 456944 429894
rect 456892 429830 456944 429836
rect 456904 402974 456932 429830
rect 457444 428460 457496 428466
rect 457444 428402 457496 428408
rect 455432 402946 455552 402974
rect 456904 402946 457024 402974
rect 454868 389292 454920 389298
rect 454868 389234 454920 389240
rect 454684 389156 454736 389162
rect 454684 389098 454736 389104
rect 454880 385914 454908 389234
rect 455524 385914 455552 402946
rect 456708 388476 456760 388482
rect 456708 388418 456760 388424
rect 454144 385886 454526 385914
rect 454880 385886 455262 385914
rect 455524 385886 455998 385914
rect 456720 385900 456748 388418
rect 456996 385914 457024 402946
rect 457456 388482 457484 428402
rect 461400 395344 461452 395350
rect 461400 395286 461452 395292
rect 458456 393984 458508 393990
rect 458456 393926 458508 393932
rect 458180 392692 458232 392698
rect 458180 392634 458232 392640
rect 457444 388476 457496 388482
rect 457444 388418 457496 388424
rect 456996 385886 457470 385914
rect 458192 385900 458220 392634
rect 458468 385914 458496 393926
rect 461124 392624 461176 392630
rect 461124 392566 461176 392572
rect 460388 391400 460440 391406
rect 460388 391342 460440 391348
rect 459652 387864 459704 387870
rect 459652 387806 459704 387812
rect 458468 385886 458942 385914
rect 459664 385900 459692 387806
rect 460400 385900 460428 391342
rect 461136 385900 461164 392566
rect 461412 385914 461440 395286
rect 461596 388550 461624 600238
rect 462424 600086 463266 600114
rect 462320 564392 462372 564398
rect 462320 564334 462372 564340
rect 461676 518016 461728 518022
rect 461676 517958 461728 517964
rect 461688 402974 461716 517958
rect 461688 402946 461808 402974
rect 461676 389904 461728 389910
rect 461676 389846 461728 389852
rect 461584 388544 461636 388550
rect 461584 388486 461636 388492
rect 461688 387870 461716 389846
rect 461780 388482 461808 402946
rect 461768 388476 461820 388482
rect 461768 388418 461820 388424
rect 461676 387864 461728 387870
rect 461676 387806 461728 387812
rect 462332 385914 462360 564334
rect 462424 518226 462452 600086
rect 463700 599888 463752 599894
rect 463700 599830 463752 599836
rect 462964 520464 463016 520470
rect 462964 520406 463016 520412
rect 462504 518764 462556 518770
rect 462504 518706 462556 518712
rect 462412 518220 462464 518226
rect 462412 518162 462464 518168
rect 462516 402974 462544 518706
rect 462516 402946 462912 402974
rect 462884 385914 462912 402946
rect 462976 387258 463004 520406
rect 463056 520056 463108 520062
rect 463056 519998 463108 520004
rect 463068 388618 463096 519998
rect 463056 388612 463108 388618
rect 463056 388554 463108 388560
rect 462964 387252 463016 387258
rect 462964 387194 463016 387200
rect 463712 385914 463740 599830
rect 465080 599752 465132 599758
rect 465080 599694 465132 599700
rect 463792 598460 463844 598466
rect 463792 598402 463844 598408
rect 463804 402974 463832 598402
rect 464344 543108 464396 543114
rect 464344 543050 464396 543056
rect 463804 402946 464292 402974
rect 464264 386050 464292 402946
rect 464356 388074 464384 543050
rect 465092 389298 465120 599694
rect 465172 598392 465224 598398
rect 465172 598334 465224 598340
rect 465080 389292 465132 389298
rect 465080 389234 465132 389240
rect 464344 388068 464396 388074
rect 464344 388010 464396 388016
rect 464264 386022 464384 386050
rect 464356 385914 464384 386022
rect 465184 385914 465212 598334
rect 468484 598256 468536 598262
rect 468484 598198 468536 598204
rect 465724 596896 465776 596902
rect 465724 596838 465776 596844
rect 465736 388006 465764 596838
rect 466460 543040 466512 543046
rect 466460 542982 466512 542988
rect 465908 389292 465960 389298
rect 465908 389234 465960 389240
rect 465724 388000 465776 388006
rect 465724 387942 465776 387948
rect 465920 385914 465948 389234
rect 466472 385914 466500 542982
rect 467102 522336 467158 522345
rect 467102 522271 467158 522280
rect 466552 518424 466604 518430
rect 466552 518366 466604 518372
rect 466564 402974 466592 518366
rect 466564 402946 466960 402974
rect 466932 386186 466960 402946
rect 467116 388686 467144 522271
rect 467932 519648 467984 519654
rect 467932 519590 467984 519596
rect 467944 402974 467972 519590
rect 467944 402946 468064 402974
rect 467104 388680 467156 388686
rect 467104 388622 467156 388628
rect 466932 386158 467328 386186
rect 467300 385914 467328 386158
rect 468036 385914 468064 402946
rect 468496 388890 468524 598198
rect 469600 596834 469628 600100
rect 469864 599684 469916 599690
rect 469864 599626 469916 599632
rect 469588 596828 469640 596834
rect 469588 596770 469640 596776
rect 468574 521112 468630 521121
rect 468574 521047 468630 521056
rect 468484 388884 468536 388890
rect 468484 388826 468536 388832
rect 468588 388822 468616 521047
rect 468576 388816 468628 388822
rect 468576 388758 468628 388764
rect 469876 388754 469904 599626
rect 469956 599616 470008 599622
rect 469956 599558 470008 599564
rect 469968 388958 469996 599558
rect 475948 598126 475976 600100
rect 482296 598262 482324 600100
rect 488644 598398 488672 600100
rect 488632 598392 488684 598398
rect 488632 598334 488684 598340
rect 494244 598392 494296 598398
rect 494244 598334 494296 598340
rect 482284 598256 482336 598262
rect 482284 598198 482336 598204
rect 494060 598256 494112 598262
rect 494060 598198 494112 598204
rect 493324 598188 493376 598194
rect 493324 598130 493376 598136
rect 473268 598120 473320 598126
rect 473268 598062 473320 598068
rect 475936 598120 475988 598126
rect 475936 598062 475988 598068
rect 473280 520402 473308 598062
rect 493336 522306 493364 598130
rect 493324 522300 493376 522306
rect 493324 522242 493376 522248
rect 488632 520464 488684 520470
rect 488632 520406 488684 520412
rect 472900 520396 472952 520402
rect 472900 520338 472952 520344
rect 473268 520396 473320 520402
rect 473268 520338 473320 520344
rect 472912 519586 472940 520338
rect 472900 519580 472952 519586
rect 472900 519522 472952 519528
rect 470692 518356 470744 518362
rect 470692 518298 470744 518304
rect 469956 388952 470008 388958
rect 469956 388894 470008 388900
rect 469864 388748 469916 388754
rect 469864 388690 469916 388696
rect 469220 388068 469272 388074
rect 469220 388010 469272 388016
rect 461412 385886 461886 385914
rect 462332 385886 462622 385914
rect 462884 385886 463358 385914
rect 463712 385886 464094 385914
rect 464356 385886 464830 385914
rect 465184 385886 465566 385914
rect 465920 385886 466302 385914
rect 466472 385886 467038 385914
rect 467300 385886 467774 385914
rect 468036 385886 468510 385914
rect 469232 385900 469260 388010
rect 469956 388000 470008 388006
rect 469956 387942 470008 387948
rect 469968 385900 469996 387942
rect 470704 385900 470732 518298
rect 470876 518288 470928 518294
rect 470876 518230 470928 518236
rect 470888 402974 470916 518230
rect 488644 517970 488672 520406
rect 488644 517942 488980 517970
rect 482664 517546 483000 517562
rect 480168 517540 480220 517546
rect 480168 517482 480220 517488
rect 482652 517540 483000 517546
rect 482704 517534 483000 517540
rect 482652 517482 482704 517488
rect 480180 461650 480208 517482
rect 491850 516216 491906 516225
rect 491850 516151 491852 516160
rect 491904 516151 491906 516160
rect 491852 516122 491904 516128
rect 494072 516066 494100 598198
rect 494256 586514 494284 598334
rect 494992 598194 495020 600100
rect 500972 600086 501354 600114
rect 506492 600086 507702 600114
rect 513392 600086 514050 600114
rect 494980 598188 495032 598194
rect 494980 598130 495032 598136
rect 493980 516038 494100 516066
rect 494164 586486 494284 586514
rect 493980 515250 494008 516038
rect 494058 515944 494114 515953
rect 494164 515930 494192 586486
rect 500972 526454 501000 600086
rect 500960 526448 501012 526454
rect 500960 526390 501012 526396
rect 506492 520946 506520 600086
rect 506480 520940 506532 520946
rect 506480 520882 506532 520888
rect 494244 520396 494296 520402
rect 494244 520338 494296 520344
rect 494114 515902 494192 515930
rect 494058 515879 494114 515888
rect 494072 515438 494100 515879
rect 494060 515432 494112 515438
rect 494060 515374 494112 515380
rect 493980 515222 494100 515250
rect 494072 513097 494100 515222
rect 494058 513088 494114 513097
rect 494058 513023 494114 513032
rect 494072 512038 494100 513023
rect 494060 512032 494112 512038
rect 494060 511974 494112 511980
rect 480272 500126 480608 500154
rect 481652 500126 481804 500154
rect 481928 500126 483000 500154
rect 483124 500126 484196 500154
rect 484412 500126 485392 500154
rect 486252 500126 486588 500154
rect 487172 500126 487784 500154
rect 488644 500126 488980 500154
rect 490176 500126 491156 500154
rect 480168 461644 480220 461650
rect 480168 461586 480220 461592
rect 480180 456822 480208 461586
rect 473728 456816 473780 456822
rect 473728 456758 473780 456764
rect 480168 456816 480220 456822
rect 480168 456758 480220 456764
rect 473740 455462 473768 456758
rect 473728 455456 473780 455462
rect 473728 455398 473780 455404
rect 473740 453900 473768 455398
rect 480272 454850 480300 500126
rect 481652 497622 481680 500126
rect 481640 497616 481692 497622
rect 481640 497558 481692 497564
rect 480996 455524 481048 455530
rect 480996 455466 481048 455472
rect 480260 454844 480312 454850
rect 480260 454786 480312 454792
rect 481008 453900 481036 455466
rect 481928 454782 481956 500126
rect 481916 454776 481968 454782
rect 481916 454718 481968 454724
rect 483124 454714 483152 500126
rect 484412 456074 484440 500126
rect 486252 497554 486280 500126
rect 486240 497548 486292 497554
rect 486240 497490 486292 497496
rect 487172 457502 487200 500126
rect 488644 497486 488672 500126
rect 488632 497480 488684 497486
rect 488632 497422 488684 497428
rect 487160 457496 487212 457502
rect 487160 457438 487212 457444
rect 484400 456068 484452 456074
rect 484400 456010 484452 456016
rect 488264 456068 488316 456074
rect 488264 456010 488316 456016
rect 483112 454708 483164 454714
rect 483112 454650 483164 454656
rect 487986 453928 488042 453937
rect 488276 453914 488304 456010
rect 488042 453900 488304 453914
rect 488042 453886 488290 453900
rect 487986 453863 488042 453872
rect 471624 428466 471652 432140
rect 474292 429894 474320 432140
rect 476132 432126 476974 432154
rect 474280 429888 474332 429894
rect 474280 429830 474332 429836
rect 471612 428460 471664 428466
rect 471612 428402 471664 428408
rect 470888 402946 471008 402974
rect 470980 385914 471008 402946
rect 476132 392698 476160 432126
rect 479628 429214 479656 432140
rect 481652 432126 482310 432154
rect 478144 429208 478196 429214
rect 478144 429150 478196 429156
rect 479616 429208 479668 429214
rect 479616 429150 479668 429156
rect 478156 393990 478184 429150
rect 478144 393984 478196 393990
rect 478144 393926 478196 393932
rect 476120 392692 476172 392698
rect 476120 392634 476172 392640
rect 472162 391232 472218 391241
rect 472162 391167 472218 391176
rect 470980 385886 471454 385914
rect 472176 385900 472204 391167
rect 481652 389910 481680 432126
rect 484964 429214 484992 432140
rect 487632 429214 487660 432140
rect 490024 432126 490314 432154
rect 482284 429208 482336 429214
rect 482284 429150 482336 429156
rect 484952 429208 485004 429214
rect 484952 429150 485004 429156
rect 486424 429208 486476 429214
rect 486424 429150 486476 429156
rect 487620 429208 487672 429214
rect 487620 429150 487672 429156
rect 482296 391406 482324 429150
rect 483020 423428 483072 423434
rect 483020 423370 483072 423376
rect 482284 391400 482336 391406
rect 482284 391342 482336 391348
rect 481640 389904 481692 389910
rect 481640 389846 481692 389852
rect 483032 389298 483060 423370
rect 485780 423360 485832 423366
rect 485780 423302 485832 423308
rect 483112 421592 483164 421598
rect 483112 421534 483164 421540
rect 483020 389292 483072 389298
rect 483020 389234 483072 389240
rect 472898 389056 472954 389065
rect 472898 388991 472954 389000
rect 474370 389056 474426 389065
rect 474370 388991 474426 389000
rect 475106 389056 475162 389065
rect 475106 388991 475162 389000
rect 476578 389056 476634 389065
rect 476578 388991 476634 389000
rect 479522 389056 479578 389065
rect 479522 388991 479578 389000
rect 472912 385900 472940 388991
rect 473634 388920 473690 388929
rect 473634 388855 473690 388864
rect 473648 385900 473676 388855
rect 474384 385900 474412 388991
rect 475120 385900 475148 388991
rect 475844 388884 475896 388890
rect 475844 388826 475896 388832
rect 475856 385900 475884 388826
rect 476592 385900 476620 388991
rect 477316 388952 477368 388958
rect 477316 388894 477368 388900
rect 477328 385900 477356 388894
rect 478052 388748 478104 388754
rect 478052 388690 478104 388696
rect 478064 385900 478092 388690
rect 478788 388544 478840 388550
rect 478788 388486 478840 388492
rect 478800 385900 478828 388486
rect 479536 385900 479564 388991
rect 481732 388816 481784 388822
rect 481732 388758 481784 388764
rect 480996 388612 481048 388618
rect 480996 388554 481048 388560
rect 480260 388476 480312 388482
rect 480260 388418 480312 388424
rect 480272 385900 480300 388418
rect 481008 385900 481036 388554
rect 481744 385900 481772 388758
rect 482468 388680 482520 388686
rect 482468 388622 482520 388628
rect 482480 385900 482508 388622
rect 483124 385914 483152 421534
rect 483572 389292 483624 389298
rect 483572 389234 483624 389240
rect 483584 385914 483612 389234
rect 484676 388952 484728 388958
rect 484676 388894 484728 388900
rect 483124 385886 483230 385914
rect 483584 385886 483966 385914
rect 484688 385900 484716 388894
rect 485412 388680 485464 388686
rect 485412 388622 485464 388628
rect 485424 385900 485452 388622
rect 485792 385914 485820 423302
rect 486436 392630 486464 429150
rect 487160 423292 487212 423298
rect 487160 423234 487212 423240
rect 486424 392624 486476 392630
rect 486424 392566 486476 392572
rect 486884 388612 486936 388618
rect 486884 388554 486936 388560
rect 485792 385886 486174 385914
rect 486896 385900 486924 388554
rect 487172 385914 487200 423234
rect 488540 423224 488592 423230
rect 488540 423166 488592 423172
rect 488552 402974 488580 423166
rect 488552 402946 488672 402974
rect 488356 388476 488408 388482
rect 488356 388418 488408 388424
rect 487172 385886 487646 385914
rect 488368 385900 488396 388418
rect 488644 385914 488672 402946
rect 490024 395350 490052 432126
rect 490012 395344 490064 395350
rect 490012 395286 490064 395292
rect 490564 392624 490616 392630
rect 490564 392566 490616 392572
rect 489828 388544 489880 388550
rect 489828 388486 489880 388492
rect 488644 385886 489118 385914
rect 489840 385900 489868 388486
rect 490576 385900 490604 392566
rect 491128 387190 491156 500126
rect 491312 500126 491372 500154
rect 491312 391338 491340 500126
rect 494072 499526 494100 511974
rect 494256 508881 494284 520338
rect 494242 508872 494298 508881
rect 494242 508807 494298 508816
rect 494256 508570 494284 508807
rect 494244 508564 494296 508570
rect 494244 508506 494296 508512
rect 494150 505200 494206 505209
rect 494150 505135 494206 505144
rect 494978 505200 495034 505209
rect 494978 505135 494980 505144
rect 494060 499520 494112 499526
rect 494060 499462 494112 499468
rect 494164 499458 494192 505135
rect 495032 505135 495034 505144
rect 494980 505106 495032 505112
rect 494702 501256 494758 501265
rect 494702 501191 494758 501200
rect 494152 499452 494204 499458
rect 494152 499394 494204 499400
rect 494716 462534 494744 501191
rect 511264 470620 511316 470626
rect 511264 470562 511316 470568
rect 494704 462528 494756 462534
rect 494704 462470 494756 462476
rect 494716 456074 494744 462470
rect 494704 456068 494756 456074
rect 494704 456010 494756 456016
rect 502984 423564 503036 423570
rect 502984 423506 503036 423512
rect 496820 423156 496872 423162
rect 496820 423098 496872 423104
rect 494060 420232 494112 420238
rect 494060 420174 494112 420180
rect 492680 398132 492732 398138
rect 492680 398074 492732 398080
rect 491576 395344 491628 395350
rect 491576 395286 491628 395292
rect 491392 393984 491444 393990
rect 491392 393926 491444 393932
rect 491300 391332 491352 391338
rect 491300 391274 491352 391280
rect 491404 389314 491432 393926
rect 491312 389286 491432 389314
rect 491116 387184 491168 387190
rect 491116 387126 491168 387132
rect 491312 385900 491340 389286
rect 491588 385914 491616 395286
rect 492692 389298 492720 398074
rect 492772 396772 492824 396778
rect 492772 396714 492824 396720
rect 492680 389292 492732 389298
rect 492680 389234 492732 389240
rect 491588 385886 492062 385914
rect 492784 385900 492812 396714
rect 494072 389298 494100 420174
rect 494152 399492 494204 399498
rect 494152 399434 494204 399440
rect 493140 389292 493192 389298
rect 493140 389234 493192 389240
rect 494060 389292 494112 389298
rect 494060 389234 494112 389240
rect 493152 385914 493180 389234
rect 494164 385914 494192 399434
rect 496452 391332 496504 391338
rect 496452 391274 496504 391280
rect 495716 389904 495768 389910
rect 495716 389846 495768 389852
rect 494612 389292 494664 389298
rect 494612 389234 494664 389240
rect 494624 385914 494652 389234
rect 493152 385886 493534 385914
rect 494164 385886 494270 385914
rect 494624 385886 495006 385914
rect 495728 385900 495756 389846
rect 496464 385900 496492 391274
rect 496832 385914 496860 423098
rect 498200 423088 498252 423094
rect 498200 423030 498252 423036
rect 497464 400920 497516 400926
rect 497464 400862 497516 400868
rect 497476 385914 497504 400862
rect 498212 385914 498240 423030
rect 499580 423020 499632 423026
rect 499580 422962 499632 422968
rect 499592 402974 499620 422962
rect 501052 422952 501104 422958
rect 501052 422894 501104 422900
rect 501064 402974 501092 422894
rect 499592 402946 499712 402974
rect 501064 402946 501184 402974
rect 499396 388816 499448 388822
rect 499396 388758 499448 388764
rect 496832 385886 497214 385914
rect 497476 385886 497950 385914
rect 498212 385886 498686 385914
rect 499408 385900 499436 388758
rect 499684 385914 499712 402946
rect 500868 388884 500920 388890
rect 500868 388826 500920 388832
rect 499684 385886 500158 385914
rect 500880 385900 500908 388826
rect 501156 385914 501184 402946
rect 502616 402280 502668 402286
rect 502616 402222 502668 402228
rect 502340 388748 502392 388754
rect 502340 388690 502392 388696
rect 501156 385886 501630 385914
rect 502352 385900 502380 388690
rect 502628 385914 502656 402222
rect 502996 388958 503024 423506
rect 507860 417784 507912 417790
rect 507860 417726 507912 417732
rect 503720 417716 503772 417722
rect 503720 417658 503772 417664
rect 502984 388952 503036 388958
rect 502984 388894 503036 388900
rect 503732 385914 503760 417658
rect 506480 417648 506532 417654
rect 506480 417590 506532 417596
rect 503996 417444 504048 417450
rect 503996 417386 504048 417392
rect 504008 402974 504036 417386
rect 504008 402946 504128 402974
rect 504100 385914 504128 402946
rect 506020 391264 506072 391270
rect 506020 391206 506072 391212
rect 505284 389836 505336 389842
rect 505284 389778 505336 389784
rect 502628 385886 503102 385914
rect 503732 385886 503838 385914
rect 504100 385886 504574 385914
rect 505296 385900 505324 389778
rect 506032 385900 506060 391206
rect 506492 389298 506520 417590
rect 506572 417580 506624 417586
rect 506572 417522 506624 417528
rect 506480 389292 506532 389298
rect 506480 389234 506532 389240
rect 506584 385914 506612 417522
rect 507872 389298 507900 417726
rect 507952 417512 508004 417518
rect 507952 417454 508004 417460
rect 507124 389292 507176 389298
rect 507124 389234 507176 389240
rect 507860 389292 507912 389298
rect 507860 389234 507912 389240
rect 507136 385914 507164 389234
rect 507964 385914 507992 417454
rect 508596 389292 508648 389298
rect 508596 389234 508648 389240
rect 508608 385914 508636 389234
rect 506584 385886 506782 385914
rect 507136 385886 507518 385914
rect 507964 385886 508254 385914
rect 508608 385886 508990 385914
rect 510710 364576 510766 364585
rect 510710 364511 510766 364520
rect 509790 362536 509846 362545
rect 509790 362471 509846 362480
rect 509330 360360 509386 360369
rect 509330 360295 509386 360304
rect 450728 334620 450780 334626
rect 450728 334562 450780 334568
rect 450740 321774 450768 334562
rect 509240 334008 509292 334014
rect 509240 333950 509292 333956
rect 509148 322244 509200 322250
rect 509148 322186 509200 322192
rect 454190 321858 454218 322116
rect 454190 321830 454264 321858
rect 450728 321768 450780 321774
rect 450728 321710 450780 321716
rect 450636 319116 450688 319122
rect 450636 319058 450688 319064
rect 453396 315512 453448 315518
rect 453396 315454 453448 315460
rect 450636 315444 450688 315450
rect 450636 315386 450688 315392
rect 450544 315376 450596 315382
rect 450544 315318 450596 315324
rect 450084 268456 450136 268462
rect 450084 268398 450136 268404
rect 450096 262818 450124 268398
rect 450084 262812 450136 262818
rect 450084 262754 450136 262760
rect 449992 195288 450044 195294
rect 449992 195230 450044 195236
rect 449912 113146 450492 113174
rect 445300 107364 445352 107370
rect 445300 107306 445352 107312
rect 439136 107296 439188 107302
rect 439136 107238 439188 107244
rect 432972 107228 433024 107234
rect 432972 107170 433024 107176
rect 426808 107160 426860 107166
rect 426808 107102 426860 107108
rect 420644 107092 420696 107098
rect 420644 107034 420696 107040
rect 414480 107024 414532 107030
rect 414480 106966 414532 106972
rect 410616 106276 410668 106282
rect 410616 106218 410668 106224
rect 410524 105596 410576 105602
rect 410524 105538 410576 105544
rect 414492 104938 414520 106966
rect 420656 104938 420684 107034
rect 426820 104938 426848 107102
rect 432984 104938 433012 107170
rect 439148 104938 439176 107238
rect 445312 104938 445340 107306
rect 450464 105346 450492 113146
rect 450556 107234 450584 315318
rect 450648 107302 450676 315386
rect 451924 314016 451976 314022
rect 451924 313958 451976 313964
rect 450728 271244 450780 271250
rect 450728 271186 450780 271192
rect 450636 107296 450688 107302
rect 450636 107238 450688 107244
rect 450544 107228 450596 107234
rect 450544 107170 450596 107176
rect 450740 107166 450768 271186
rect 450820 269952 450872 269958
rect 450820 269894 450872 269900
rect 450728 107160 450780 107166
rect 450728 107102 450780 107108
rect 450832 107098 450860 269894
rect 450912 160200 450964 160206
rect 450912 160142 450964 160148
rect 450924 142866 450952 160142
rect 450912 142860 450964 142866
rect 450912 142802 450964 142808
rect 451556 136536 451608 136542
rect 451554 136504 451556 136513
rect 451608 136504 451610 136513
rect 451554 136439 451610 136448
rect 451936 123593 451964 313958
rect 452108 311228 452160 311234
rect 452108 311170 452160 311176
rect 452016 286816 452068 286822
rect 452016 286758 452068 286764
rect 452028 124953 452056 286758
rect 452120 150385 452148 311170
rect 453304 309868 453356 309874
rect 453304 309810 453356 309816
rect 452292 283756 452344 283762
rect 452292 283698 452344 283704
rect 452200 268388 452252 268394
rect 452200 268330 452252 268336
rect 452106 150376 452162 150385
rect 452106 150311 452162 150320
rect 452212 126313 452240 268330
rect 452304 151745 452332 283698
rect 452384 278044 452436 278050
rect 452384 277986 452436 277992
rect 452396 171134 452424 277986
rect 452396 171106 452516 171134
rect 452384 157344 452436 157350
rect 452382 157312 452384 157321
rect 452436 157312 452438 157321
rect 452382 157247 452438 157256
rect 452384 155848 452436 155854
rect 452382 155816 452384 155825
rect 452436 155816 452438 155825
rect 452382 155751 452438 155760
rect 452384 154352 452436 154358
rect 452382 154320 452384 154329
rect 452436 154320 452438 154329
rect 452382 154255 452438 154264
rect 452488 153105 452516 171106
rect 452568 158432 452620 158438
rect 452566 158400 452568 158409
rect 452620 158400 452622 158409
rect 452566 158335 452622 158344
rect 452474 153096 452530 153105
rect 452474 153031 452530 153040
rect 452290 151736 452346 151745
rect 452290 151671 452346 151680
rect 452568 149048 452620 149054
rect 452566 149016 452568 149025
rect 452620 149016 452622 149025
rect 452566 148951 452622 148960
rect 452568 147552 452620 147558
rect 452566 147520 452568 147529
rect 452620 147520 452622 147529
rect 452566 147455 452622 147464
rect 452568 146192 452620 146198
rect 452566 146160 452568 146169
rect 452620 146160 452622 146169
rect 452566 146095 452622 146104
rect 452568 144832 452620 144838
rect 452566 144800 452568 144809
rect 452620 144800 452622 144809
rect 452566 144735 452622 144744
rect 452568 143472 452620 143478
rect 452566 143440 452568 143449
rect 452620 143440 452622 143449
rect 452566 143375 452622 143384
rect 452568 142112 452620 142118
rect 452566 142080 452568 142089
rect 452620 142080 452622 142089
rect 452566 142015 452622 142024
rect 452568 140752 452620 140758
rect 452566 140720 452568 140729
rect 452620 140720 452622 140729
rect 452566 140655 452622 140664
rect 452568 139392 452620 139398
rect 452566 139360 452568 139369
rect 452620 139360 452622 139369
rect 452566 139295 452622 139304
rect 452568 137896 452620 137902
rect 452566 137864 452568 137873
rect 452620 137864 452622 137873
rect 452566 137799 452622 137808
rect 452568 135176 452620 135182
rect 452566 135144 452568 135153
rect 452620 135144 452622 135153
rect 452566 135079 452622 135088
rect 452568 133816 452620 133822
rect 452566 133784 452568 133793
rect 452620 133784 452622 133793
rect 452566 133719 452622 133728
rect 452568 132456 452620 132462
rect 452566 132424 452568 132433
rect 452620 132424 452622 132433
rect 452566 132359 452622 132368
rect 452568 131096 452620 131102
rect 452566 131064 452568 131073
rect 452620 131064 452622 131073
rect 452566 130999 452622 131008
rect 452568 129736 452620 129742
rect 452566 129704 452568 129713
rect 452620 129704 452622 129713
rect 452566 129639 452622 129648
rect 452290 128344 452346 128353
rect 453316 128314 453344 309810
rect 453408 157350 453436 315454
rect 454236 305794 454264 321830
rect 454316 318980 454368 318986
rect 454316 318922 454368 318928
rect 454224 305788 454276 305794
rect 454224 305730 454276 305736
rect 454328 294438 454356 318922
rect 454420 296002 454448 322116
rect 454696 318986 454724 322116
rect 454684 318980 454736 318986
rect 454684 318922 454736 318928
rect 454776 316804 454828 316810
rect 454776 316746 454828 316752
rect 454684 316668 454736 316674
rect 454684 316610 454736 316616
rect 454408 295996 454460 296002
rect 454408 295938 454460 295944
rect 454316 294432 454368 294438
rect 454316 294374 454368 294380
rect 453580 285116 453632 285122
rect 453580 285058 453632 285064
rect 453488 275324 453540 275330
rect 453488 275266 453540 275272
rect 453396 157344 453448 157350
rect 453396 157286 453448 157292
rect 452290 128279 452292 128288
rect 452344 128279 452346 128288
rect 453304 128308 453356 128314
rect 452292 128250 452344 128256
rect 453304 128250 453356 128256
rect 452382 126984 452438 126993
rect 453500 126954 453528 275266
rect 453592 155854 453620 285058
rect 453672 273964 453724 273970
rect 453672 273906 453724 273912
rect 453580 155848 453632 155854
rect 453580 155790 453632 155796
rect 453684 154358 453712 273906
rect 453764 268524 453816 268530
rect 453764 268466 453816 268472
rect 453776 232558 453804 268466
rect 454040 232620 454092 232626
rect 454040 232562 454092 232568
rect 453764 232552 453816 232558
rect 453764 232494 453816 232500
rect 454052 221474 454080 232562
rect 454040 221468 454092 221474
rect 454040 221410 454092 221416
rect 453672 154352 453724 154358
rect 453672 154294 453724 154300
rect 452382 126919 452384 126928
rect 452436 126919 452438 126928
rect 453488 126948 453540 126954
rect 452384 126890 452436 126896
rect 453488 126890 453540 126896
rect 452198 126304 452254 126313
rect 452198 126239 452254 126248
rect 452014 124944 452070 124953
rect 452014 124879 452070 124888
rect 451922 123584 451978 123593
rect 451922 123519 451978 123528
rect 451924 122188 451976 122194
rect 451924 122130 451976 122136
rect 451936 121553 451964 122130
rect 451922 121544 451978 121553
rect 451922 121479 451978 121488
rect 450820 107092 450872 107098
rect 450820 107034 450872 107040
rect 454696 107030 454724 316610
rect 454684 107024 454736 107030
rect 454684 106966 454736 106972
rect 454788 106962 454816 316746
rect 454972 291718 455000 322116
rect 454960 291712 455012 291718
rect 454960 291654 455012 291660
rect 455248 290494 455276 322116
rect 455524 315314 455552 322116
rect 455512 315308 455564 315314
rect 455512 315250 455564 315256
rect 455800 304502 455828 322116
rect 456076 316742 456104 322116
rect 456352 321502 456380 322116
rect 456628 321570 456656 322116
rect 456616 321564 456668 321570
rect 456616 321506 456668 321512
rect 456340 321496 456392 321502
rect 456340 321438 456392 321444
rect 456904 318782 456932 322116
rect 457180 319326 457208 322116
rect 457168 319320 457220 319326
rect 457168 319262 457220 319268
rect 456892 318776 456944 318782
rect 456892 318718 456944 318724
rect 457456 318714 457484 322116
rect 457444 318708 457496 318714
rect 457444 318650 457496 318656
rect 457732 318646 457760 322116
rect 458008 321434 458036 322116
rect 458284 321473 458312 322116
rect 458270 321464 458326 321473
rect 457996 321428 458048 321434
rect 458270 321399 458326 321408
rect 457996 321370 458048 321376
rect 458560 320142 458588 322116
rect 458836 321230 458864 322116
rect 459112 321298 459140 322116
rect 459388 321366 459416 322116
rect 459376 321360 459428 321366
rect 459376 321302 459428 321308
rect 459100 321292 459152 321298
rect 459100 321234 459152 321240
rect 458824 321224 458876 321230
rect 458824 321166 458876 321172
rect 459664 320929 459692 322116
rect 459940 321065 459968 322116
rect 460216 321094 460244 322116
rect 460492 321162 460520 322116
rect 460768 321201 460796 322116
rect 460754 321192 460810 321201
rect 460480 321156 460532 321162
rect 460754 321127 460810 321136
rect 460480 321098 460532 321104
rect 460204 321088 460256 321094
rect 459926 321056 459982 321065
rect 460204 321030 460256 321036
rect 459926 320991 459982 321000
rect 459650 320920 459706 320929
rect 459650 320855 459706 320864
rect 458548 320136 458600 320142
rect 458548 320078 458600 320084
rect 461044 320074 461072 322116
rect 461320 320113 461348 322116
rect 461306 320104 461362 320113
rect 461032 320068 461084 320074
rect 461306 320039 461362 320048
rect 461032 320010 461084 320016
rect 461596 319938 461624 322116
rect 461872 320006 461900 322116
rect 462148 321842 462176 322116
rect 462136 321836 462188 321842
rect 462136 321778 462188 321784
rect 461860 320000 461912 320006
rect 461860 319942 461912 319948
rect 461584 319932 461636 319938
rect 461584 319874 461636 319880
rect 460204 319456 460256 319462
rect 460204 319398 460256 319404
rect 457720 318640 457772 318646
rect 457720 318582 457772 318588
rect 458824 318164 458876 318170
rect 458824 318106 458876 318112
rect 457444 318096 457496 318102
rect 457444 318038 457496 318044
rect 456064 316736 456116 316742
rect 456064 316678 456116 316684
rect 456892 315580 456944 315586
rect 456892 315522 456944 315528
rect 455788 304496 455840 304502
rect 455788 304438 455840 304444
rect 455236 290488 455288 290494
rect 455236 290430 455288 290436
rect 456800 286748 456852 286754
rect 456800 286690 456852 286696
rect 456248 282192 456300 282198
rect 456248 282134 456300 282140
rect 456156 274032 456208 274038
rect 456156 273974 456208 273980
rect 456064 272604 456116 272610
rect 456064 272546 456116 272552
rect 454960 272536 455012 272542
rect 454960 272478 455012 272484
rect 454868 271312 454920 271318
rect 454868 271254 454920 271260
rect 454880 107370 454908 271254
rect 454972 146198 455000 272478
rect 455052 270020 455104 270026
rect 455052 269962 455104 269968
rect 455064 158438 455092 269962
rect 455052 158432 455104 158438
rect 455052 158374 455104 158380
rect 454960 146192 455012 146198
rect 454960 146134 455012 146140
rect 456076 135182 456104 272546
rect 456168 137902 456196 273974
rect 456260 149054 456288 282134
rect 456340 271380 456392 271386
rect 456340 271322 456392 271328
rect 456248 149048 456300 149054
rect 456248 148990 456300 148996
rect 456352 142118 456380 271322
rect 456706 234968 456762 234977
rect 456706 234903 456762 234912
rect 456720 233918 456748 234903
rect 456708 233912 456760 233918
rect 456708 233854 456760 233860
rect 456706 207224 456762 207233
rect 456706 207159 456762 207168
rect 456720 206310 456748 207159
rect 456708 206304 456760 206310
rect 456708 206246 456760 206252
rect 456340 142112 456392 142118
rect 456340 142054 456392 142060
rect 456156 137896 456208 137902
rect 456156 137838 456208 137844
rect 456064 135176 456116 135182
rect 456064 135118 456116 135124
rect 456812 113174 456840 286690
rect 456904 234977 456932 315522
rect 456984 274712 457036 274718
rect 456984 274654 457036 274660
rect 456996 268598 457024 274654
rect 456984 268592 457036 268598
rect 456984 268534 457036 268540
rect 456984 263560 457036 263566
rect 456984 263502 457036 263508
rect 456996 262721 457024 263502
rect 456982 262712 457038 262721
rect 456982 262647 457038 262656
rect 456890 234968 456946 234977
rect 456890 234903 456946 234912
rect 457456 132462 457484 318038
rect 457628 314696 457680 314702
rect 457628 314638 457680 314644
rect 457536 305448 457588 305454
rect 457536 305390 457588 305396
rect 457548 136542 457576 305390
rect 457640 283626 457668 314638
rect 457628 283620 457680 283626
rect 457628 283562 457680 283568
rect 457720 276752 457772 276758
rect 457720 276694 457772 276700
rect 457628 275392 457680 275398
rect 457628 275334 457680 275340
rect 457640 140758 457668 275334
rect 457732 144838 457760 276694
rect 458088 249076 458140 249082
rect 458088 249018 458140 249024
rect 458100 248849 458128 249018
rect 458086 248840 458142 248849
rect 458086 248775 458142 248784
rect 457904 221468 457956 221474
rect 457904 221410 457956 221416
rect 457916 221105 457944 221410
rect 457902 221096 457958 221105
rect 457902 221031 457958 221040
rect 458100 200190 458128 248775
rect 458088 200184 458140 200190
rect 458088 200126 458140 200132
rect 457720 144832 457772 144838
rect 457720 144774 457772 144780
rect 457628 140752 457680 140758
rect 457628 140694 457680 140700
rect 457536 136536 457588 136542
rect 457536 136478 457588 136484
rect 457444 132456 457496 132462
rect 457444 132398 457496 132404
rect 458836 122194 458864 318106
rect 459008 316872 459060 316878
rect 459008 316814 459060 316820
rect 458916 308508 458968 308514
rect 458916 308450 458968 308456
rect 458928 129742 458956 308450
rect 459020 147558 459048 316814
rect 459100 293344 459152 293350
rect 459100 293286 459152 293292
rect 459008 147552 459060 147558
rect 459008 147494 459060 147500
rect 459112 131102 459140 293286
rect 459284 280832 459336 280838
rect 459284 280774 459336 280780
rect 459192 279472 459244 279478
rect 459192 279414 459244 279420
rect 459204 139398 459232 279414
rect 459296 143478 459324 280774
rect 459466 221096 459522 221105
rect 459466 221031 459522 221040
rect 459374 207224 459430 207233
rect 459374 207159 459430 207168
rect 459388 199442 459416 207159
rect 459480 200802 459508 221031
rect 459468 200796 459520 200802
rect 459468 200738 459520 200744
rect 459376 199436 459428 199442
rect 459376 199378 459428 199384
rect 459284 143472 459336 143478
rect 459284 143414 459336 143420
rect 459192 139392 459244 139398
rect 459192 139334 459244 139340
rect 459100 131096 459152 131102
rect 459100 131038 459152 131044
rect 458916 129736 458968 129742
rect 458916 129678 458968 129684
rect 458824 122188 458876 122194
rect 458824 122130 458876 122136
rect 456812 113146 456932 113174
rect 454868 107364 454920 107370
rect 454868 107306 454920 107312
rect 454776 106956 454828 106962
rect 454776 106898 454828 106904
rect 450464 105318 450768 105346
rect 407592 104910 408020 104938
rect 414184 104910 414520 104938
rect 420348 104910 420684 104938
rect 426512 104910 426848 104938
rect 432676 104910 433012 104938
rect 438840 104910 439176 104938
rect 445004 104910 445340 104938
rect 450740 104938 450768 105318
rect 456904 104938 456932 113146
rect 450740 104910 451168 104938
rect 456904 104910 457332 104938
rect 386328 62076 386380 62082
rect 386328 62018 386380 62024
rect 386236 33652 386288 33658
rect 386236 33594 386288 33600
rect 460216 31754 460244 319398
rect 461584 316736 461636 316742
rect 461584 316678 461636 316684
rect 461596 299470 461624 316678
rect 462424 314702 462452 322116
rect 462412 314696 462464 314702
rect 462412 314638 462464 314644
rect 461584 299464 461636 299470
rect 461584 299406 461636 299412
rect 462700 285734 462728 322116
rect 462976 302734 463004 322116
rect 463252 302802 463280 322116
rect 463528 306338 463556 322116
rect 463516 306332 463568 306338
rect 463516 306274 463568 306280
rect 463804 305522 463832 322116
rect 464080 305590 464108 322116
rect 464068 305584 464120 305590
rect 464068 305526 464120 305532
rect 463792 305516 463844 305522
rect 463792 305458 463844 305464
rect 463240 302796 463292 302802
rect 463240 302738 463292 302744
rect 462964 302728 463016 302734
rect 462964 302670 463016 302676
rect 464356 301578 464384 322116
rect 464632 308446 464660 322116
rect 464620 308440 464672 308446
rect 464620 308382 464672 308388
rect 464344 301572 464396 301578
rect 464344 301514 464396 301520
rect 464344 297220 464396 297226
rect 464344 297162 464396 297168
rect 464356 288930 464384 297162
rect 464344 288924 464396 288930
rect 464344 288866 464396 288872
rect 460388 285728 460440 285734
rect 460388 285670 460440 285676
rect 462688 285728 462740 285734
rect 462688 285670 462740 285676
rect 460296 276820 460348 276826
rect 460296 276762 460348 276768
rect 460308 133822 460336 276762
rect 460400 274718 460428 285670
rect 464908 285054 464936 322116
rect 465184 312594 465212 322116
rect 465172 312588 465224 312594
rect 465172 312530 465224 312536
rect 464896 285048 464948 285054
rect 464896 284990 464948 284996
rect 460388 274712 460440 274718
rect 460388 274654 460440 274660
rect 465460 269890 465488 322116
rect 465736 301578 465764 322116
rect 465724 301572 465776 301578
rect 465724 301514 465776 301520
rect 466012 287706 466040 322116
rect 466000 287700 466052 287706
rect 466000 287642 466052 287648
rect 466288 271182 466316 322116
rect 466564 313274 466592 322116
rect 466840 321366 466868 322116
rect 466828 321360 466880 321366
rect 466828 321302 466880 321308
rect 467116 320074 467144 322116
rect 467392 321094 467420 322116
rect 467668 321162 467696 322116
rect 467656 321156 467708 321162
rect 467656 321098 467708 321104
rect 467380 321088 467432 321094
rect 467380 321030 467432 321036
rect 467104 320068 467156 320074
rect 467104 320010 467156 320016
rect 467944 319734 467972 322116
rect 468220 321298 468248 322116
rect 468208 321292 468260 321298
rect 468208 321234 468260 321240
rect 467932 319728 467984 319734
rect 467932 319670 467984 319676
rect 468496 319666 468524 322116
rect 468772 319802 468800 322116
rect 469048 320958 469076 322116
rect 469036 320952 469088 320958
rect 469036 320894 469088 320900
rect 469220 320884 469272 320890
rect 469220 320826 469272 320832
rect 469232 320142 469260 320826
rect 469220 320136 469272 320142
rect 469220 320078 469272 320084
rect 468760 319796 468812 319802
rect 468760 319738 468812 319744
rect 469324 319682 469352 322116
rect 468484 319660 468536 319666
rect 468484 319602 468536 319608
rect 469140 319654 469352 319682
rect 469140 319530 469168 319654
rect 469600 319598 469628 322116
rect 469876 320686 469904 322116
rect 469864 320680 469916 320686
rect 469864 320622 469916 320628
rect 469588 319592 469640 319598
rect 469588 319534 469640 319540
rect 469128 319524 469180 319530
rect 469128 319466 469180 319472
rect 469220 319524 469272 319530
rect 469220 319466 469272 319472
rect 469232 317218 469260 319466
rect 470152 319054 470180 322116
rect 470140 319048 470192 319054
rect 470140 318990 470192 318996
rect 470428 318510 470456 322116
rect 470704 318578 470732 322116
rect 470980 319841 471008 322116
rect 470966 319832 471022 319841
rect 470966 319767 471022 319776
rect 471256 319705 471284 322116
rect 471242 319696 471298 319705
rect 471242 319631 471298 319640
rect 471532 319394 471560 322116
rect 471808 319870 471836 322116
rect 471796 319864 471848 319870
rect 471796 319806 471848 319812
rect 471520 319388 471572 319394
rect 471520 319330 471572 319336
rect 470692 318572 470744 318578
rect 470692 318514 470744 318520
rect 470416 318504 470468 318510
rect 470416 318446 470468 318452
rect 472084 318442 472112 322116
rect 472360 321706 472388 322116
rect 472348 321700 472400 321706
rect 472348 321642 472400 321648
rect 472636 320142 472664 322116
rect 472624 320136 472676 320142
rect 472624 320078 472676 320084
rect 472912 319530 472940 322116
rect 472900 319524 472952 319530
rect 472900 319466 472952 319472
rect 472072 318436 472124 318442
rect 472072 318378 472124 318384
rect 467104 317212 467156 317218
rect 467104 317154 467156 317160
rect 469220 317212 469272 317218
rect 469220 317154 469272 317160
rect 466552 313268 466604 313274
rect 466552 313210 466604 313216
rect 467116 297226 467144 317154
rect 472624 316940 472676 316946
rect 472624 316882 472676 316888
rect 467104 297220 467156 297226
rect 467104 297162 467156 297168
rect 471244 282260 471296 282266
rect 471244 282202 471296 282208
rect 466276 271176 466328 271182
rect 466276 271118 466328 271124
rect 465448 269884 465500 269890
rect 465448 269826 465500 269832
rect 471256 268462 471284 282202
rect 472636 268530 472664 316882
rect 473188 299946 473216 322116
rect 473464 317218 473492 322116
rect 473452 317212 473504 317218
rect 473452 317154 473504 317160
rect 473740 306134 473768 322116
rect 473912 317212 473964 317218
rect 473912 317154 473964 317160
rect 473728 306128 473780 306134
rect 473728 306070 473780 306076
rect 473924 302870 473952 317154
rect 474016 306202 474044 322116
rect 474292 306270 474320 322116
rect 474568 319462 474596 322116
rect 474556 319456 474608 319462
rect 474556 319398 474608 319404
rect 474280 306264 474332 306270
rect 474280 306206 474332 306212
rect 474004 306196 474056 306202
rect 474004 306138 474056 306144
rect 473912 302864 473964 302870
rect 473912 302806 473964 302812
rect 473176 299940 473228 299946
rect 473176 299882 473228 299888
rect 474004 288856 474056 288862
rect 474004 288798 474056 288804
rect 474016 282266 474044 288798
rect 474844 284986 474872 322116
rect 475120 309806 475148 322116
rect 475396 311166 475424 322116
rect 475384 311160 475436 311166
rect 475384 311102 475436 311108
rect 475108 309800 475160 309806
rect 475108 309742 475160 309748
rect 475672 286686 475700 322116
rect 475948 293282 475976 322116
rect 476224 297226 476252 322116
rect 476212 297220 476264 297226
rect 476212 297162 476264 297168
rect 475936 293276 475988 293282
rect 475936 293218 475988 293224
rect 475660 286680 475712 286686
rect 475660 286622 475712 286628
rect 474832 284980 474884 284986
rect 474832 284922 474884 284928
rect 476500 283626 476528 322116
rect 476488 283620 476540 283626
rect 476488 283562 476540 283568
rect 474004 282260 474056 282266
rect 474004 282202 474056 282208
rect 476776 273222 476804 322116
rect 477052 320142 477080 322116
rect 477040 320136 477092 320142
rect 477040 320078 477092 320084
rect 477328 319598 477356 322116
rect 477604 321230 477632 322116
rect 477592 321224 477644 321230
rect 477592 321166 477644 321172
rect 477880 320006 477908 322116
rect 477868 320000 477920 320006
rect 477868 319942 477920 319948
rect 477316 319592 477368 319598
rect 477316 319534 477368 319540
rect 478156 319394 478184 322116
rect 478432 319870 478460 322116
rect 478708 319938 478736 322116
rect 478696 319932 478748 319938
rect 478696 319874 478748 319880
rect 478420 319864 478472 319870
rect 478420 319806 478472 319812
rect 478984 319530 479012 322116
rect 479260 320113 479288 322116
rect 479246 320104 479302 320113
rect 479246 320039 479302 320048
rect 478972 319524 479024 319530
rect 478972 319466 479024 319472
rect 478144 319388 478196 319394
rect 478144 319330 478196 319336
rect 479536 319122 479564 322116
rect 479812 321026 479840 322116
rect 479800 321020 479852 321026
rect 479800 320962 479852 320968
rect 480088 320822 480116 322116
rect 480076 320816 480128 320822
rect 480076 320758 480128 320764
rect 480364 319258 480392 322116
rect 480640 319977 480668 322116
rect 480916 321337 480944 322116
rect 480902 321328 480958 321337
rect 480902 321263 480958 321272
rect 480626 319968 480682 319977
rect 480626 319903 480682 319912
rect 480812 319456 480864 319462
rect 480812 319398 480864 319404
rect 480352 319252 480404 319258
rect 480352 319194 480404 319200
rect 479524 319116 479576 319122
rect 479524 319058 479576 319064
rect 480260 317280 480312 317286
rect 480260 317222 480312 317228
rect 480272 312458 480300 317222
rect 480824 316946 480852 319398
rect 481192 317354 481220 322116
rect 481468 319569 481496 322116
rect 481454 319560 481510 319569
rect 481454 319495 481510 319504
rect 481744 317422 481772 322116
rect 482020 319190 482048 322116
rect 482296 321638 482324 322116
rect 482572 321774 482600 322116
rect 482560 321768 482612 321774
rect 482560 321710 482612 321716
rect 482284 321632 482336 321638
rect 482284 321574 482336 321580
rect 482848 320754 482876 322116
rect 482836 320748 482888 320754
rect 482836 320690 482888 320696
rect 483124 319462 483152 322116
rect 483112 319456 483164 319462
rect 483112 319398 483164 319404
rect 482008 319184 482060 319190
rect 482008 319126 482060 319132
rect 481732 317416 481784 317422
rect 481732 317358 481784 317364
rect 481180 317348 481232 317354
rect 481180 317290 481232 317296
rect 483400 317286 483428 322116
rect 483388 317280 483440 317286
rect 483388 317222 483440 317228
rect 480812 316940 480864 316946
rect 480812 316882 480864 316888
rect 478144 312452 478196 312458
rect 478144 312394 478196 312400
rect 480260 312452 480312 312458
rect 480260 312394 480312 312400
rect 478156 288862 478184 312394
rect 483676 300014 483704 322116
rect 483952 303618 483980 322116
rect 484228 305930 484256 322116
rect 484504 305998 484532 322116
rect 484780 306066 484808 322116
rect 484768 306060 484820 306066
rect 484768 306002 484820 306008
rect 484492 305992 484544 305998
rect 484492 305934 484544 305940
rect 484216 305924 484268 305930
rect 484216 305866 484268 305872
rect 483940 303612 483992 303618
rect 483940 303554 483992 303560
rect 483664 300008 483716 300014
rect 483664 299950 483716 299956
rect 485056 298858 485084 322116
rect 485332 305862 485360 322116
rect 485608 313954 485636 322116
rect 485596 313948 485648 313954
rect 485596 313890 485648 313896
rect 485320 305856 485372 305862
rect 485320 305798 485372 305804
rect 485884 303618 485912 322116
rect 485872 303612 485924 303618
rect 485872 303554 485924 303560
rect 485044 298852 485096 298858
rect 485044 298794 485096 298800
rect 478144 288856 478196 288862
rect 478144 288798 478196 288804
rect 486160 284986 486188 322116
rect 486436 301646 486464 322116
rect 486424 301640 486476 301646
rect 486424 301582 486476 301588
rect 486148 284980 486200 284986
rect 486148 284922 486200 284928
rect 476764 273216 476816 273222
rect 476764 273158 476816 273164
rect 486712 270026 486740 322116
rect 486988 318170 487016 322116
rect 486976 318164 487028 318170
rect 486976 318106 487028 318112
rect 487264 314022 487292 322116
rect 487252 314016 487304 314022
rect 487252 313958 487304 313964
rect 487540 286822 487568 322116
rect 487528 286816 487580 286822
rect 487528 286758 487580 286764
rect 486700 270020 486752 270026
rect 486700 269962 486752 269968
rect 472624 268524 472676 268530
rect 472624 268466 472676 268472
rect 471244 268456 471296 268462
rect 471244 268398 471296 268404
rect 487816 268394 487844 322116
rect 488092 275330 488120 322116
rect 488368 309874 488396 322116
rect 488356 309868 488408 309874
rect 488356 309810 488408 309816
rect 488644 308514 488672 322116
rect 488632 308508 488684 308514
rect 488632 308450 488684 308456
rect 488920 293350 488948 322116
rect 489196 318102 489224 322116
rect 489184 318096 489236 318102
rect 489184 318038 489236 318044
rect 488908 293344 488960 293350
rect 488908 293286 488960 293292
rect 489472 276826 489500 322116
rect 489460 276820 489512 276826
rect 489460 276762 489512 276768
rect 488080 275324 488132 275330
rect 488080 275266 488132 275272
rect 489748 272610 489776 322116
rect 490024 305454 490052 322116
rect 490300 316034 490328 322116
rect 490300 316006 490420 316034
rect 490012 305448 490064 305454
rect 490012 305390 490064 305396
rect 490392 274038 490420 316006
rect 490576 279478 490604 322116
rect 490564 279472 490616 279478
rect 490564 279414 490616 279420
rect 490852 275398 490880 322116
rect 490840 275392 490892 275398
rect 490840 275334 490892 275340
rect 490380 274032 490432 274038
rect 490380 273974 490432 273980
rect 489736 272604 489788 272610
rect 489736 272546 489788 272552
rect 491128 271386 491156 322116
rect 491404 280838 491432 322116
rect 491392 280832 491444 280838
rect 491392 280774 491444 280780
rect 491680 276758 491708 322116
rect 491668 276752 491720 276758
rect 491668 276694 491720 276700
rect 491956 272542 491984 322116
rect 492232 316878 492260 322116
rect 492220 316872 492272 316878
rect 492220 316814 492272 316820
rect 492508 282198 492536 322116
rect 492784 311234 492812 322116
rect 492772 311228 492824 311234
rect 492772 311170 492824 311176
rect 493060 283762 493088 322116
rect 493048 283756 493100 283762
rect 493048 283698 493100 283704
rect 492496 282192 492548 282198
rect 492496 282134 492548 282140
rect 493336 278050 493364 322116
rect 493324 278044 493376 278050
rect 493324 277986 493376 277992
rect 493612 273970 493640 322116
rect 493888 285122 493916 322116
rect 494164 315518 494192 322116
rect 494440 318102 494468 322116
rect 494428 318096 494480 318102
rect 494428 318038 494480 318044
rect 494152 315512 494204 315518
rect 494152 315454 494204 315460
rect 493876 285116 493928 285122
rect 493876 285058 493928 285064
rect 493600 273964 493652 273970
rect 493600 273906 493652 273912
rect 491944 272536 491996 272542
rect 491944 272478 491996 272484
rect 491116 271380 491168 271386
rect 491116 271322 491168 271328
rect 494716 268394 494744 322116
rect 494992 271386 495020 322116
rect 495268 275398 495296 322116
rect 495256 275392 495308 275398
rect 495256 275334 495308 275340
rect 495544 273970 495572 322116
rect 495820 275330 495848 322116
rect 496096 316878 496124 322116
rect 496084 316872 496136 316878
rect 496084 316814 496136 316820
rect 495808 275324 495860 275330
rect 495808 275266 495860 275272
rect 495532 273964 495584 273970
rect 495532 273906 495584 273912
rect 496372 272542 496400 322116
rect 496648 314022 496676 322116
rect 496636 314016 496688 314022
rect 496636 313958 496688 313964
rect 496924 276758 496952 322116
rect 497200 316946 497228 322116
rect 497188 316940 497240 316946
rect 497188 316882 497240 316888
rect 496912 276752 496964 276758
rect 496912 276694 496964 276700
rect 497476 274038 497504 322116
rect 497752 275466 497780 322116
rect 498028 276826 498056 322116
rect 498304 315518 498332 322116
rect 498292 315512 498344 315518
rect 498292 315454 498344 315460
rect 498016 276820 498068 276826
rect 498016 276762 498068 276768
rect 497740 275460 497792 275466
rect 497740 275402 497792 275408
rect 497464 274032 497516 274038
rect 497464 273974 497516 273980
rect 498580 272610 498608 322116
rect 498856 278050 498884 322116
rect 498844 278044 498896 278050
rect 498844 277986 498896 277992
rect 499132 274106 499160 322116
rect 499120 274100 499172 274106
rect 499120 274042 499172 274048
rect 498568 272604 498620 272610
rect 498568 272546 498620 272552
rect 496360 272536 496412 272542
rect 496360 272478 496412 272484
rect 494980 271380 495032 271386
rect 494980 271322 495032 271328
rect 499408 268462 499436 322116
rect 499684 317014 499712 322116
rect 499672 317008 499724 317014
rect 499672 316950 499724 316956
rect 499960 270026 499988 322116
rect 499948 270020 500000 270026
rect 499948 269962 500000 269968
rect 500236 268530 500264 322116
rect 500512 270094 500540 322116
rect 500788 313993 500816 322116
rect 501064 315586 501092 322116
rect 501052 315580 501104 315586
rect 501052 315522 501104 315528
rect 500774 313984 500830 313993
rect 500774 313919 500830 313928
rect 501340 271454 501368 322116
rect 501616 317082 501644 322116
rect 501604 317076 501656 317082
rect 501604 317018 501656 317024
rect 501892 283762 501920 322116
rect 502168 319462 502196 322116
rect 502156 319456 502208 319462
rect 502156 319398 502208 319404
rect 502444 316810 502472 322116
rect 502432 316804 502484 316810
rect 502432 316746 502484 316752
rect 502720 301510 502748 322116
rect 502996 316742 503024 322116
rect 502984 316736 503036 316742
rect 502984 316678 503036 316684
rect 502708 301504 502760 301510
rect 502708 301446 502760 301452
rect 501880 283756 501932 283762
rect 501880 283698 501932 283704
rect 501328 271448 501380 271454
rect 501328 271390 501380 271396
rect 500500 270088 500552 270094
rect 500500 270030 500552 270036
rect 503272 269958 503300 322116
rect 503548 271250 503576 322116
rect 503824 315382 503852 322116
rect 504100 315450 504128 322116
rect 504088 315444 504140 315450
rect 504088 315386 504140 315392
rect 503812 315376 503864 315382
rect 503812 315318 503864 315324
rect 504376 271318 504404 322116
rect 504652 283694 504680 322116
rect 504928 286754 504956 322116
rect 507216 321904 507268 321910
rect 507216 321846 507268 321852
rect 507766 321872 507822 321881
rect 507122 321736 507178 321745
rect 507122 321671 507178 321680
rect 506940 320884 506992 320890
rect 506940 320826 506992 320832
rect 506952 303414 506980 320826
rect 507032 320544 507084 320550
rect 507032 320486 507084 320492
rect 506940 303408 506992 303414
rect 506940 303350 506992 303356
rect 507044 300626 507072 320486
rect 507032 300620 507084 300626
rect 507032 300562 507084 300568
rect 504916 286748 504968 286754
rect 504916 286690 504968 286696
rect 507136 286618 507164 321671
rect 507228 288998 507256 321846
rect 507584 321836 507636 321842
rect 507766 321807 507822 321816
rect 507584 321778 507636 321784
rect 507400 320952 507452 320958
rect 507306 320920 507362 320929
rect 507400 320894 507452 320900
rect 507306 320855 507362 320864
rect 507320 289270 507348 320855
rect 507412 292534 507440 320894
rect 507490 320784 507546 320793
rect 507490 320719 507546 320728
rect 507400 292528 507452 292534
rect 507400 292470 507452 292476
rect 507308 289264 507360 289270
rect 507308 289206 507360 289212
rect 507504 289066 507532 320719
rect 507596 298110 507624 321778
rect 507674 321328 507730 321337
rect 507674 321263 507730 321272
rect 507584 298104 507636 298110
rect 507584 298046 507636 298052
rect 507688 291786 507716 321263
rect 507780 297362 507808 321807
rect 507952 321768 508004 321774
rect 507952 321710 508004 321716
rect 507860 321700 507912 321706
rect 507860 321642 507912 321648
rect 507872 319666 507900 321642
rect 507964 319734 507992 321710
rect 509160 320142 509188 322186
rect 509252 321910 509280 333950
rect 509240 321904 509292 321910
rect 509240 321846 509292 321852
rect 509148 320136 509200 320142
rect 509148 320078 509200 320084
rect 507952 319728 508004 319734
rect 507952 319670 508004 319676
rect 507860 319660 507912 319666
rect 507860 319602 507912 319608
rect 509344 300082 509372 360295
rect 509422 358864 509478 358873
rect 509422 358799 509478 358808
rect 509436 303210 509464 358799
rect 509514 357640 509570 357649
rect 509514 357575 509570 357584
rect 509528 303482 509556 357575
rect 509606 344040 509662 344049
rect 509606 343975 509662 343984
rect 509516 303476 509568 303482
rect 509516 303418 509568 303424
rect 509620 303249 509648 343975
rect 509698 334248 509754 334257
rect 509698 334183 509754 334192
rect 509712 334014 509740 334183
rect 509700 334008 509752 334014
rect 509700 333950 509752 333956
rect 509698 329352 509754 329361
rect 509698 329287 509754 329296
rect 509606 303240 509662 303249
rect 509424 303204 509476 303210
rect 509606 303175 509662 303184
rect 509424 303146 509476 303152
rect 509712 300257 509740 329287
rect 509698 300248 509754 300257
rect 509698 300183 509754 300192
rect 509332 300076 509384 300082
rect 509332 300018 509384 300024
rect 507768 297356 507820 297362
rect 507768 297298 507820 297304
rect 509804 294506 509832 362471
rect 509974 331528 510030 331537
rect 509974 331463 510030 331472
rect 509882 326632 509938 326641
rect 509882 326567 509938 326576
rect 509896 321842 509924 326567
rect 509884 321836 509936 321842
rect 509884 321778 509936 321784
rect 509988 320550 510016 331463
rect 510158 324320 510214 324329
rect 510158 324255 510214 324264
rect 510068 322380 510120 322386
rect 510068 322322 510120 322328
rect 510080 321774 510108 322322
rect 510068 321768 510120 321774
rect 510068 321710 510120 321716
rect 509976 320544 510028 320550
rect 509976 320486 510028 320492
rect 510172 306105 510200 324255
rect 510618 323232 510674 323241
rect 510618 323167 510674 323176
rect 510528 322448 510580 322454
rect 510528 322390 510580 322396
rect 510540 319394 510568 322390
rect 510528 319388 510580 319394
rect 510528 319330 510580 319336
rect 510158 306096 510214 306105
rect 510158 306031 510214 306040
rect 509792 294500 509844 294506
rect 509792 294442 509844 294448
rect 507676 291780 507728 291786
rect 507676 291722 507728 291728
rect 507492 289060 507544 289066
rect 507492 289002 507544 289008
rect 507216 288992 507268 288998
rect 507216 288934 507268 288940
rect 507124 286612 507176 286618
rect 507124 286554 507176 286560
rect 504640 283688 504692 283694
rect 504640 283630 504692 283636
rect 504364 271312 504416 271318
rect 504364 271254 504416 271260
rect 503536 271244 503588 271250
rect 503536 271186 503588 271192
rect 503260 269952 503312 269958
rect 503260 269894 503312 269900
rect 510632 269822 510660 323167
rect 510724 294574 510752 364511
rect 510986 362400 511042 362409
rect 510986 362335 511042 362344
rect 510894 356416 510950 356425
rect 510894 356351 510950 356360
rect 510908 295050 510936 356351
rect 511000 300830 511028 362335
rect 511078 352608 511134 352617
rect 511078 352543 511134 352552
rect 511092 303346 511120 352543
rect 511170 346080 511226 346089
rect 511170 346015 511226 346024
rect 511080 303340 511132 303346
rect 511080 303282 511132 303288
rect 511184 303113 511212 346015
rect 511276 321094 511304 470562
rect 513392 387122 513420 600086
rect 520384 598194 520412 600100
rect 526732 598330 526760 600100
rect 526720 598324 526772 598330
rect 526720 598266 526772 598272
rect 519544 598188 519596 598194
rect 519544 598130 519596 598136
rect 520372 598188 520424 598194
rect 520372 598130 520424 598136
rect 515404 524476 515456 524482
rect 515404 524418 515456 524424
rect 513380 387116 513432 387122
rect 513380 387058 513432 387064
rect 512276 386572 512328 386578
rect 512276 386514 512328 386520
rect 512184 386504 512236 386510
rect 512184 386446 512236 386452
rect 512092 386436 512144 386442
rect 512092 386378 512144 386384
rect 512000 385076 512052 385082
rect 512000 385018 512052 385024
rect 512012 383874 512040 385018
rect 511920 383846 512040 383874
rect 511920 383466 511948 383846
rect 512104 383738 512132 386378
rect 512012 383710 512132 383738
rect 512012 383586 512040 383710
rect 512000 383580 512052 383586
rect 512000 383522 512052 383528
rect 511920 383438 512040 383466
rect 512012 378185 512040 383438
rect 512090 380352 512146 380361
rect 512090 380287 512146 380296
rect 512104 379914 512132 380287
rect 512092 379908 512144 379914
rect 512092 379850 512144 379856
rect 512196 378842 512224 386446
rect 512104 378814 512224 378842
rect 511998 378176 512054 378185
rect 511998 378111 512054 378120
rect 512104 376553 512132 378814
rect 512182 378720 512238 378729
rect 512182 378655 512238 378664
rect 512196 378350 512224 378655
rect 512184 378344 512236 378350
rect 512184 378286 512236 378292
rect 512288 377641 512316 386514
rect 512734 384704 512790 384713
rect 512734 384639 512790 384648
rect 512748 383790 512776 384639
rect 513286 384160 513342 384169
rect 513286 384095 513342 384104
rect 512736 383784 512788 383790
rect 512736 383726 512788 383732
rect 513300 383722 513328 384095
rect 513288 383716 513340 383722
rect 513288 383658 513340 383664
rect 513010 383616 513066 383625
rect 512552 383580 512604 383586
rect 513010 383551 513066 383560
rect 512552 383522 512604 383528
rect 512458 382528 512514 382537
rect 512458 382463 512460 382472
rect 512512 382463 512514 382472
rect 512460 382434 512512 382440
rect 512366 381984 512422 381993
rect 512366 381919 512422 381928
rect 512274 377632 512330 377641
rect 512274 377567 512330 377576
rect 512090 376544 512146 376553
rect 512090 376479 512146 376488
rect 512380 376038 512408 381919
rect 512368 376032 512420 376038
rect 512368 375974 512420 375980
rect 512458 376000 512514 376009
rect 512458 375935 512514 375944
rect 512472 375562 512500 375935
rect 512460 375556 512512 375562
rect 512460 375498 512512 375504
rect 512564 374921 512592 383522
rect 512826 383072 512882 383081
rect 512826 383007 512828 383016
rect 512880 383007 512882 383016
rect 512828 382978 512880 382984
rect 513024 382430 513052 383551
rect 513012 382424 513064 382430
rect 513012 382366 513064 382372
rect 513286 381440 513342 381449
rect 513286 381375 513342 381384
rect 513300 380934 513328 381375
rect 513288 380928 513340 380934
rect 512826 380896 512882 380905
rect 513288 380870 513340 380876
rect 512826 380831 512882 380840
rect 512840 377466 512868 380831
rect 514116 379908 514168 379914
rect 514116 379850 514168 379856
rect 513286 379808 513342 379817
rect 513286 379743 513342 379752
rect 513300 379574 513328 379743
rect 513288 379568 513340 379574
rect 513288 379510 513340 379516
rect 513286 379264 513342 379273
rect 513286 379199 513342 379208
rect 513300 378282 513328 379199
rect 513288 378276 513340 378282
rect 513288 378218 513340 378224
rect 514024 378208 514076 378214
rect 514024 378150 514076 378156
rect 512828 377460 512880 377466
rect 512828 377402 512880 377408
rect 513286 377088 513342 377097
rect 513286 377023 513342 377032
rect 513300 376854 513328 377023
rect 513288 376848 513340 376854
rect 513288 376790 513340 376796
rect 512734 375456 512790 375465
rect 512734 375391 512736 375400
rect 512788 375391 512790 375400
rect 512736 375362 512788 375368
rect 512550 374912 512606 374921
rect 512550 374847 512606 374856
rect 513286 374368 513342 374377
rect 513286 374303 513342 374312
rect 513300 374066 513328 374303
rect 513288 374060 513340 374066
rect 513288 374002 513340 374008
rect 512642 373824 512698 373833
rect 512642 373759 512698 373768
rect 512656 373386 512684 373759
rect 512644 373380 512696 373386
rect 512644 373322 512696 373328
rect 512642 373280 512698 373289
rect 512642 373215 512698 373224
rect 512656 372638 512684 373215
rect 513286 372736 513342 372745
rect 513286 372671 513288 372680
rect 513340 372671 513342 372680
rect 513288 372642 513340 372648
rect 512644 372632 512696 372638
rect 512644 372574 512696 372580
rect 512090 372192 512146 372201
rect 512090 372127 512146 372136
rect 512104 371414 512132 372127
rect 512182 371648 512238 371657
rect 512182 371583 512238 371592
rect 512092 371408 512144 371414
rect 512092 371350 512144 371356
rect 512090 371104 512146 371113
rect 512090 371039 512146 371048
rect 512104 371006 512132 371039
rect 512092 371000 512144 371006
rect 512092 370942 512144 370948
rect 512090 370016 512146 370025
rect 512090 369951 512146 369960
rect 511998 367840 512054 367849
rect 511998 367775 512054 367784
rect 512012 367198 512040 367775
rect 512000 367192 512052 367198
rect 512000 367134 512052 367140
rect 511538 365664 511594 365673
rect 511538 365599 511594 365608
rect 511446 347712 511502 347721
rect 511446 347647 511502 347656
rect 511356 333260 511408 333266
rect 511356 333202 511408 333208
rect 511264 321088 511316 321094
rect 511264 321030 511316 321036
rect 511368 319530 511396 333202
rect 511356 319524 511408 319530
rect 511356 319466 511408 319472
rect 511460 303550 511488 347647
rect 511448 303544 511500 303550
rect 511448 303486 511500 303492
rect 511170 303104 511226 303113
rect 511170 303039 511226 303048
rect 510988 300824 511040 300830
rect 510988 300766 511040 300772
rect 511552 300762 511580 365599
rect 511998 364032 512054 364041
rect 511998 363967 512054 363976
rect 512012 363390 512040 363967
rect 512000 363384 512052 363390
rect 512000 363326 512052 363332
rect 511998 361312 512054 361321
rect 511998 361247 512000 361256
rect 512052 361247 512054 361256
rect 512000 361218 512052 361224
rect 511998 358592 512054 358601
rect 511998 358527 512054 358536
rect 511540 300756 511592 300762
rect 511540 300698 511592 300704
rect 510896 295044 510948 295050
rect 510896 294986 510948 294992
rect 510712 294568 510764 294574
rect 510712 294510 510764 294516
rect 512012 276690 512040 358527
rect 512104 297770 512132 369951
rect 512196 305726 512224 371583
rect 513286 370560 513342 370569
rect 513342 370518 513604 370546
rect 513286 370495 513342 370504
rect 512734 369472 512790 369481
rect 512734 369407 512790 369416
rect 512274 368928 512330 368937
rect 512274 368863 512276 368872
rect 512328 368863 512330 368872
rect 512276 368834 512328 368840
rect 512748 368558 512776 369407
rect 512736 368552 512788 368558
rect 512736 368494 512788 368500
rect 513286 368384 513342 368393
rect 513286 368319 513342 368328
rect 513300 367402 513328 368319
rect 513288 367396 513340 367402
rect 513288 367338 513340 367344
rect 513286 367296 513342 367305
rect 513342 367254 513420 367282
rect 513286 367231 513342 367240
rect 513010 366752 513066 366761
rect 513010 366687 513066 366696
rect 513024 365770 513052 366687
rect 513286 366208 513342 366217
rect 513286 366143 513342 366152
rect 513300 365906 513328 366143
rect 513288 365900 513340 365906
rect 513288 365842 513340 365848
rect 513012 365764 513064 365770
rect 513012 365706 513064 365712
rect 512366 365120 512422 365129
rect 512366 365055 512422 365064
rect 512380 364334 512408 365055
rect 513392 364334 513420 367254
rect 512380 364306 512592 364334
rect 513392 364306 513512 364334
rect 512458 361856 512514 361865
rect 512458 361791 512514 361800
rect 512274 355872 512330 355881
rect 512274 355807 512330 355816
rect 512288 355434 512316 355807
rect 512276 355428 512328 355434
rect 512276 355370 512328 355376
rect 512472 355178 512500 361791
rect 512288 355150 512500 355178
rect 512184 305720 512236 305726
rect 512184 305662 512236 305668
rect 512288 297974 512316 355150
rect 512564 354674 512592 364306
rect 513286 363488 513342 363497
rect 513286 363423 513342 363432
rect 513300 363322 513328 363423
rect 513288 363316 513340 363322
rect 513288 363258 513340 363264
rect 513288 360256 513340 360262
rect 513286 360224 513288 360233
rect 513340 360224 513342 360233
rect 513286 360159 513342 360168
rect 512642 359680 512698 359689
rect 512642 359615 512698 359624
rect 512656 358902 512684 359615
rect 512644 358896 512696 358902
rect 512644 358838 512696 358844
rect 513194 358048 513250 358057
rect 513194 357983 513250 357992
rect 513208 357746 513236 357983
rect 513196 357740 513248 357746
rect 513196 357682 513248 357688
rect 513286 356960 513342 356969
rect 513286 356895 513342 356904
rect 513300 356386 513328 356895
rect 513288 356380 513340 356386
rect 513288 356322 513340 356328
rect 513286 355328 513342 355337
rect 513286 355263 513342 355272
rect 513300 355026 513328 355263
rect 513288 355020 513340 355026
rect 513288 354962 513340 354968
rect 513286 354784 513342 354793
rect 513286 354719 513288 354728
rect 513340 354719 513342 354728
rect 513288 354690 513340 354696
rect 512380 354646 512592 354674
rect 512380 304298 512408 354646
rect 512458 354240 512514 354249
rect 512458 354175 512514 354184
rect 512472 353394 512500 354175
rect 512826 353696 512882 353705
rect 512826 353631 512882 353640
rect 512840 353530 512868 353631
rect 512828 353524 512880 353530
rect 512828 353466 512880 353472
rect 512460 353388 512512 353394
rect 512460 353330 512512 353336
rect 513010 353152 513066 353161
rect 513010 353087 513066 353096
rect 513024 352714 513052 353087
rect 513012 352708 513064 352714
rect 513012 352650 513064 352656
rect 512458 352064 512514 352073
rect 512458 351999 512460 352008
rect 512512 351999 512514 352008
rect 512460 351970 512512 351976
rect 513286 351520 513342 351529
rect 513286 351455 513342 351464
rect 512458 350976 512514 350985
rect 513300 350946 513328 351455
rect 512458 350911 512514 350920
rect 513288 350940 513340 350946
rect 512472 350810 512500 350911
rect 513288 350882 513340 350888
rect 512460 350804 512512 350810
rect 512460 350746 512512 350752
rect 512826 350432 512882 350441
rect 512826 350367 512882 350376
rect 512458 349888 512514 349897
rect 512840 349858 512868 350367
rect 512458 349823 512514 349832
rect 512828 349852 512880 349858
rect 512472 349314 512500 349823
rect 512828 349794 512880 349800
rect 512550 349344 512606 349353
rect 512460 349308 512512 349314
rect 512550 349279 512606 349288
rect 512460 349250 512512 349256
rect 512564 349246 512592 349279
rect 512552 349240 512604 349246
rect 512552 349182 512604 349188
rect 513286 348800 513342 348809
rect 513286 348735 513342 348744
rect 513102 348256 513158 348265
rect 513102 348191 513158 348200
rect 513116 347818 513144 348191
rect 513300 347954 513328 348735
rect 513288 347948 513340 347954
rect 513288 347890 513340 347896
rect 513104 347812 513156 347818
rect 513104 347754 513156 347760
rect 513194 347168 513250 347177
rect 513194 347103 513250 347112
rect 512550 346624 512606 346633
rect 512550 346559 512606 346568
rect 512458 343360 512514 343369
rect 512458 343295 512514 343304
rect 512472 342582 512500 343295
rect 512460 342576 512512 342582
rect 512460 342518 512512 342524
rect 512458 334656 512514 334665
rect 512458 334591 512514 334600
rect 512472 334558 512500 334591
rect 512460 334552 512512 334558
rect 512460 334494 512512 334500
rect 512564 305658 512592 346559
rect 513102 341184 513158 341193
rect 513102 341119 513104 341128
rect 513156 341119 513158 341128
rect 513104 341090 513156 341096
rect 512642 340640 512698 340649
rect 512642 340575 512698 340584
rect 512552 305652 512604 305658
rect 512552 305594 512604 305600
rect 512368 304292 512420 304298
rect 512368 304234 512420 304240
rect 512656 302841 512684 340575
rect 513010 339008 513066 339017
rect 513010 338943 513066 338952
rect 513024 338162 513052 338943
rect 513012 338156 513064 338162
rect 513012 338098 513064 338104
rect 513010 337920 513066 337929
rect 513010 337855 513066 337864
rect 513024 337210 513052 337855
rect 513102 337376 513158 337385
rect 513102 337311 513158 337320
rect 513012 337204 513064 337210
rect 513012 337146 513064 337152
rect 513116 336802 513144 337311
rect 513104 336796 513156 336802
rect 513104 336738 513156 336744
rect 512826 335200 512882 335209
rect 512826 335135 512882 335144
rect 512840 334218 512868 335135
rect 512828 334212 512880 334218
rect 512828 334154 512880 334160
rect 512826 332480 512882 332489
rect 512826 332415 512882 332424
rect 512840 331498 512868 332415
rect 512828 331492 512880 331498
rect 512828 331434 512880 331440
rect 512734 328672 512790 328681
rect 512734 328607 512790 328616
rect 512748 305697 512776 328607
rect 512826 325408 512882 325417
rect 512826 325343 512882 325352
rect 512734 305688 512790 305697
rect 512734 305623 512790 305632
rect 512840 304366 512868 325343
rect 512918 323232 512974 323241
rect 512918 323167 512974 323176
rect 512932 322998 512960 323167
rect 512920 322992 512972 322998
rect 512920 322934 512972 322940
rect 512828 304360 512880 304366
rect 512828 304302 512880 304308
rect 512642 302832 512698 302841
rect 512642 302767 512698 302776
rect 513208 298790 513236 347103
rect 513286 345536 513342 345545
rect 513286 345471 513342 345480
rect 513300 345234 513328 345471
rect 513288 345228 513340 345234
rect 513288 345170 513340 345176
rect 513286 344992 513342 345001
rect 513286 344927 513342 344936
rect 513300 344282 513328 344927
rect 513288 344276 513340 344282
rect 513288 344218 513340 344224
rect 513286 343904 513342 343913
rect 513286 343839 513288 343848
rect 513340 343839 513342 343848
rect 513288 343810 513340 343816
rect 513288 342304 513340 342310
rect 513286 342272 513288 342281
rect 513340 342272 513342 342281
rect 513286 342207 513342 342216
rect 513286 341728 513342 341737
rect 513286 341663 513342 341672
rect 513300 341290 513328 341663
rect 513288 341284 513340 341290
rect 513288 341226 513340 341232
rect 513286 340096 513342 340105
rect 513286 340031 513342 340040
rect 513300 339658 513328 340031
rect 513288 339652 513340 339658
rect 513288 339594 513340 339600
rect 513286 339552 513342 339561
rect 513286 339487 513288 339496
rect 513340 339487 513342 339496
rect 513288 339458 513340 339464
rect 513286 338464 513342 338473
rect 513286 338399 513342 338408
rect 513300 338298 513328 338399
rect 513288 338292 513340 338298
rect 513288 338234 513340 338240
rect 513288 336932 513340 336938
rect 513288 336874 513340 336880
rect 513300 336841 513328 336874
rect 513286 336832 513342 336841
rect 513286 336767 513342 336776
rect 513286 336288 513342 336297
rect 513286 336223 513342 336232
rect 513300 336122 513328 336223
rect 513288 336116 513340 336122
rect 513288 336058 513340 336064
rect 513286 335744 513342 335753
rect 513286 335679 513342 335688
rect 513300 335374 513328 335679
rect 513288 335368 513340 335374
rect 513288 335310 513340 335316
rect 513286 333568 513342 333577
rect 513286 333503 513342 333512
rect 513300 332722 513328 333503
rect 513288 332716 513340 332722
rect 513288 332658 513340 332664
rect 513286 331936 513342 331945
rect 513342 331894 513420 331922
rect 513286 331871 513342 331880
rect 513392 320958 513420 331894
rect 513380 320952 513432 320958
rect 513380 320894 513432 320900
rect 513484 300558 513512 364306
rect 513576 302938 513604 370518
rect 513748 363384 513800 363390
rect 513748 363326 513800 363332
rect 513656 361276 513708 361282
rect 513656 361218 513708 361224
rect 513564 302932 513616 302938
rect 513564 302874 513616 302880
rect 513472 300552 513524 300558
rect 513472 300494 513524 300500
rect 513196 298784 513248 298790
rect 513196 298726 513248 298732
rect 512276 297968 512328 297974
rect 512276 297910 512328 297916
rect 512092 297764 512144 297770
rect 512092 297706 512144 297712
rect 513668 295118 513696 361218
rect 513760 300694 513788 363326
rect 513932 350804 513984 350810
rect 513932 350746 513984 350752
rect 513840 349308 513892 349314
rect 513840 349250 513892 349256
rect 513748 300688 513800 300694
rect 513748 300630 513800 300636
rect 513852 297566 513880 349250
rect 513944 303142 513972 350746
rect 514036 322522 514064 378150
rect 514128 358834 514156 379850
rect 514852 371408 514904 371414
rect 514852 371350 514904 371356
rect 514760 371000 514812 371006
rect 514760 370942 514812 370948
rect 514208 367192 514260 367198
rect 514208 367134 514260 367140
rect 514116 358828 514168 358834
rect 514116 358770 514168 358776
rect 514116 334552 514168 334558
rect 514116 334494 514168 334500
rect 514024 322516 514076 322522
rect 514024 322458 514076 322464
rect 514024 322312 514076 322318
rect 514024 322254 514076 322260
rect 514036 321706 514064 322254
rect 514024 321700 514076 321706
rect 514024 321642 514076 321648
rect 513932 303136 513984 303142
rect 513932 303078 513984 303084
rect 514128 298042 514156 334494
rect 514116 298036 514168 298042
rect 514116 297978 514168 297984
rect 513840 297560 513892 297566
rect 513840 297502 513892 297508
rect 514220 295254 514248 367134
rect 514300 322516 514352 322522
rect 514300 322458 514352 322464
rect 514312 319598 514340 322458
rect 514300 319592 514352 319598
rect 514300 319534 514352 319540
rect 514772 295322 514800 370942
rect 514864 300422 514892 371350
rect 514944 368892 514996 368898
rect 514944 368834 514996 368840
rect 514956 300490 514984 368834
rect 515128 355428 515180 355434
rect 515128 355370 515180 355376
rect 515036 352028 515088 352034
rect 515036 351970 515088 351976
rect 514944 300484 514996 300490
rect 514944 300426 514996 300432
rect 514852 300416 514904 300422
rect 514852 300358 514904 300364
rect 514760 295316 514812 295322
rect 514760 295258 514812 295264
rect 514208 295248 514260 295254
rect 514208 295190 514260 295196
rect 513656 295112 513708 295118
rect 513656 295054 513708 295060
rect 515048 289678 515076 351970
rect 515140 303074 515168 355370
rect 515220 353388 515272 353394
rect 515220 353330 515272 353336
rect 515128 303068 515180 303074
rect 515128 303010 515180 303016
rect 515232 303006 515260 353330
rect 515312 349240 515364 349246
rect 515312 349182 515364 349188
rect 515324 303278 515352 349182
rect 515416 321162 515444 524418
rect 515496 461712 515548 461718
rect 515496 461654 515548 461660
rect 515404 321156 515456 321162
rect 515404 321098 515456 321104
rect 515508 319802 515536 461654
rect 518164 383036 518216 383042
rect 518164 382978 518216 382984
rect 515588 382492 515640 382498
rect 515588 382434 515640 382440
rect 515600 358494 515628 382434
rect 517520 376848 517572 376854
rect 517520 376790 517572 376796
rect 516140 375420 516192 375426
rect 516140 375362 516192 375368
rect 515588 358488 515640 358494
rect 515588 358430 515640 358436
rect 515588 342576 515640 342582
rect 515588 342518 515640 342524
rect 515496 319796 515548 319802
rect 515496 319738 515548 319744
rect 515312 303272 515364 303278
rect 515312 303214 515364 303220
rect 515220 303000 515272 303006
rect 515220 302942 515272 302948
rect 515600 297838 515628 342518
rect 516152 300354 516180 375362
rect 516232 368552 516284 368558
rect 516232 368494 516284 368500
rect 516140 300348 516192 300354
rect 516140 300290 516192 300296
rect 515588 297832 515640 297838
rect 515588 297774 515640 297780
rect 516244 295186 516272 368494
rect 516784 365764 516836 365770
rect 516784 365706 516836 365712
rect 516416 358896 516468 358902
rect 516416 358838 516468 358844
rect 516324 353524 516376 353530
rect 516324 353466 516376 353472
rect 516232 295180 516284 295186
rect 516232 295122 516284 295128
rect 516336 289814 516364 353466
rect 516428 294846 516456 358838
rect 516600 352708 516652 352714
rect 516600 352650 516652 352656
rect 516508 349852 516560 349858
rect 516508 349794 516560 349800
rect 516416 294840 516468 294846
rect 516416 294782 516468 294788
rect 516324 289808 516376 289814
rect 516324 289750 516376 289756
rect 515036 289672 515088 289678
rect 515036 289614 515088 289620
rect 516520 289542 516548 349794
rect 516612 294710 516640 352650
rect 516692 347812 516744 347818
rect 516692 347754 516744 347760
rect 516704 297634 516732 347754
rect 516796 320890 516824 365706
rect 516876 341148 516928 341154
rect 516876 341090 516928 341096
rect 516784 320884 516836 320890
rect 516784 320826 516836 320832
rect 516888 297702 516916 341090
rect 516968 337204 517020 337210
rect 516968 337146 517020 337152
rect 516980 297906 517008 337146
rect 517532 300218 517560 376790
rect 517704 373380 517756 373386
rect 517704 373322 517756 373328
rect 517612 363316 517664 363322
rect 517612 363258 517664 363264
rect 517520 300212 517572 300218
rect 517520 300154 517572 300160
rect 516968 297900 517020 297906
rect 516968 297842 517020 297848
rect 516876 297696 516928 297702
rect 516876 297638 516928 297644
rect 516692 297628 516744 297634
rect 516692 297570 516744 297576
rect 516600 294704 516652 294710
rect 516600 294646 516652 294652
rect 516508 289536 516560 289542
rect 516508 289478 516560 289484
rect 517624 289338 517652 363258
rect 517716 300286 517744 373322
rect 517796 365900 517848 365906
rect 517796 365842 517848 365848
rect 517704 300280 517756 300286
rect 517704 300222 517756 300228
rect 517808 294914 517836 365842
rect 518176 358698 518204 382978
rect 518900 374060 518952 374066
rect 518900 374002 518952 374008
rect 518164 358692 518216 358698
rect 518164 358634 518216 358640
rect 517888 357740 517940 357746
rect 517888 357682 517940 357688
rect 517796 294908 517848 294914
rect 517796 294850 517848 294856
rect 517900 294778 517928 357682
rect 517980 354748 518032 354754
rect 517980 354690 518032 354696
rect 517888 294772 517940 294778
rect 517888 294714 517940 294720
rect 517992 294642 518020 354690
rect 518072 350940 518124 350946
rect 518072 350882 518124 350888
rect 518084 297430 518112 350882
rect 518164 344276 518216 344282
rect 518164 344218 518216 344224
rect 518072 297424 518124 297430
rect 518072 297366 518124 297372
rect 518176 297294 518204 344218
rect 518256 339516 518308 339522
rect 518256 339458 518308 339464
rect 518268 297498 518296 339458
rect 518348 336116 518400 336122
rect 518348 336058 518400 336064
rect 518360 300150 518388 336058
rect 518348 300144 518400 300150
rect 518348 300086 518400 300092
rect 518256 297492 518308 297498
rect 518256 297434 518308 297440
rect 518164 297288 518216 297294
rect 518164 297230 518216 297236
rect 517980 294636 518032 294642
rect 517980 294578 518032 294584
rect 518912 291922 518940 374002
rect 518992 372700 519044 372706
rect 518992 372642 519044 372648
rect 519004 294982 519032 372642
rect 519084 356380 519136 356386
rect 519084 356322 519136 356328
rect 518992 294976 519044 294982
rect 518992 294918 519044 294924
rect 518900 291916 518952 291922
rect 518900 291858 518952 291864
rect 519096 289610 519124 356322
rect 519176 347948 519228 347954
rect 519176 347890 519228 347896
rect 519188 292466 519216 347890
rect 519268 341284 519320 341290
rect 519268 341226 519320 341232
rect 519176 292460 519228 292466
rect 519176 292402 519228 292408
rect 519280 292262 519308 341226
rect 519452 334212 519504 334218
rect 519452 334154 519504 334160
rect 519360 331492 519412 331498
rect 519360 331434 519412 331440
rect 519268 292256 519320 292262
rect 519268 292198 519320 292204
rect 519084 289604 519136 289610
rect 519084 289546 519136 289552
rect 519372 289474 519400 331434
rect 519464 292126 519492 334154
rect 519556 322998 519584 598130
rect 538220 515432 538272 515438
rect 538220 515374 538272 515380
rect 535460 512032 535512 512038
rect 535460 511974 535512 511980
rect 532700 508564 532752 508570
rect 532700 508506 532752 508512
rect 529940 505164 529992 505170
rect 529940 505106 529992 505112
rect 529952 480254 529980 505106
rect 532712 480254 532740 508506
rect 535472 480254 535500 511974
rect 538232 480254 538260 515374
rect 529952 480226 530256 480254
rect 532712 480226 533200 480254
rect 535472 480226 536144 480254
rect 538232 480226 539088 480254
rect 527640 462528 527692 462534
rect 527640 462470 527692 462476
rect 521752 461644 521804 461650
rect 521752 461586 521804 461592
rect 521764 460972 521792 461586
rect 524432 460970 524722 460986
rect 527652 460972 527680 462470
rect 530228 460986 530256 480226
rect 533172 460986 533200 480226
rect 536116 460986 536144 480226
rect 539060 460986 539088 480226
rect 542372 461718 542400 702406
rect 559668 699825 559696 703520
rect 559654 699816 559710 699825
rect 559654 699751 559710 699760
rect 580262 697232 580318 697241
rect 580262 697167 580318 697176
rect 579618 644056 579674 644065
rect 579618 643991 579674 644000
rect 579632 643142 579660 643991
rect 569224 643136 569276 643142
rect 569224 643078 569276 643084
rect 579620 643136 579672 643142
rect 579620 643078 579672 643084
rect 567844 630692 567896 630698
rect 567844 630634 567896 630640
rect 545120 500268 545172 500274
rect 545120 500210 545172 500216
rect 542452 498908 542504 498914
rect 542452 498850 542504 498856
rect 542360 461712 542412 461718
rect 542360 461654 542412 461660
rect 542464 460986 542492 498850
rect 524420 460964 524722 460970
rect 524472 460958 524722 460964
rect 530228 460958 530610 460986
rect 533172 460958 533554 460986
rect 536116 460958 536498 460986
rect 539060 460958 539442 460986
rect 542386 460958 542492 460986
rect 545132 460986 545160 500210
rect 547880 498840 547932 498846
rect 547880 498782 547932 498788
rect 547892 460986 547920 498782
rect 554136 462460 554188 462466
rect 554136 462402 554188 462408
rect 551192 462392 551244 462398
rect 551192 462334 551244 462340
rect 545132 460958 545330 460986
rect 547892 460958 548274 460986
rect 551204 460972 551232 462334
rect 554148 460972 554176 462402
rect 524420 460906 524472 460912
rect 557538 442912 557594 442921
rect 557538 442847 557594 442856
rect 521212 421598 521240 425068
rect 522304 423496 522356 423502
rect 522304 423438 522356 423444
rect 521200 421592 521252 421598
rect 521200 421534 521252 421540
rect 522316 388822 522344 423438
rect 522500 423434 522528 425068
rect 523788 423570 523816 425068
rect 524708 425054 525090 425082
rect 523776 423564 523828 423570
rect 523776 423506 523828 423512
rect 522488 423428 522540 423434
rect 522488 423370 522540 423376
rect 523684 423428 523736 423434
rect 523684 423370 523736 423376
rect 523696 388890 523724 423370
rect 524708 412634 524736 425054
rect 526364 423366 526392 425068
rect 527284 425054 527666 425082
rect 526352 423360 526404 423366
rect 526352 423302 526404 423308
rect 526444 423360 526496 423366
rect 526444 423302 526496 423308
rect 524432 412606 524736 412634
rect 523684 388884 523736 388890
rect 523684 388826 523736 388832
rect 522304 388816 522356 388822
rect 522304 388758 522356 388764
rect 524432 388686 524460 412606
rect 526456 388754 526484 423302
rect 527284 412634 527312 425054
rect 528940 423298 528968 425068
rect 530228 423638 530256 425068
rect 529204 423632 529256 423638
rect 529204 423574 529256 423580
rect 530216 423632 530268 423638
rect 530216 423574 530268 423580
rect 530584 423632 530636 423638
rect 530584 423574 530636 423580
rect 528928 423292 528980 423298
rect 528928 423234 528980 423240
rect 527192 412606 527312 412634
rect 526444 388748 526496 388754
rect 526444 388690 526496 388696
rect 524420 388680 524472 388686
rect 524420 388622 524472 388628
rect 527192 388618 527220 412606
rect 527180 388612 527232 388618
rect 527180 388554 527232 388560
rect 529216 388482 529244 423574
rect 530596 388550 530624 423574
rect 531516 423230 531544 425068
rect 532804 423638 532832 425068
rect 532792 423632 532844 423638
rect 532792 423574 532844 423580
rect 531504 423224 531556 423230
rect 531504 423166 531556 423172
rect 534092 392630 534120 425068
rect 535012 425054 535394 425082
rect 536300 425054 536682 425082
rect 537588 425054 537970 425082
rect 538876 425054 539258 425082
rect 540164 425054 540546 425082
rect 535012 412634 535040 425054
rect 536300 412634 536328 425054
rect 537588 412634 537616 425054
rect 538876 412634 538904 425054
rect 540164 412634 540192 425054
rect 541820 420238 541848 425068
rect 542740 425054 543122 425082
rect 544028 425054 544410 425082
rect 541808 420232 541860 420238
rect 541808 420174 541860 420180
rect 542740 412634 542768 425054
rect 544028 412634 544056 425054
rect 545684 423162 545712 425068
rect 546604 425054 546986 425082
rect 545672 423156 545724 423162
rect 545672 423098 545724 423104
rect 546604 412634 546632 425054
rect 548260 423094 548288 425068
rect 549548 423502 549576 425068
rect 549536 423496 549588 423502
rect 549536 423438 549588 423444
rect 548248 423088 548300 423094
rect 548248 423030 548300 423036
rect 550836 423026 550864 425068
rect 552124 423434 552152 425068
rect 552112 423428 552164 423434
rect 552112 423370 552164 423376
rect 550824 423020 550876 423026
rect 550824 422962 550876 422968
rect 553412 422958 553440 425068
rect 554700 423366 554728 425068
rect 554688 423360 554740 423366
rect 554688 423302 554740 423308
rect 553400 422952 553452 422958
rect 553400 422894 553452 422900
rect 534184 412606 535040 412634
rect 535472 412606 536328 412634
rect 536852 412606 537616 412634
rect 538232 412606 538904 412634
rect 539612 412606 540192 412634
rect 542372 412606 542768 412634
rect 543752 412606 544056 412634
rect 546512 412606 546632 412634
rect 534184 393990 534212 412606
rect 535472 395350 535500 412606
rect 536852 396778 536880 412606
rect 538232 398138 538260 412606
rect 539612 399498 539640 412606
rect 539600 399492 539652 399498
rect 539600 399434 539652 399440
rect 538220 398132 538272 398138
rect 538220 398074 538272 398080
rect 536840 396772 536892 396778
rect 536840 396714 536892 396720
rect 535460 395344 535512 395350
rect 535460 395286 535512 395292
rect 534172 393984 534224 393990
rect 534172 393926 534224 393932
rect 534080 392624 534132 392630
rect 534080 392566 534132 392572
rect 542372 389910 542400 412606
rect 543752 391338 543780 412606
rect 546512 400926 546540 412606
rect 557552 402286 557580 442847
rect 557540 402280 557592 402286
rect 557540 402222 557592 402228
rect 546500 400920 546552 400926
rect 546500 400862 546552 400868
rect 543740 391332 543792 391338
rect 543740 391274 543792 391280
rect 542360 389904 542412 389910
rect 542360 389846 542412 389852
rect 530584 388544 530636 388550
rect 530584 388486 530636 388492
rect 529204 388476 529256 388482
rect 529204 388418 529256 388424
rect 553952 386640 554004 386646
rect 553952 386582 554004 386588
rect 530584 383784 530636 383790
rect 530584 383726 530636 383732
rect 519636 382424 519688 382430
rect 519636 382366 519688 382372
rect 519648 358630 519676 382366
rect 522304 378344 522356 378350
rect 522304 378286 522356 378292
rect 520280 375556 520332 375562
rect 520280 375498 520332 375504
rect 519636 358624 519688 358630
rect 519636 358566 519688 358572
rect 519728 338292 519780 338298
rect 519728 338234 519780 338240
rect 519636 332716 519688 332722
rect 519636 332658 519688 332664
rect 519544 322992 519596 322998
rect 519544 322934 519596 322940
rect 519452 292120 519504 292126
rect 519452 292062 519504 292068
rect 519648 292058 519676 332658
rect 519740 304434 519768 338234
rect 519728 304428 519780 304434
rect 519728 304370 519780 304376
rect 519636 292052 519688 292058
rect 519636 291994 519688 292000
rect 520292 291854 520320 375498
rect 520372 367396 520424 367402
rect 520372 367338 520424 367344
rect 520280 291848 520332 291854
rect 520280 291790 520332 291796
rect 519360 289468 519412 289474
rect 519360 289410 519412 289416
rect 517612 289332 517664 289338
rect 517612 289274 517664 289280
rect 520384 289202 520412 367338
rect 520464 360256 520516 360262
rect 520464 360198 520516 360204
rect 520476 289746 520504 360198
rect 522316 358970 522344 378286
rect 523040 372632 523092 372638
rect 523040 372574 523092 372580
rect 522304 358964 522356 358970
rect 522304 358906 522356 358912
rect 520556 355020 520608 355026
rect 520556 354962 520608 354968
rect 520464 289740 520516 289746
rect 520464 289682 520516 289688
rect 520568 289406 520596 354962
rect 520648 345228 520700 345234
rect 520648 345170 520700 345176
rect 520660 292398 520688 345170
rect 520740 343868 520792 343874
rect 520740 343810 520792 343816
rect 520648 292392 520700 292398
rect 520648 292334 520700 292340
rect 520752 292330 520780 343810
rect 521660 342304 521712 342310
rect 521660 342246 521712 342252
rect 520832 339652 520884 339658
rect 520832 339594 520884 339600
rect 520740 292324 520792 292330
rect 520740 292266 520792 292272
rect 520844 292194 520872 339594
rect 520924 336932 520976 336938
rect 520924 336874 520976 336880
rect 520832 292188 520884 292194
rect 520832 292130 520884 292136
rect 520936 291990 520964 336874
rect 520924 291984 520976 291990
rect 520924 291926 520976 291932
rect 520556 289400 520608 289406
rect 520556 289342 520608 289348
rect 520372 289196 520424 289202
rect 520372 289138 520424 289144
rect 521672 286482 521700 342246
rect 521752 338156 521804 338162
rect 521752 338098 521804 338104
rect 521660 286476 521712 286482
rect 521660 286418 521712 286424
rect 521764 286414 521792 338098
rect 521844 335368 521896 335374
rect 521844 335310 521896 335316
rect 521856 286550 521884 335310
rect 523052 289134 523080 372574
rect 530596 358902 530624 383726
rect 547144 383716 547196 383722
rect 547144 383658 547196 383664
rect 544384 379568 544436 379574
rect 544384 379510 544436 379516
rect 544396 359106 544424 379510
rect 544384 359100 544436 359106
rect 544384 359042 544436 359048
rect 547156 359038 547184 383658
rect 549904 380928 549956 380934
rect 549904 380870 549956 380876
rect 548524 378276 548576 378282
rect 548524 378218 548576 378224
rect 547236 376032 547288 376038
rect 547236 375974 547288 375980
rect 547144 359032 547196 359038
rect 547144 358974 547196 358980
rect 530584 358896 530636 358902
rect 530584 358838 530636 358844
rect 547248 358562 547276 375974
rect 548536 360194 548564 378218
rect 548524 360188 548576 360194
rect 548524 360130 548576 360136
rect 549916 359174 549944 380870
rect 553964 377890 553992 386582
rect 563428 385144 563480 385150
rect 563428 385086 563480 385092
rect 553964 377862 554438 377890
rect 563440 377876 563468 385086
rect 549996 377460 550048 377466
rect 549996 377402 550048 377408
rect 549904 359168 549956 359174
rect 549904 359110 549956 359116
rect 550008 358766 550036 377402
rect 552032 360194 552322 360210
rect 552020 360188 552322 360194
rect 552072 360182 552322 360188
rect 552020 360130 552072 360136
rect 550836 358970 550864 360060
rect 553780 359106 553808 360060
rect 553768 359100 553820 359106
rect 553768 359042 553820 359048
rect 550824 358964 550876 358970
rect 550824 358906 550876 358912
rect 555252 358834 555280 360060
rect 555240 358828 555292 358834
rect 555240 358770 555292 358776
rect 556724 358766 556752 360060
rect 558196 359174 558224 360060
rect 558184 359168 558236 359174
rect 558184 359110 558236 359116
rect 549996 358760 550048 358766
rect 549996 358702 550048 358708
rect 556712 358760 556764 358766
rect 556712 358702 556764 358708
rect 559668 358562 559696 360060
rect 547236 358556 547288 358562
rect 547236 358498 547288 358504
rect 559656 358556 559708 358562
rect 559656 358498 559708 358504
rect 561140 358494 561168 360060
rect 562612 358698 562640 360060
rect 562600 358692 562652 358698
rect 562600 358634 562652 358640
rect 564084 358630 564112 360060
rect 565556 359038 565584 360060
rect 565544 359032 565596 359038
rect 565544 358974 565596 358980
rect 567028 358902 567056 360060
rect 567016 358896 567068 358902
rect 567016 358838 567068 358844
rect 564072 358624 564124 358630
rect 564072 358566 564124 358572
rect 561128 358488 561180 358494
rect 561128 358430 561180 358436
rect 523132 336796 523184 336802
rect 523132 336738 523184 336744
rect 523040 289128 523092 289134
rect 523040 289070 523092 289076
rect 521844 286544 521896 286550
rect 521844 286486 521896 286492
rect 521752 286408 521804 286414
rect 521752 286350 521804 286356
rect 523144 286346 523172 336738
rect 567856 321298 567884 630634
rect 567936 590708 567988 590714
rect 567936 590650 567988 590656
rect 567844 321292 567896 321298
rect 567844 321234 567896 321240
rect 567948 319870 567976 590650
rect 569236 319938 569264 643078
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 571984 616888 572036 616894
rect 571984 616830 572036 616836
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 569316 484424 569368 484430
rect 569316 484366 569368 484372
rect 569328 320006 569356 484366
rect 569408 430636 569460 430642
rect 569408 430578 569460 430584
rect 569420 321230 569448 430578
rect 569500 364404 569552 364410
rect 569500 364346 569552 364352
rect 569512 321366 569540 364346
rect 569500 321360 569552 321366
rect 569500 321302 569552 321308
rect 569408 321224 569460 321230
rect 569408 321166 569460 321172
rect 569316 320000 569368 320006
rect 569316 319942 569368 319948
rect 569224 319932 569276 319938
rect 569224 319874 569276 319880
rect 567936 319864 567988 319870
rect 567936 319806 567988 319812
rect 543740 319456 543792 319462
rect 543740 319398 543792 319404
rect 540980 318096 541032 318102
rect 540980 318038 541032 318044
rect 539140 317076 539192 317082
rect 539140 317018 539192 317024
rect 529940 313948 529992 313954
rect 529940 313890 529992 313896
rect 529204 301640 529256 301646
rect 529204 301582 529256 301588
rect 529216 287054 529244 301582
rect 529216 287026 529336 287054
rect 523132 286340 523184 286346
rect 523132 286282 523184 286288
rect 512000 276684 512052 276690
rect 512000 276626 512052 276632
rect 510620 269816 510672 269822
rect 510620 269758 510672 269764
rect 500224 268524 500276 268530
rect 500224 268466 500276 268472
rect 499396 268456 499448 268462
rect 499396 268398 499448 268404
rect 487804 268388 487856 268394
rect 487804 268330 487856 268336
rect 494704 268388 494756 268394
rect 494704 268330 494756 268336
rect 529308 261633 529336 287026
rect 529294 261624 529350 261633
rect 529294 261559 529350 261568
rect 529952 209273 529980 313890
rect 530032 303612 530084 303618
rect 530032 303554 530084 303560
rect 530044 226250 530072 303554
rect 537484 301572 537536 301578
rect 537484 301514 537536 301520
rect 536104 293276 536156 293282
rect 536104 293218 536156 293224
rect 533344 290488 533396 290494
rect 533344 290430 533396 290436
rect 531320 284980 531372 284986
rect 531320 284922 531372 284928
rect 531332 243681 531360 284922
rect 531318 243672 531374 243681
rect 531318 243607 531374 243616
rect 530122 226264 530178 226273
rect 530044 226222 530122 226250
rect 530122 226199 530178 226208
rect 529938 209264 529994 209273
rect 529938 209199 529994 209208
rect 485780 200796 485832 200802
rect 485780 200738 485832 200744
rect 462964 200184 463016 200190
rect 462964 200126 463016 200132
rect 461584 196648 461636 196654
rect 461584 196590 461636 196596
rect 460296 133816 460348 133822
rect 460296 133758 460348 133764
rect 461596 41410 461624 196590
rect 461676 160132 461728 160138
rect 461676 160074 461728 160080
rect 461688 142934 461716 160074
rect 461676 142928 461728 142934
rect 461676 142870 461728 142876
rect 462504 67584 462556 67590
rect 462318 67552 462374 67561
rect 462318 67487 462374 67496
rect 462502 67552 462504 67561
rect 462556 67552 462558 67561
rect 462502 67487 462558 67496
rect 461584 41404 461636 41410
rect 461584 41346 461636 41352
rect 460204 31748 460256 31754
rect 460204 31690 460256 31696
rect 462332 31686 462360 67487
rect 462976 34474 463004 200126
rect 481640 199436 481692 199442
rect 481640 199378 481692 199384
rect 481652 140826 481680 199378
rect 464344 140820 464396 140826
rect 464344 140762 464396 140768
rect 481640 140820 481692 140826
rect 481640 140762 481692 140768
rect 464356 67590 464384 140762
rect 481652 139890 481680 140762
rect 485792 139890 485820 200738
rect 528560 195288 528612 195294
rect 528560 195230 528612 195236
rect 524420 171828 524472 171834
rect 524420 171770 524472 171776
rect 496820 161900 496872 161906
rect 496820 161842 496872 161848
rect 494060 161764 494112 161770
rect 494060 161706 494112 161712
rect 489920 142928 489972 142934
rect 489920 142870 489972 142876
rect 489932 139890 489960 142870
rect 494072 139890 494100 161706
rect 496832 151814 496860 161842
rect 500960 161832 501012 161838
rect 500960 161774 501012 161780
rect 500972 151814 501000 161774
rect 505100 161696 505152 161702
rect 505100 161638 505152 161644
rect 505112 151814 505140 161638
rect 513380 161628 513432 161634
rect 513380 161570 513432 161576
rect 513392 151814 513420 161570
rect 517520 161560 517572 161566
rect 517520 161502 517572 161508
rect 496832 151786 497688 151814
rect 500972 151786 501644 151814
rect 505112 151786 505600 151814
rect 513392 151786 513512 151814
rect 497660 139890 497688 151786
rect 501616 139890 501644 151786
rect 505572 139890 505600 151786
rect 509608 142860 509660 142866
rect 509608 142802 509660 142808
rect 509620 139890 509648 142802
rect 513484 139890 513512 151786
rect 517532 139890 517560 161502
rect 521660 160744 521712 160750
rect 521660 160686 521712 160692
rect 521672 139890 521700 160686
rect 524432 151814 524460 171770
rect 528572 151814 528600 195230
rect 533356 167006 533384 290430
rect 533344 167000 533396 167006
rect 533344 166942 533396 166948
rect 532700 161492 532752 161498
rect 532700 161434 532752 161440
rect 532712 151814 532740 161434
rect 536116 153202 536144 293218
rect 537496 179382 537524 301514
rect 537484 179376 537536 179382
rect 537484 179318 537536 179324
rect 536840 159384 536892 159390
rect 536840 159326 536892 159332
rect 536104 153196 536156 153202
rect 536104 153138 536156 153144
rect 536852 151814 536880 159326
rect 524432 151786 525380 151814
rect 528572 151786 529336 151814
rect 532712 151786 533292 151814
rect 536852 151786 537248 151814
rect 525352 139890 525380 151786
rect 529308 139890 529336 151786
rect 533264 139890 533292 151786
rect 537220 139890 537248 151786
rect 481652 139862 482264 139890
rect 485792 139862 486220 139890
rect 489932 139862 490176 139890
rect 494072 139862 494132 139890
rect 497660 139862 498088 139890
rect 501616 139862 502044 139890
rect 505572 139862 506000 139890
rect 509620 139862 509956 139890
rect 513484 139862 513912 139890
rect 517532 139862 517868 139890
rect 521672 139862 521824 139890
rect 525352 139862 525780 139890
rect 529308 139862 529736 139890
rect 533264 139862 533692 139890
rect 537220 139862 537648 139890
rect 539152 135674 539180 317018
rect 539600 314016 539652 314022
rect 539600 313958 539652 313964
rect 539232 283756 539284 283762
rect 539232 283698 539284 283704
rect 539244 151814 539272 283698
rect 539244 151786 539364 151814
rect 539336 137737 539364 151786
rect 539322 137728 539378 137737
rect 539322 137663 539378 137672
rect 539322 135688 539378 135697
rect 539152 135646 539322 135674
rect 539322 135623 539378 135632
rect 539612 99249 539640 313958
rect 539876 276820 539928 276826
rect 539876 276762 539928 276768
rect 539784 276752 539836 276758
rect 539784 276694 539836 276700
rect 539692 271380 539744 271386
rect 539692 271322 539744 271328
rect 539598 99240 539654 99249
rect 539598 99175 539654 99184
rect 539704 86873 539732 271322
rect 539796 100609 539824 276694
rect 539888 109177 539916 276762
rect 540060 274100 540112 274106
rect 540060 274042 540112 274048
rect 539968 272604 540020 272610
rect 539968 272546 540020 272552
rect 539980 112849 540008 272546
rect 540072 117337 540100 274042
rect 540336 271448 540388 271454
rect 540336 271390 540388 271396
rect 540244 270088 540296 270094
rect 540244 270030 540296 270036
rect 540152 268524 540204 268530
rect 540152 268466 540204 268472
rect 540164 125225 540192 268466
rect 540256 127265 540284 270030
rect 540348 133385 540376 271390
rect 540334 133376 540390 133385
rect 540334 133311 540390 133320
rect 540242 127256 540298 127265
rect 540242 127191 540298 127200
rect 540150 125216 540206 125225
rect 540150 125151 540206 125160
rect 540058 117328 540114 117337
rect 540058 117263 540114 117272
rect 539966 112840 540022 112849
rect 539966 112775 540022 112784
rect 539874 109168 539930 109177
rect 539874 109103 539930 109112
rect 539782 100600 539838 100609
rect 539782 100535 539838 100544
rect 539690 86864 539746 86873
rect 539690 86799 539746 86808
rect 540992 82385 541020 318038
rect 542452 317008 542504 317014
rect 542452 316950 542504 316956
rect 541072 316940 541124 316946
rect 541072 316882 541124 316888
rect 541084 102785 541112 316882
rect 541164 315512 541216 315518
rect 541164 315454 541216 315460
rect 541176 110945 541204 315454
rect 541532 278044 541584 278050
rect 541532 277986 541584 277992
rect 541440 275460 541492 275466
rect 541440 275402 541492 275408
rect 541256 275392 541308 275398
rect 541256 275334 541308 275340
rect 541162 110936 541218 110945
rect 541162 110871 541218 110880
rect 541070 102776 541126 102785
rect 541070 102711 541126 102720
rect 541268 88505 541296 275334
rect 541348 274032 541400 274038
rect 541348 273974 541400 273980
rect 541360 104825 541388 273974
rect 541452 106865 541480 275402
rect 541544 115025 541572 277986
rect 542464 121145 542492 316950
rect 543188 316872 543240 316878
rect 543188 316814 543240 316820
rect 542728 315580 542780 315586
rect 542728 315522 542780 315528
rect 542636 273964 542688 273970
rect 542636 273906 542688 273912
rect 542544 268388 542596 268394
rect 542544 268330 542596 268336
rect 542450 121136 542506 121145
rect 542450 121071 542506 121080
rect 541530 115016 541586 115025
rect 541530 114951 541586 114960
rect 541438 106856 541494 106865
rect 541438 106791 541494 106800
rect 541346 104816 541402 104825
rect 541346 104751 541402 104760
rect 541254 88496 541310 88505
rect 541254 88431 541310 88440
rect 542556 84425 542584 268330
rect 542648 90545 542676 273906
rect 542740 131345 542768 315522
rect 542820 275324 542872 275330
rect 542820 275266 542872 275272
rect 542726 131336 542782 131345
rect 542726 131271 542782 131280
rect 542832 92585 542860 275266
rect 542912 272536 542964 272542
rect 542912 272478 542964 272484
rect 542924 96665 542952 272478
rect 543096 270020 543148 270026
rect 543096 269962 543148 269968
rect 543004 268456 543056 268462
rect 543004 268398 543056 268404
rect 543016 119105 543044 268398
rect 543108 123185 543136 269962
rect 543094 123176 543150 123185
rect 543094 123111 543150 123120
rect 543002 119096 543058 119105
rect 543002 119031 543058 119040
rect 542910 96656 542966 96665
rect 542910 96591 542966 96600
rect 543200 94625 543228 316814
rect 543186 94616 543242 94625
rect 543186 94551 543242 94560
rect 542818 92576 542874 92585
rect 542818 92511 542874 92520
rect 542634 90536 542690 90545
rect 542634 90471 542690 90480
rect 542542 84416 542598 84425
rect 542542 84351 542598 84360
rect 540978 82376 541034 82385
rect 540978 82311 541034 82320
rect 464344 67584 464396 67590
rect 464344 67526 464396 67532
rect 543752 51134 543780 319398
rect 571996 318646 572024 616830
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 590714 580212 590951
rect 580172 590708 580224 590714
rect 580172 590650 580224 590656
rect 579618 564360 579674 564369
rect 579618 564295 579674 564304
rect 579632 563106 579660 564295
rect 577504 563100 577556 563106
rect 577504 563042 577556 563048
rect 579620 563100 579672 563106
rect 579620 563042 579672 563048
rect 577516 318714 577544 563042
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 578882 458144 578938 458153
rect 578882 458079 578938 458088
rect 578896 318782 578924 458079
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 579802 378448 579858 378457
rect 579802 378383 579858 378392
rect 579816 378214 579844 378383
rect 579804 378208 579856 378214
rect 579804 378150 579856 378156
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580184 364410 580212 365055
rect 580172 364404 580224 364410
rect 580172 364346 580224 364352
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 580184 325694 580212 351863
rect 580276 333266 580304 697167
rect 580354 683904 580410 683913
rect 580354 683839 580410 683848
rect 580264 333260 580316 333266
rect 580264 333202 580316 333208
rect 580092 325666 580212 325694
rect 580092 321502 580120 325666
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 322250 580212 325207
rect 580368 322318 580396 683839
rect 580446 670712 580502 670721
rect 580446 670647 580502 670656
rect 580356 322312 580408 322318
rect 580356 322254 580408 322260
rect 580172 322244 580224 322250
rect 580172 322186 580224 322192
rect 580080 321496 580132 321502
rect 580080 321438 580132 321444
rect 580460 321434 580488 670647
rect 580538 577688 580594 577697
rect 580538 577623 580594 577632
rect 580552 322386 580580 577623
rect 580630 537840 580686 537849
rect 580630 537775 580686 537784
rect 580644 322454 580672 537775
rect 580722 511320 580778 511329
rect 580722 511255 580778 511264
rect 580632 322448 580684 322454
rect 580632 322390 580684 322396
rect 580540 322380 580592 322386
rect 580540 322322 580592 322328
rect 580448 321428 580500 321434
rect 580448 321370 580500 321376
rect 580736 319326 580764 511255
rect 580814 418296 580870 418305
rect 580814 418231 580870 418240
rect 580828 320074 580856 418231
rect 580906 404968 580962 404977
rect 580906 404903 580962 404912
rect 580920 321570 580948 404903
rect 580908 321564 580960 321570
rect 580908 321506 580960 321512
rect 580816 320068 580868 320074
rect 580816 320010 580868 320016
rect 580724 319320 580776 319326
rect 580724 319262 580776 319268
rect 578884 318776 578936 318782
rect 578884 318718 578936 318724
rect 577504 318708 577556 318714
rect 577504 318650 577556 318656
rect 571984 318640 572036 318646
rect 571984 318582 572036 318588
rect 570604 315308 570656 315314
rect 570604 315250 570656 315256
rect 551284 312588 551336 312594
rect 551284 312530 551336 312536
rect 544384 311160 544436 311166
rect 544384 311102 544436 311108
rect 544396 73166 544424 311102
rect 548524 297220 548576 297226
rect 548524 297162 548576 297168
rect 547144 285048 547196 285054
rect 547144 284990 547196 284996
rect 544384 73160 544436 73166
rect 544384 73102 544436 73108
rect 547156 60722 547184 284990
rect 548536 193186 548564 297162
rect 548524 193180 548576 193186
rect 548524 193122 548576 193128
rect 551296 100706 551324 312530
rect 563704 309800 563756 309806
rect 563704 309742 563756 309748
rect 562324 308440 562376 308446
rect 562324 308382 562376 308388
rect 554044 269884 554096 269890
rect 554044 269826 554096 269832
rect 554056 139398 554084 269826
rect 554044 139392 554096 139398
rect 554044 139334 554096 139340
rect 551284 100700 551336 100706
rect 551284 100642 551336 100648
rect 547144 60716 547196 60722
rect 547144 60658 547196 60664
rect 540612 51128 540664 51134
rect 540612 51070 540664 51076
rect 543740 51128 543792 51134
rect 543740 51070 543792 51076
rect 540624 48929 540652 51070
rect 540610 48920 540666 48929
rect 540610 48855 540666 48864
rect 536840 41404 536892 41410
rect 536840 41346 536892 41352
rect 536852 41041 536880 41346
rect 536838 41032 536894 41041
rect 536838 40967 536894 40976
rect 462964 34468 463016 34474
rect 462964 34410 463016 34416
rect 536840 34468 536892 34474
rect 536840 34410 536892 34416
rect 536852 33697 536880 34410
rect 536838 33688 536894 33697
rect 536838 33623 536894 33632
rect 462320 31680 462372 31686
rect 462320 31622 462372 31628
rect 386052 31476 386104 31482
rect 386052 31418 386104 31424
rect 385960 31068 386012 31074
rect 385960 31010 386012 31016
rect 562336 20670 562364 308382
rect 563716 33114 563744 309742
rect 565084 305788 565136 305794
rect 565084 305730 565136 305736
rect 563704 33108 563756 33114
rect 563704 33050 563756 33056
rect 562324 20664 562376 20670
rect 562324 20606 562376 20612
rect 565096 6866 565124 305730
rect 569224 287700 569276 287706
rect 569224 287642 569276 287648
rect 566464 283620 566516 283626
rect 566464 283562 566516 283568
rect 566476 233238 566504 283562
rect 566464 233232 566516 233238
rect 566464 233174 566516 233180
rect 569236 219434 569264 287642
rect 569224 219428 569276 219434
rect 569224 219370 569276 219376
rect 570616 206990 570644 315250
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 573364 304496 573416 304502
rect 573364 304438 573416 304444
rect 571984 286680 572036 286686
rect 571984 286622 572036 286628
rect 570604 206984 570656 206990
rect 570604 206926 570656 206932
rect 571996 113150 572024 286622
rect 573376 245614 573404 304438
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 578884 295996 578936 296002
rect 578884 295938 578936 295944
rect 576124 294432 576176 294438
rect 576124 294374 576176 294380
rect 574744 291712 574796 291718
rect 574744 291654 574796 291660
rect 573364 245608 573416 245614
rect 573364 245550 573416 245556
rect 574756 126954 574784 291654
rect 574744 126948 574796 126954
rect 574744 126890 574796 126896
rect 571984 113144 572036 113150
rect 571984 113086 572036 113092
rect 576136 86970 576164 294374
rect 576124 86964 576176 86970
rect 576124 86906 576176 86912
rect 578896 46345 578924 295938
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580264 271176 580316 271182
rect 580264 271118 580316 271124
rect 580276 258913 580304 271118
rect 580262 258904 580318 258913
rect 580262 258839 580318 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 578882 46336 578938 46345
rect 578882 46271 578938 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 565084 6860 565136 6866
rect 565084 6802 565136 6808
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 385684 3460 385736 3466
rect 385684 3402 385736 3408
rect 384486 3360 384542 3369
rect 384486 3295 384542 3304
rect 384304 2100 384356 2106
rect 384304 2042 384356 2048
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3238 684256 3294 684312
rect 3054 682760 3110 682816
rect 3146 658180 3148 658200
rect 3148 658180 3200 658200
rect 3200 658180 3202 658200
rect 3146 658144 3202 658180
rect 3238 579944 3294 580000
rect 3330 566888 3386 566944
rect 3698 632032 3754 632088
rect 3606 475632 3662 475688
rect 3514 462576 3570 462632
rect 3422 449520 3478 449576
rect 6918 683712 6974 683768
rect 170310 700440 170366 700496
rect 137834 700304 137890 700360
rect 235170 700576 235226 700632
rect 201498 683984 201554 684040
rect 23478 683848 23534 683904
rect 4066 553832 4122 553888
rect 3974 527856 4030 527912
rect 3882 514800 3938 514856
rect 361762 678988 361764 679008
rect 361764 678988 361816 679008
rect 361816 678988 361818 679008
rect 361762 678952 361818 678988
rect 361762 667956 361818 667992
rect 361762 667936 361764 667956
rect 361764 667936 361816 667956
rect 361816 667936 361818 667956
rect 361762 656940 361818 656976
rect 361762 656920 361764 656940
rect 361764 656920 361816 656940
rect 361816 656920 361818 656940
rect 361762 645924 361818 645960
rect 361762 645904 361764 645924
rect 361764 645904 361816 645924
rect 361816 645904 361818 645924
rect 361578 634888 361634 634944
rect 361578 623872 361634 623928
rect 361578 612856 361634 612912
rect 361762 601840 361818 601896
rect 361762 590824 361818 590880
rect 361762 579808 361818 579864
rect 361762 568792 361818 568848
rect 361578 557796 361634 557832
rect 361578 557776 361580 557796
rect 361580 557776 361632 557796
rect 361632 557776 361634 557796
rect 361578 546760 361634 546816
rect 361578 535764 361634 535800
rect 361578 535744 361580 535764
rect 361580 535744 361632 535764
rect 361632 535744 361634 535764
rect 361762 524728 361818 524784
rect 3790 501744 3846 501800
rect 3698 423544 3754 423600
rect 361762 513712 361818 513768
rect 361762 502696 361818 502752
rect 362222 491680 362278 491736
rect 361762 480664 361818 480720
rect 361762 469648 361818 469704
rect 361762 458632 361818 458688
rect 361762 436600 361818 436656
rect 361578 414568 361634 414624
rect 3974 410488 4030 410544
rect 361578 403552 361634 403608
rect 3882 397432 3938 397488
rect 3422 358400 3478 358456
rect 3514 345344 3570 345400
rect 3422 293120 3478 293176
rect 3330 162832 3386 162888
rect 3238 149776 3294 149832
rect 3146 84632 3202 84688
rect 3146 71576 3202 71632
rect 3790 319232 3846 319288
rect 3698 306176 3754 306232
rect 3514 267144 3570 267200
rect 3422 59880 3478 59936
rect 3422 58520 3478 58576
rect 3606 254088 3662 254144
rect 361578 392536 361634 392592
rect 3974 371320 4030 371376
rect 3790 241032 3846 241088
rect 3698 97552 3754 97608
rect 3882 214920 3938 214976
rect 3974 201864 4030 201920
rect 4066 188808 4122 188864
rect 19338 49544 19394 49600
rect 3514 45484 3570 45520
rect 3514 45464 3516 45484
rect 3516 45464 3568 45484
rect 3568 45464 3570 45484
rect 21362 46688 21418 46744
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 46938 44784 46994 44840
rect 3422 6432 3478 6488
rect 1674 3304 1730 3360
rect 5262 3848 5318 3904
rect 8758 3712 8814 3768
rect 13542 3576 13598 3632
rect 17038 3984 17094 4040
rect 24214 3440 24270 3496
rect 361578 381520 361634 381576
rect 362314 447616 362370 447672
rect 362406 425584 362462 425640
rect 361578 370504 361634 370560
rect 362314 359488 362370 359544
rect 361762 348472 361818 348528
rect 361762 337456 361818 337512
rect 362222 326440 362278 326496
rect 361762 315424 361818 315480
rect 361762 304408 361818 304464
rect 361118 302776 361174 302832
rect 361026 3848 361082 3904
rect 361762 293392 361818 293448
rect 361762 282376 361818 282432
rect 361762 271360 361818 271416
rect 361762 260344 361818 260400
rect 361762 249328 361818 249384
rect 361762 238312 361818 238368
rect 361762 227296 361818 227352
rect 361670 216316 361672 216336
rect 361672 216316 361724 216336
rect 361724 216316 361726 216336
rect 361670 216280 361726 216316
rect 361762 205264 361818 205320
rect 361762 194248 361818 194304
rect 361762 183232 361818 183288
rect 361762 172216 361818 172272
rect 361762 161200 361818 161256
rect 361762 139168 361818 139224
rect 361762 128152 361818 128208
rect 361762 117136 361818 117192
rect 361762 106120 361818 106176
rect 361762 84124 361764 84144
rect 361764 84124 361816 84144
rect 361816 84124 361818 84144
rect 361762 84088 361818 84124
rect 361762 73108 361764 73128
rect 361764 73108 361816 73128
rect 361816 73108 361818 73128
rect 361762 73072 361818 73108
rect 361762 62076 361818 62112
rect 361762 62056 361764 62076
rect 361764 62056 361816 62076
rect 361816 62056 361818 62076
rect 361762 51076 361764 51096
rect 361764 51076 361816 51096
rect 361816 51076 361818 51096
rect 361762 51040 361818 51076
rect 361394 46416 361450 46472
rect 362590 150184 362646 150240
rect 362682 95104 362738 95160
rect 370502 305632 370558 305688
rect 368018 300056 368074 300112
rect 365166 3712 365222 3768
rect 370686 300192 370742 300248
rect 370686 3984 370742 4040
rect 372158 291760 372214 291816
rect 370502 3576 370558 3632
rect 376114 302912 376170 302968
rect 378598 46552 378654 46608
rect 384486 306176 384542 306232
rect 384302 306040 384358 306096
rect 381910 303048 381966 303104
rect 382186 303184 382242 303240
rect 383014 3440 383070 3496
rect 384670 305904 384726 305960
rect 384854 46960 384910 47016
rect 384762 46688 384818 46744
rect 385774 46824 385830 46880
rect 420274 682896 420330 682952
rect 420090 334600 420146 334656
rect 420734 334736 420790 334792
rect 420734 334464 420790 334520
rect 428094 334464 428150 334520
rect 421746 162696 421802 162752
rect 432602 332832 432658 332888
rect 432418 329160 432474 329216
rect 428646 162696 428702 162752
rect 432694 325488 432750 325544
rect 432878 321816 432934 321872
rect 432786 318144 432842 318200
rect 433246 314508 433248 314528
rect 433248 314508 433300 314528
rect 433300 314508 433302 314528
rect 433246 314472 433302 314508
rect 432602 310800 432658 310856
rect 432234 307128 432290 307184
rect 442446 334736 442502 334792
rect 445298 683304 445354 683360
rect 445482 321136 445538 321192
rect 446770 683168 446826 683224
rect 446770 319640 446826 319696
rect 447322 516160 447378 516216
rect 447690 507184 447746 507240
rect 447874 503376 447930 503432
rect 448518 516160 448574 516216
rect 448334 514256 448390 514312
rect 448242 512760 448298 512816
rect 448150 510448 448206 510504
rect 448058 505144 448114 505200
rect 447966 501880 448022 501936
rect 447138 383832 447194 383888
rect 447138 383152 447194 383208
rect 447230 382472 447286 382528
rect 447138 381792 447194 381848
rect 447230 381112 447286 381168
rect 447138 380432 447194 380488
rect 447230 379752 447286 379808
rect 447138 379072 447194 379128
rect 447230 378392 447286 378448
rect 447138 377712 447194 377768
rect 447230 377032 447286 377088
rect 447138 376352 447194 376408
rect 447230 375672 447286 375728
rect 447138 374992 447194 375048
rect 447230 374312 447286 374368
rect 447138 373632 447194 373688
rect 447230 372952 447286 373008
rect 447138 372272 447194 372328
rect 447230 371592 447286 371648
rect 447138 370912 447194 370968
rect 447230 370232 447286 370288
rect 447138 369552 447194 369608
rect 447230 368872 447286 368928
rect 447138 368192 447194 368248
rect 447230 367512 447286 367568
rect 447230 366832 447286 366888
rect 447138 366152 447194 366208
rect 447230 365472 447286 365528
rect 447138 364792 447194 364848
rect 447230 364112 447286 364168
rect 447138 363432 447194 363488
rect 447230 362752 447286 362808
rect 447138 362072 447194 362128
rect 447230 361392 447286 361448
rect 447138 360712 447194 360768
rect 447230 360032 447286 360088
rect 447138 359352 447194 359408
rect 447138 351908 447140 351928
rect 447140 351908 447192 351928
rect 447192 351908 447194 351928
rect 447138 351872 447194 351908
rect 447138 350548 447140 350568
rect 447140 350548 447192 350568
rect 447192 350548 447194 350568
rect 447138 350512 447194 350548
rect 447138 347112 447194 347168
rect 447690 353232 447746 353288
rect 447782 349152 447838 349208
rect 447322 343712 447378 343768
rect 447138 341672 447194 341728
rect 447230 341012 447286 341048
rect 447230 340992 447232 341012
rect 447232 340992 447284 341012
rect 447284 340992 447286 341012
rect 447138 340312 447194 340368
rect 447230 339632 447286 339688
rect 447230 338952 447286 339008
rect 447138 338272 447194 338328
rect 447230 337592 447286 337648
rect 447138 336912 447194 336968
rect 447230 336232 447286 336288
rect 447322 335552 447378 335608
rect 447322 334872 447378 334928
rect 447230 334192 447286 334248
rect 447322 333512 447378 333568
rect 447230 332832 447286 332888
rect 447230 331472 447286 331528
rect 447230 330792 447286 330848
rect 447230 330132 447286 330168
rect 447230 330112 447232 330132
rect 447232 330112 447284 330132
rect 447284 330112 447286 330132
rect 447230 329432 447286 329488
rect 447782 344392 447838 344448
rect 447598 332152 447654 332208
rect 447230 328752 447286 328808
rect 447230 328072 447286 328128
rect 447230 326032 447286 326088
rect 447322 323992 447378 324048
rect 448426 510448 448482 510504
rect 448978 357992 449034 358048
rect 448426 357312 448482 357368
rect 448426 351192 448482 351248
rect 448334 328072 448390 328128
rect 448242 327392 448298 327448
rect 448150 326712 448206 326768
rect 448058 325352 448114 325408
rect 447966 324672 448022 324728
rect 448242 324672 448298 324728
rect 448334 323992 448390 324048
rect 449070 342352 449126 342408
rect 527178 699760 527234 699816
rect 449806 503376 449862 503432
rect 449346 385600 449402 385656
rect 449438 356632 449494 356688
rect 449530 355272 449586 355328
rect 449622 354592 449678 354648
rect 449806 355952 449862 356008
rect 449714 353912 449770 353968
rect 449622 349832 449678 349888
rect 449346 323992 449402 324048
rect 450266 352960 450322 353016
rect 450174 348880 450230 348936
rect 450450 358808 450506 358864
rect 450358 348200 450414 348256
rect 449990 346840 450046 346896
rect 449898 346160 449954 346216
rect 449806 345072 449862 345128
rect 449714 343068 449716 343088
rect 449716 343068 449768 343088
rect 449768 343068 449770 343088
rect 449714 343032 449770 343068
rect 450542 334600 450598 334656
rect 449990 331608 450046 331664
rect 459650 667936 459706 667992
rect 458086 659912 458142 659968
rect 457994 657464 458050 657520
rect 457626 652840 457682 652896
rect 457534 650120 457590 650176
rect 457442 647672 457498 647728
rect 457350 623872 457406 623928
rect 457258 618296 457314 618352
rect 457902 643184 457958 643240
rect 457718 621016 457774 621072
rect 457810 615984 457866 616040
rect 459190 655696 459246 655752
rect 459006 645904 459062 645960
rect 458914 640328 458970 640384
rect 458822 611360 458878 611416
rect 458638 608640 458694 608696
rect 459098 628088 459154 628144
rect 459006 603608 459062 603664
rect 458914 599528 458970 599584
rect 458730 598168 458786 598224
rect 459466 637880 459522 637936
rect 459374 635432 459430 635488
rect 459282 633392 459338 633448
rect 459190 542952 459246 543008
rect 459282 519560 459338 519616
rect 459558 626252 459614 626308
rect 459466 520920 459522 520976
rect 459374 519424 459430 519480
rect 459834 614080 459890 614136
rect 459742 601840 459798 601896
rect 459926 606328 459982 606384
rect 467102 522280 467158 522336
rect 468574 521056 468630 521112
rect 491850 516180 491906 516216
rect 491850 516160 491852 516180
rect 491852 516160 491904 516180
rect 491904 516160 491906 516180
rect 494058 515888 494114 515944
rect 494058 513032 494114 513088
rect 487986 453872 488042 453928
rect 472162 391176 472218 391232
rect 472898 389000 472954 389056
rect 474370 389000 474426 389056
rect 475106 389000 475162 389056
rect 476578 389000 476634 389056
rect 479522 389000 479578 389056
rect 473634 388864 473690 388920
rect 494242 508816 494298 508872
rect 494150 505144 494206 505200
rect 494978 505164 495034 505200
rect 494978 505144 494980 505164
rect 494980 505144 495032 505164
rect 495032 505144 495034 505164
rect 494702 501200 494758 501256
rect 510710 364520 510766 364576
rect 509790 362480 509846 362536
rect 509330 360304 509386 360360
rect 451554 136484 451556 136504
rect 451556 136484 451608 136504
rect 451608 136484 451610 136504
rect 451554 136448 451610 136484
rect 452106 150320 452162 150376
rect 452382 157292 452384 157312
rect 452384 157292 452436 157312
rect 452436 157292 452438 157312
rect 452382 157256 452438 157292
rect 452382 155796 452384 155816
rect 452384 155796 452436 155816
rect 452436 155796 452438 155816
rect 452382 155760 452438 155796
rect 452382 154300 452384 154320
rect 452384 154300 452436 154320
rect 452436 154300 452438 154320
rect 452382 154264 452438 154300
rect 452566 158380 452568 158400
rect 452568 158380 452620 158400
rect 452620 158380 452622 158400
rect 452566 158344 452622 158380
rect 452474 153040 452530 153096
rect 452290 151680 452346 151736
rect 452566 148996 452568 149016
rect 452568 148996 452620 149016
rect 452620 148996 452622 149016
rect 452566 148960 452622 148996
rect 452566 147500 452568 147520
rect 452568 147500 452620 147520
rect 452620 147500 452622 147520
rect 452566 147464 452622 147500
rect 452566 146140 452568 146160
rect 452568 146140 452620 146160
rect 452620 146140 452622 146160
rect 452566 146104 452622 146140
rect 452566 144780 452568 144800
rect 452568 144780 452620 144800
rect 452620 144780 452622 144800
rect 452566 144744 452622 144780
rect 452566 143420 452568 143440
rect 452568 143420 452620 143440
rect 452620 143420 452622 143440
rect 452566 143384 452622 143420
rect 452566 142060 452568 142080
rect 452568 142060 452620 142080
rect 452620 142060 452622 142080
rect 452566 142024 452622 142060
rect 452566 140700 452568 140720
rect 452568 140700 452620 140720
rect 452620 140700 452622 140720
rect 452566 140664 452622 140700
rect 452566 139340 452568 139360
rect 452568 139340 452620 139360
rect 452620 139340 452622 139360
rect 452566 139304 452622 139340
rect 452566 137844 452568 137864
rect 452568 137844 452620 137864
rect 452620 137844 452622 137864
rect 452566 137808 452622 137844
rect 452566 135124 452568 135144
rect 452568 135124 452620 135144
rect 452620 135124 452622 135144
rect 452566 135088 452622 135124
rect 452566 133764 452568 133784
rect 452568 133764 452620 133784
rect 452620 133764 452622 133784
rect 452566 133728 452622 133764
rect 452566 132404 452568 132424
rect 452568 132404 452620 132424
rect 452620 132404 452622 132424
rect 452566 132368 452622 132404
rect 452566 131044 452568 131064
rect 452568 131044 452620 131064
rect 452620 131044 452622 131064
rect 452566 131008 452622 131044
rect 452566 129684 452568 129704
rect 452568 129684 452620 129704
rect 452620 129684 452622 129704
rect 452566 129648 452622 129684
rect 452290 128308 452346 128344
rect 452290 128288 452292 128308
rect 452292 128288 452344 128308
rect 452344 128288 452346 128308
rect 452382 126948 452438 126984
rect 452382 126928 452384 126948
rect 452384 126928 452436 126948
rect 452436 126928 452438 126948
rect 452198 126248 452254 126304
rect 452014 124888 452070 124944
rect 451922 123528 451978 123584
rect 451922 121488 451978 121544
rect 458270 321408 458326 321464
rect 460754 321136 460810 321192
rect 459926 321000 459982 321056
rect 459650 320864 459706 320920
rect 461306 320048 461362 320104
rect 456706 234912 456762 234968
rect 456706 207168 456762 207224
rect 456982 262656 457038 262712
rect 456890 234912 456946 234968
rect 458086 248784 458142 248840
rect 457902 221040 457958 221096
rect 459466 221040 459522 221096
rect 459374 207168 459430 207224
rect 470966 319776 471022 319832
rect 471242 319640 471298 319696
rect 479246 320048 479302 320104
rect 480902 321272 480958 321328
rect 480626 319912 480682 319968
rect 481454 319504 481510 319560
rect 500774 313928 500830 313984
rect 507122 321680 507178 321736
rect 507766 321816 507822 321872
rect 507306 320864 507362 320920
rect 507490 320728 507546 320784
rect 507674 321272 507730 321328
rect 509422 358808 509478 358864
rect 509514 357584 509570 357640
rect 509606 343984 509662 344040
rect 509698 334192 509754 334248
rect 509698 329296 509754 329352
rect 509606 303184 509662 303240
rect 509698 300192 509754 300248
rect 509974 331472 510030 331528
rect 509882 326576 509938 326632
rect 510158 324264 510214 324320
rect 510618 323176 510674 323232
rect 510158 306040 510214 306096
rect 510986 362344 511042 362400
rect 510894 356360 510950 356416
rect 511078 352552 511134 352608
rect 511170 346024 511226 346080
rect 512090 380296 512146 380352
rect 511998 378120 512054 378176
rect 512182 378664 512238 378720
rect 512734 384648 512790 384704
rect 513286 384104 513342 384160
rect 513010 383560 513066 383616
rect 512458 382492 512514 382528
rect 512458 382472 512460 382492
rect 512460 382472 512512 382492
rect 512512 382472 512514 382492
rect 512366 381928 512422 381984
rect 512274 377576 512330 377632
rect 512090 376488 512146 376544
rect 512458 375944 512514 376000
rect 512826 383036 512882 383072
rect 512826 383016 512828 383036
rect 512828 383016 512880 383036
rect 512880 383016 512882 383036
rect 513286 381384 513342 381440
rect 512826 380840 512882 380896
rect 513286 379752 513342 379808
rect 513286 379208 513342 379264
rect 513286 377032 513342 377088
rect 512734 375420 512790 375456
rect 512734 375400 512736 375420
rect 512736 375400 512788 375420
rect 512788 375400 512790 375420
rect 512550 374856 512606 374912
rect 513286 374312 513342 374368
rect 512642 373768 512698 373824
rect 512642 373224 512698 373280
rect 513286 372700 513342 372736
rect 513286 372680 513288 372700
rect 513288 372680 513340 372700
rect 513340 372680 513342 372700
rect 512090 372136 512146 372192
rect 512182 371592 512238 371648
rect 512090 371048 512146 371104
rect 512090 369960 512146 370016
rect 511998 367784 512054 367840
rect 511538 365608 511594 365664
rect 511446 347656 511502 347712
rect 511170 303048 511226 303104
rect 511998 363976 512054 364032
rect 511998 361276 512054 361312
rect 511998 361256 512000 361276
rect 512000 361256 512052 361276
rect 512052 361256 512054 361276
rect 511998 358536 512054 358592
rect 513286 370504 513342 370560
rect 512734 369416 512790 369472
rect 512274 368892 512330 368928
rect 512274 368872 512276 368892
rect 512276 368872 512328 368892
rect 512328 368872 512330 368892
rect 513286 368328 513342 368384
rect 513286 367240 513342 367296
rect 513010 366696 513066 366752
rect 513286 366152 513342 366208
rect 512366 365064 512422 365120
rect 512458 361800 512514 361856
rect 512274 355816 512330 355872
rect 513286 363432 513342 363488
rect 513286 360204 513288 360224
rect 513288 360204 513340 360224
rect 513340 360204 513342 360224
rect 513286 360168 513342 360204
rect 512642 359624 512698 359680
rect 513194 357992 513250 358048
rect 513286 356904 513342 356960
rect 513286 355272 513342 355328
rect 513286 354748 513342 354784
rect 513286 354728 513288 354748
rect 513288 354728 513340 354748
rect 513340 354728 513342 354748
rect 512458 354184 512514 354240
rect 512826 353640 512882 353696
rect 513010 353096 513066 353152
rect 512458 352028 512514 352064
rect 512458 352008 512460 352028
rect 512460 352008 512512 352028
rect 512512 352008 512514 352028
rect 513286 351464 513342 351520
rect 512458 350920 512514 350976
rect 512826 350376 512882 350432
rect 512458 349832 512514 349888
rect 512550 349288 512606 349344
rect 513286 348744 513342 348800
rect 513102 348200 513158 348256
rect 513194 347112 513250 347168
rect 512550 346568 512606 346624
rect 512458 343304 512514 343360
rect 512458 334600 512514 334656
rect 513102 341148 513158 341184
rect 513102 341128 513104 341148
rect 513104 341128 513156 341148
rect 513156 341128 513158 341148
rect 512642 340584 512698 340640
rect 513010 338952 513066 339008
rect 513010 337864 513066 337920
rect 513102 337320 513158 337376
rect 512826 335144 512882 335200
rect 512826 332424 512882 332480
rect 512734 328616 512790 328672
rect 512826 325352 512882 325408
rect 512734 305632 512790 305688
rect 512918 323176 512974 323232
rect 512642 302776 512698 302832
rect 513286 345480 513342 345536
rect 513286 344936 513342 344992
rect 513286 343868 513342 343904
rect 513286 343848 513288 343868
rect 513288 343848 513340 343868
rect 513340 343848 513342 343868
rect 513286 342252 513288 342272
rect 513288 342252 513340 342272
rect 513340 342252 513342 342272
rect 513286 342216 513342 342252
rect 513286 341672 513342 341728
rect 513286 340040 513342 340096
rect 513286 339516 513342 339552
rect 513286 339496 513288 339516
rect 513288 339496 513340 339516
rect 513340 339496 513342 339516
rect 513286 338408 513342 338464
rect 513286 336776 513342 336832
rect 513286 336232 513342 336288
rect 513286 335688 513342 335744
rect 513286 333512 513342 333568
rect 513286 331880 513342 331936
rect 559654 699760 559710 699816
rect 580262 697176 580318 697232
rect 579618 644000 579674 644056
rect 557538 442856 557594 442912
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 529294 261568 529350 261624
rect 531318 243616 531374 243672
rect 530122 226208 530178 226264
rect 529938 209208 529994 209264
rect 462318 67496 462374 67552
rect 462502 67532 462504 67552
rect 462504 67532 462556 67552
rect 462556 67532 462558 67552
rect 462502 67496 462558 67532
rect 539322 137672 539378 137728
rect 539322 135632 539378 135688
rect 539598 99184 539654 99240
rect 540334 133320 540390 133376
rect 540242 127200 540298 127256
rect 540150 125160 540206 125216
rect 540058 117272 540114 117328
rect 539966 112784 540022 112840
rect 539874 109112 539930 109168
rect 539782 100544 539838 100600
rect 539690 86808 539746 86864
rect 541162 110880 541218 110936
rect 541070 102720 541126 102776
rect 542450 121080 542506 121136
rect 541530 114960 541586 115016
rect 541438 106800 541494 106856
rect 541346 104760 541402 104816
rect 541254 88440 541310 88496
rect 542726 131280 542782 131336
rect 543094 123120 543150 123176
rect 543002 119040 543058 119096
rect 542910 96600 542966 96656
rect 543186 94560 543242 94616
rect 542818 92520 542874 92576
rect 542634 90480 542690 90536
rect 542542 84360 542598 84416
rect 540978 82320 541034 82376
rect 580170 590960 580226 591016
rect 579618 564304 579674 564360
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 578882 458088 578938 458144
rect 580170 431568 580226 431624
rect 579802 378392 579858 378448
rect 580170 365064 580226 365120
rect 580170 351872 580226 351928
rect 580354 683848 580410 683904
rect 580170 325216 580226 325272
rect 580446 670656 580502 670712
rect 580538 577632 580594 577688
rect 580630 537784 580686 537840
rect 580722 511264 580778 511320
rect 580814 418240 580870 418296
rect 580906 404912 580962 404968
rect 540610 48864 540666 48920
rect 536838 40976 536894 41032
rect 536838 33632 536894 33688
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 580262 258848 580318 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 579986 232328 580042 232384
rect 580170 219000 580226 219056
rect 579802 205672 579858 205728
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 578882 46280 578938 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
rect 384486 3304 384542 3360
<< metal3 >>
rect 235165 700634 235231 700637
rect 450486 700634 450492 700636
rect 235165 700632 450492 700634
rect 235165 700576 235170 700632
rect 235226 700576 450492 700632
rect 235165 700574 450492 700576
rect 235165 700571 235231 700574
rect 450486 700572 450492 700574
rect 450556 700572 450562 700636
rect 170305 700498 170371 700501
rect 444230 700498 444236 700500
rect 170305 700496 444236 700498
rect 170305 700440 170310 700496
rect 170366 700440 444236 700496
rect 170305 700438 444236 700440
rect 170305 700435 170371 700438
rect 444230 700436 444236 700438
rect 444300 700436 444306 700500
rect 137829 700362 137895 700365
rect 447726 700362 447732 700364
rect 137829 700360 447732 700362
rect 137829 700304 137834 700360
rect 137890 700304 447732 700360
rect 137829 700302 447732 700304
rect 137829 700299 137895 700302
rect 447726 700300 447732 700302
rect 447796 700300 447802 700364
rect 526294 699756 526300 699820
rect 526364 699818 526370 699820
rect 527173 699818 527239 699821
rect 526364 699816 527239 699818
rect 526364 699760 527178 699816
rect 527234 699760 527239 699816
rect 526364 699758 527239 699760
rect 526364 699756 526370 699758
rect 527173 699755 527239 699758
rect 559414 699756 559420 699820
rect 559484 699818 559490 699820
rect 559649 699818 559715 699821
rect 559484 699816 559715 699818
rect 559484 699760 559654 699816
rect 559710 699760 559715 699816
rect 559484 699758 559715 699760
rect 559484 699756 559490 699758
rect 559649 699755 559715 699758
rect -960 697220 480 697460
rect 580257 697234 580323 697237
rect 583520 697234 584960 697324
rect 580257 697232 584960 697234
rect 580257 697176 580262 697232
rect 580318 697176 584960 697232
rect 580257 697174 584960 697176
rect 580257 697171 580323 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3233 684314 3299 684317
rect -960 684312 3299 684314
rect -960 684256 3238 684312
rect 3294 684256 3299 684312
rect -960 684254 3299 684256
rect -960 684164 480 684254
rect 3233 684251 3299 684254
rect 201493 684042 201559 684045
rect 450670 684042 450676 684044
rect 201493 684040 450676 684042
rect 201493 683984 201498 684040
rect 201554 683984 450676 684040
rect 201493 683982 450676 683984
rect 201493 683979 201559 683982
rect 450670 683980 450676 683982
rect 450740 683980 450746 684044
rect 23473 683906 23539 683909
rect 446254 683906 446260 683908
rect 23473 683904 446260 683906
rect 23473 683848 23478 683904
rect 23534 683848 446260 683904
rect 23473 683846 446260 683848
rect 23473 683843 23539 683846
rect 446254 683844 446260 683846
rect 446324 683844 446330 683908
rect 580349 683906 580415 683909
rect 583520 683906 584960 683996
rect 580349 683904 584960 683906
rect 580349 683848 580354 683904
rect 580410 683848 584960 683904
rect 580349 683846 584960 683848
rect 580349 683843 580415 683846
rect 6913 683770 6979 683773
rect 446438 683770 446444 683772
rect 6913 683768 446444 683770
rect 6913 683712 6918 683768
rect 6974 683712 446444 683768
rect 6913 683710 446444 683712
rect 6913 683707 6979 683710
rect 446438 683708 446444 683710
rect 446508 683708 446514 683772
rect 583520 683756 584960 683846
rect 3550 683300 3556 683364
rect 3620 683362 3626 683364
rect 445293 683362 445359 683365
rect 3620 683360 445359 683362
rect 3620 683304 445298 683360
rect 445354 683304 445359 683360
rect 3620 683302 445359 683304
rect 3620 683300 3626 683302
rect 445293 683299 445359 683302
rect 3734 683164 3740 683228
rect 3804 683226 3810 683228
rect 446765 683226 446831 683229
rect 3804 683224 446831 683226
rect 3804 683168 446770 683224
rect 446826 683168 446831 683224
rect 3804 683166 446831 683168
rect 3804 683164 3810 683166
rect 446765 683163 446831 683166
rect 3366 682892 3372 682956
rect 3436 682954 3442 682956
rect 420269 682954 420335 682957
rect 3436 682952 420335 682954
rect 3436 682896 420274 682952
rect 420330 682896 420335 682952
rect 3436 682894 420335 682896
rect 3436 682892 3442 682894
rect 420269 682891 420335 682894
rect 3049 682818 3115 682821
rect 447910 682818 447916 682820
rect 3049 682816 447916 682818
rect 3049 682760 3054 682816
rect 3110 682760 447916 682816
rect 3049 682758 447916 682760
rect 3049 682755 3115 682758
rect 447910 682756 447916 682758
rect 447980 682756 447986 682820
rect 361757 679010 361823 679013
rect 359812 679008 361823 679010
rect 359812 678952 361762 679008
rect 361818 678952 361823 679008
rect 359812 678950 361823 678952
rect 361757 678947 361823 678950
rect -960 671258 480 671348
rect 3734 671258 3740 671260
rect -960 671198 3740 671258
rect -960 671108 480 671198
rect 3734 671196 3740 671198
rect 3804 671196 3810 671260
rect 580441 670714 580507 670717
rect 583520 670714 584960 670804
rect 580441 670712 584960 670714
rect 580441 670656 580446 670712
rect 580502 670656 584960 670712
rect 580441 670654 584960 670656
rect 580441 670651 580507 670654
rect 583520 670564 584960 670654
rect 361757 667994 361823 667997
rect 359812 667992 361823 667994
rect 359812 667936 361762 667992
rect 361818 667936 361823 667992
rect 359812 667934 361823 667936
rect 361757 667931 361823 667934
rect 459645 667994 459711 667997
rect 459645 667992 460092 667994
rect 459645 667936 459650 667992
rect 459706 667936 460092 667992
rect 459645 667934 460092 667936
rect 459645 667931 459711 667934
rect 458030 665212 458036 665276
rect 458100 665274 458106 665276
rect 460062 665274 460122 665448
rect 458100 665214 460122 665274
rect 458100 665212 458106 665214
rect 457846 662492 457852 662556
rect 457916 662554 457922 662556
rect 460062 662554 460122 663000
rect 457916 662494 460122 662554
rect 457916 662492 457922 662494
rect 458081 659970 458147 659973
rect 460062 659970 460122 660552
rect 458081 659968 460122 659970
rect 458081 659912 458086 659968
rect 458142 659912 460122 659968
rect 458081 659910 460122 659912
rect 458081 659907 458147 659910
rect -960 658202 480 658292
rect 3141 658202 3207 658205
rect -960 658200 3207 658202
rect -960 658144 3146 658200
rect 3202 658144 3207 658200
rect -960 658142 3207 658144
rect -960 658052 480 658142
rect 3141 658139 3207 658142
rect 457989 657522 458055 657525
rect 460062 657522 460122 658104
rect 457989 657520 460122 657522
rect 457989 657464 457994 657520
rect 458050 657464 460122 657520
rect 457989 657462 460122 657464
rect 457989 657459 458055 657462
rect 583520 657236 584960 657476
rect 361757 656978 361823 656981
rect 359812 656976 361823 656978
rect 359812 656920 361762 656976
rect 361818 656920 361823 656976
rect 359812 656918 361823 656920
rect 361757 656915 361823 656918
rect 459185 655754 459251 655757
rect 459185 655752 460092 655754
rect 459185 655696 459190 655752
rect 459246 655696 460092 655752
rect 459185 655694 460092 655696
rect 459185 655691 459251 655694
rect 457621 652898 457687 652901
rect 460062 652898 460122 653208
rect 457621 652896 460122 652898
rect 457621 652840 457626 652896
rect 457682 652840 460122 652896
rect 457621 652838 460122 652840
rect 457621 652835 457687 652838
rect 457529 650178 457595 650181
rect 460062 650178 460122 650760
rect 457529 650176 460122 650178
rect 457529 650120 457534 650176
rect 457590 650120 460122 650176
rect 457529 650118 460122 650120
rect 457529 650115 457595 650118
rect 457437 647730 457503 647733
rect 460062 647730 460122 648312
rect 457437 647728 460122 647730
rect 457437 647672 457442 647728
rect 457498 647672 460122 647728
rect 457437 647670 460122 647672
rect 457437 647667 457503 647670
rect 361757 645962 361823 645965
rect 359812 645960 361823 645962
rect 359812 645904 361762 645960
rect 361818 645904 361823 645960
rect 359812 645902 361823 645904
rect 361757 645899 361823 645902
rect 459001 645962 459067 645965
rect 459001 645960 460092 645962
rect 459001 645904 459006 645960
rect 459062 645904 460092 645960
rect 459001 645902 460092 645904
rect 459001 645899 459067 645902
rect -960 644996 480 645236
rect 579613 644058 579679 644061
rect 583520 644058 584960 644148
rect 579613 644056 584960 644058
rect 579613 644000 579618 644056
rect 579674 644000 584960 644056
rect 579613 643998 584960 644000
rect 579613 643995 579679 643998
rect 583520 643908 584960 643998
rect 457897 643242 457963 643245
rect 460062 643242 460122 643416
rect 457897 643240 460122 643242
rect 457897 643184 457902 643240
rect 457958 643184 460122 643240
rect 457897 643182 460122 643184
rect 457897 643179 457963 643182
rect 458909 640386 458975 640389
rect 460062 640386 460122 640968
rect 458909 640384 460122 640386
rect 458909 640328 458914 640384
rect 458970 640328 460122 640384
rect 458909 640326 460122 640328
rect 458909 640323 458975 640326
rect 459461 637938 459527 637941
rect 460062 637938 460122 638520
rect 459461 637936 460122 637938
rect 459461 637880 459466 637936
rect 459522 637880 460122 637936
rect 459461 637878 460122 637880
rect 459461 637875 459527 637878
rect 459369 635490 459435 635493
rect 460062 635490 460122 636072
rect 459369 635488 460122 635490
rect 459369 635432 459374 635488
rect 459430 635432 460122 635488
rect 459369 635430 460122 635432
rect 459369 635427 459435 635430
rect 361573 634946 361639 634949
rect 359812 634944 361639 634946
rect 359812 634888 361578 634944
rect 361634 634888 361639 634944
rect 359812 634886 361639 634888
rect 361573 634883 361639 634886
rect 459277 633450 459343 633453
rect 460062 633450 460122 633624
rect 459277 633448 460122 633450
rect 459277 633392 459282 633448
rect 459338 633392 460122 633448
rect 459277 633390 460122 633392
rect 459277 633387 459343 633390
rect -960 632090 480 632180
rect 3693 632090 3759 632093
rect -960 632088 3759 632090
rect -960 632032 3698 632088
rect 3754 632032 3759 632088
rect -960 632030 3759 632032
rect -960 631940 480 632030
rect 3693 632027 3759 632030
rect 459134 630668 459140 630732
rect 459204 630730 459210 630732
rect 460062 630730 460122 631176
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 459204 630670 460122 630730
rect 583520 630716 584960 630806
rect 459204 630668 459210 630670
rect 459093 628146 459159 628149
rect 460062 628146 460122 628728
rect 459093 628144 460122 628146
rect 459093 628088 459098 628144
rect 459154 628088 460122 628144
rect 459093 628086 460122 628088
rect 459093 628083 459159 628086
rect 459553 626310 459619 626313
rect 459553 626308 460092 626310
rect 459553 626252 459558 626308
rect 459614 626252 460092 626308
rect 459553 626250 460092 626252
rect 459553 626247 459619 626250
rect 361573 623930 361639 623933
rect 359812 623928 361639 623930
rect 359812 623872 361578 623928
rect 361634 623872 361639 623928
rect 359812 623870 361639 623872
rect 361573 623867 361639 623870
rect 457345 623930 457411 623933
rect 457345 623928 460092 623930
rect 457345 623872 457350 623928
rect 457406 623872 460092 623928
rect 457345 623870 460092 623872
rect 457345 623867 457411 623870
rect 457713 621074 457779 621077
rect 460062 621074 460122 621384
rect 457713 621072 460122 621074
rect 457713 621016 457718 621072
rect 457774 621016 460122 621072
rect 457713 621014 460122 621016
rect 457713 621011 457779 621014
rect -960 619170 480 619260
rect 3550 619170 3556 619172
rect -960 619110 3556 619170
rect -960 619020 480 619110
rect 3550 619108 3556 619110
rect 3620 619108 3626 619172
rect 457253 618354 457319 618357
rect 460062 618354 460122 618936
rect 457253 618352 460122 618354
rect 457253 618296 457258 618352
rect 457314 618296 460122 618352
rect 457253 618294 460122 618296
rect 457253 618291 457319 618294
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect 457805 616042 457871 616045
rect 460062 616042 460122 616488
rect 457805 616040 460122 616042
rect 457805 615984 457810 616040
rect 457866 615984 460122 616040
rect 457805 615982 460122 615984
rect 457805 615979 457871 615982
rect 459829 614138 459895 614141
rect 459829 614136 460092 614138
rect 459829 614080 459834 614136
rect 459890 614080 460092 614136
rect 459829 614078 460092 614080
rect 459829 614075 459895 614078
rect 361573 612914 361639 612917
rect 359812 612912 361639 612914
rect 359812 612856 361578 612912
rect 361634 612856 361639 612912
rect 359812 612854 361639 612856
rect 361573 612851 361639 612854
rect 458817 611418 458883 611421
rect 460062 611418 460122 611592
rect 458817 611416 460122 611418
rect 458817 611360 458822 611416
rect 458878 611360 460122 611416
rect 458817 611358 460122 611360
rect 458817 611355 458883 611358
rect 458633 608698 458699 608701
rect 460062 608698 460122 609144
rect 458633 608696 460122 608698
rect 458633 608640 458638 608696
rect 458694 608640 460122 608696
rect 458633 608638 460122 608640
rect 458633 608635 458699 608638
rect 459921 606386 459987 606389
rect 460062 606386 460122 606696
rect 459921 606384 460122 606386
rect 459921 606328 459926 606384
rect 459982 606328 460122 606384
rect 459921 606326 460122 606328
rect 459921 606323 459987 606326
rect -960 606114 480 606204
rect 3366 606114 3372 606116
rect -960 606054 3372 606114
rect -960 605964 480 606054
rect 3366 606052 3372 606054
rect 3436 606052 3442 606116
rect 459001 603666 459067 603669
rect 460062 603666 460122 604248
rect 583520 604060 584960 604300
rect 459001 603664 460122 603666
rect 459001 603608 459006 603664
rect 459062 603608 460122 603664
rect 459001 603606 460122 603608
rect 459001 603603 459067 603606
rect 361757 601898 361823 601901
rect 359812 601896 361823 601898
rect 359812 601840 361762 601896
rect 361818 601840 361823 601896
rect 359812 601838 361823 601840
rect 361757 601835 361823 601838
rect 459737 601898 459803 601901
rect 459737 601896 460092 601898
rect 459737 601840 459742 601896
rect 459798 601840 460092 601896
rect 459737 601838 460092 601840
rect 459737 601835 459803 601838
rect 458909 599586 458975 599589
rect 474774 599586 474780 599588
rect 458909 599584 474780 599586
rect 458909 599528 458914 599584
rect 458970 599528 474780 599584
rect 458909 599526 474780 599528
rect 458909 599523 458975 599526
rect 474774 599524 474780 599526
rect 474844 599524 474850 599588
rect 458725 598226 458791 598229
rect 476430 598226 476436 598228
rect 458725 598224 476436 598226
rect 458725 598168 458730 598224
rect 458786 598168 476436 598224
rect 458725 598166 476436 598168
rect 458725 598163 458791 598166
rect 476430 598164 476436 598166
rect 476500 598164 476506 598228
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 361757 590882 361823 590885
rect 359812 590880 361823 590882
rect 359812 590824 361762 590880
rect 361818 590824 361823 590880
rect 583520 590868 584960 590958
rect 359812 590822 361823 590824
rect 361757 590819 361823 590822
rect -960 580002 480 580092
rect 3233 580002 3299 580005
rect -960 580000 3299 580002
rect -960 579944 3238 580000
rect 3294 579944 3299 580000
rect -960 579942 3299 579944
rect -960 579852 480 579942
rect 3233 579939 3299 579942
rect 361757 579866 361823 579869
rect 359812 579864 361823 579866
rect 359812 579808 361762 579864
rect 361818 579808 361823 579864
rect 359812 579806 361823 579808
rect 361757 579803 361823 579806
rect 580533 577690 580599 577693
rect 583520 577690 584960 577780
rect 580533 577688 584960 577690
rect 580533 577632 580538 577688
rect 580594 577632 584960 577688
rect 580533 577630 584960 577632
rect 580533 577627 580599 577630
rect 583520 577540 584960 577630
rect 361757 568850 361823 568853
rect 359812 568848 361823 568850
rect 359812 568792 361762 568848
rect 361818 568792 361823 568848
rect 359812 568790 361823 568792
rect 361757 568787 361823 568790
rect -960 566946 480 567036
rect 3325 566946 3391 566949
rect -960 566944 3391 566946
rect -960 566888 3330 566944
rect 3386 566888 3391 566944
rect -960 566886 3391 566888
rect -960 566796 480 566886
rect 3325 566883 3391 566886
rect 579613 564362 579679 564365
rect 583520 564362 584960 564452
rect 579613 564360 584960 564362
rect 579613 564304 579618 564360
rect 579674 564304 584960 564360
rect 579613 564302 584960 564304
rect 579613 564299 579679 564302
rect 583520 564212 584960 564302
rect 361573 557834 361639 557837
rect 359812 557832 361639 557834
rect 359812 557776 361578 557832
rect 361634 557776 361639 557832
rect 359812 557774 361639 557776
rect 361573 557771 361639 557774
rect -960 553890 480 553980
rect 4061 553890 4127 553893
rect -960 553888 4127 553890
rect -960 553832 4066 553888
rect 4122 553832 4127 553888
rect -960 553830 4127 553832
rect -960 553740 480 553830
rect 4061 553827 4127 553830
rect 583520 551020 584960 551260
rect 361573 546818 361639 546821
rect 359812 546816 361639 546818
rect 359812 546760 361578 546816
rect 361634 546760 361639 546816
rect 359812 546758 361639 546760
rect 361573 546755 361639 546758
rect 459185 543010 459251 543013
rect 478822 543010 478828 543012
rect 459185 543008 478828 543010
rect 459185 542952 459190 543008
rect 459246 542952 478828 543008
rect 459185 542950 478828 542952
rect 459185 542947 459251 542950
rect 478822 542948 478828 542950
rect 478892 542948 478898 543012
rect -960 540684 480 540924
rect 580625 537842 580691 537845
rect 583520 537842 584960 537932
rect 580625 537840 584960 537842
rect 580625 537784 580630 537840
rect 580686 537784 584960 537840
rect 580625 537782 584960 537784
rect 580625 537779 580691 537782
rect 583520 537692 584960 537782
rect 361573 535802 361639 535805
rect 359812 535800 361639 535802
rect 359812 535744 361578 535800
rect 361634 535744 361639 535800
rect 359812 535742 361639 535744
rect 361573 535739 361639 535742
rect -960 527914 480 528004
rect 3969 527914 4035 527917
rect -960 527912 4035 527914
rect -960 527856 3974 527912
rect 4030 527856 4035 527912
rect -960 527854 4035 527856
rect -960 527764 480 527854
rect 3969 527851 4035 527854
rect 361757 524786 361823 524789
rect 359812 524784 361823 524786
rect 359812 524728 361762 524784
rect 361818 524728 361823 524784
rect 359812 524726 361823 524728
rect 361757 524723 361823 524726
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect 458030 522276 458036 522340
rect 458100 522338 458106 522340
rect 467097 522338 467163 522341
rect 458100 522336 467163 522338
rect 458100 522280 467102 522336
rect 467158 522280 467163 522336
rect 458100 522278 467163 522280
rect 458100 522276 458106 522278
rect 467097 522275 467163 522278
rect 457846 521052 457852 521116
rect 457916 521114 457922 521116
rect 468569 521114 468635 521117
rect 457916 521112 468635 521114
rect 457916 521056 468574 521112
rect 468630 521056 468635 521112
rect 457916 521054 468635 521056
rect 457916 521052 457922 521054
rect 468569 521051 468635 521054
rect 459461 520978 459527 520981
rect 474406 520978 474412 520980
rect 459461 520976 474412 520978
rect 459461 520920 459466 520976
rect 459522 520920 474412 520976
rect 459461 520918 474412 520920
rect 459461 520915 459527 520918
rect 474406 520916 474412 520918
rect 474476 520916 474482 520980
rect 459277 519618 459343 519621
rect 472014 519618 472020 519620
rect 459277 519616 472020 519618
rect 459277 519560 459282 519616
rect 459338 519560 472020 519616
rect 459277 519558 472020 519560
rect 459277 519555 459343 519558
rect 472014 519556 472020 519558
rect 472084 519556 472090 519620
rect 459369 519482 459435 519485
rect 474590 519482 474596 519484
rect 459369 519480 474596 519482
rect 459369 519424 459374 519480
rect 459430 519424 474596 519480
rect 459369 519422 474596 519424
rect 459369 519419 459435 519422
rect 474590 519420 474596 519422
rect 474660 519420 474666 519484
rect 447317 516218 447383 516221
rect 448513 516218 448579 516221
rect 450126 516218 450186 516528
rect 447317 516216 450186 516218
rect 447317 516160 447322 516216
rect 447378 516160 448518 516216
rect 448574 516160 450186 516216
rect 447317 516158 450186 516160
rect 491845 516218 491911 516221
rect 491845 516216 491954 516218
rect 491845 516160 491850 516216
rect 491906 516160 491954 516216
rect 447317 516155 447383 516158
rect 448513 516155 448579 516158
rect 491845 516155 491954 516160
rect 491894 515946 491954 516155
rect 494053 515946 494119 515949
rect 491894 515944 494119 515946
rect 491894 515888 494058 515944
rect 494114 515888 494119 515944
rect 491894 515886 494119 515888
rect 494053 515883 494119 515886
rect -960 514858 480 514948
rect 3877 514858 3943 514861
rect -960 514856 3943 514858
rect -960 514800 3882 514856
rect 3938 514800 3943 514856
rect -960 514798 3943 514800
rect -960 514708 480 514798
rect 3877 514795 3943 514798
rect 448329 514314 448395 514317
rect 450126 514314 450186 514352
rect 448329 514312 450186 514314
rect 448329 514256 448334 514312
rect 448390 514256 450186 514312
rect 448329 514254 450186 514256
rect 448329 514251 448395 514254
rect 361757 513770 361823 513773
rect 359812 513768 361823 513770
rect 359812 513712 361762 513768
rect 361818 513712 361823 513768
rect 359812 513710 361823 513712
rect 361757 513707 361823 513710
rect 494053 513090 494119 513093
rect 491894 513088 494119 513090
rect 491894 513032 494058 513088
rect 494114 513032 494119 513088
rect 491894 513030 494119 513032
rect 448237 512818 448303 512821
rect 448237 512816 450186 512818
rect 448237 512760 448242 512816
rect 448298 512760 450186 512816
rect 448237 512758 450186 512760
rect 448237 512755 448303 512758
rect 450126 512176 450186 512758
rect 491894 512448 491954 513030
rect 494053 513027 494119 513030
rect 580717 511322 580783 511325
rect 583520 511322 584960 511412
rect 580717 511320 584960 511322
rect 580717 511264 580722 511320
rect 580778 511264 584960 511320
rect 580717 511262 584960 511264
rect 580717 511259 580783 511262
rect 583520 511172 584960 511262
rect 448145 510506 448211 510509
rect 448421 510506 448487 510509
rect 448145 510504 450186 510506
rect 448145 510448 448150 510504
rect 448206 510448 448426 510504
rect 448482 510448 450186 510504
rect 448145 510446 450186 510448
rect 448145 510443 448211 510446
rect 448421 510443 448487 510446
rect 450126 510000 450186 510446
rect 491894 508874 491954 508912
rect 494237 508874 494303 508877
rect 491894 508872 494303 508874
rect 491894 508816 494242 508872
rect 494298 508816 494303 508872
rect 491894 508814 494303 508816
rect 494237 508811 494303 508814
rect 447685 507242 447751 507245
rect 450126 507242 450186 507824
rect 447685 507240 450186 507242
rect 447685 507184 447690 507240
rect 447746 507184 450186 507240
rect 447685 507182 450186 507184
rect 447685 507179 447751 507182
rect 448053 505202 448119 505205
rect 450126 505202 450186 505648
rect 448053 505200 450186 505202
rect 448053 505144 448058 505200
rect 448114 505144 450186 505200
rect 448053 505142 450186 505144
rect 491894 505202 491954 505376
rect 494145 505202 494211 505205
rect 494973 505202 495039 505205
rect 491894 505200 495039 505202
rect 491894 505144 494150 505200
rect 494206 505144 494978 505200
rect 495034 505144 495039 505200
rect 491894 505142 495039 505144
rect 448053 505139 448119 505142
rect 494145 505139 494211 505142
rect 494973 505139 495039 505142
rect 447869 503434 447935 503437
rect 449801 503434 449867 503437
rect 450126 503434 450186 503472
rect 447869 503432 450186 503434
rect 447869 503376 447874 503432
rect 447930 503376 449806 503432
rect 449862 503376 450186 503432
rect 447869 503374 450186 503376
rect 447869 503371 447935 503374
rect 449801 503371 449867 503374
rect 361757 502754 361823 502757
rect 359812 502752 361823 502754
rect 359812 502696 361762 502752
rect 361818 502696 361823 502752
rect 359812 502694 361823 502696
rect 361757 502691 361823 502694
rect 447961 501938 448027 501941
rect 447961 501936 450186 501938
rect -960 501802 480 501892
rect 447961 501880 447966 501936
rect 448022 501880 450186 501936
rect 447961 501878 450186 501880
rect 447961 501875 448027 501878
rect 3785 501802 3851 501805
rect -960 501800 3851 501802
rect -960 501744 3790 501800
rect 3846 501744 3851 501800
rect -960 501742 3851 501744
rect -960 501652 480 501742
rect 3785 501739 3851 501742
rect 450126 500986 450186 501878
rect 491894 501258 491954 501840
rect 494697 501258 494763 501261
rect 489870 501256 494763 501258
rect 489870 501200 494702 501256
rect 494758 501200 494763 501256
rect 489870 501198 494763 501200
rect 489870 501122 489930 501198
rect 494697 501195 494763 501198
rect 470550 501062 489930 501122
rect 470550 500986 470610 501062
rect 450126 500926 470610 500986
rect 583520 497844 584960 498084
rect 362217 491738 362283 491741
rect 359812 491736 362283 491738
rect 359812 491680 362222 491736
rect 362278 491680 362283 491736
rect 359812 491678 362283 491680
rect 362217 491675 362283 491678
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect 361757 480722 361823 480725
rect 359812 480720 361823 480722
rect 359812 480664 361762 480720
rect 361818 480664 361823 480720
rect 359812 480662 361823 480664
rect 361757 480659 361823 480662
rect -960 475690 480 475780
rect 3601 475690 3667 475693
rect -960 475688 3667 475690
rect -960 475632 3606 475688
rect 3662 475632 3667 475688
rect -960 475630 3667 475632
rect -960 475540 480 475630
rect 3601 475627 3667 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect 361757 469706 361823 469709
rect 359812 469704 361823 469706
rect 359812 469648 361762 469704
rect 361818 469648 361823 469704
rect 359812 469646 361823 469648
rect 361757 469643 361823 469646
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 361757 458690 361823 458693
rect 359812 458688 361823 458690
rect 359812 458632 361762 458688
rect 361818 458632 361823 458688
rect 359812 458630 361823 458632
rect 361757 458627 361823 458630
rect 578877 458146 578943 458149
rect 583520 458146 584960 458236
rect 578877 458144 584960 458146
rect 578877 458088 578882 458144
rect 578938 458088 584960 458144
rect 578877 458086 584960 458088
rect 578877 458083 578943 458086
rect 583520 457996 584960 458086
rect 487102 453868 487108 453932
rect 487172 453930 487178 453932
rect 487981 453930 488047 453933
rect 487172 453928 488047 453930
rect 487172 453872 487986 453928
rect 488042 453872 488047 453928
rect 487172 453870 488047 453872
rect 487172 453868 487178 453870
rect 487981 453867 488047 453870
rect -960 449578 480 449668
rect 3417 449578 3483 449581
rect -960 449576 3483 449578
rect -960 449520 3422 449576
rect 3478 449520 3483 449576
rect -960 449518 3483 449520
rect -960 449428 480 449518
rect 3417 449515 3483 449518
rect 362309 447674 362375 447677
rect 359812 447672 362375 447674
rect 359812 447616 362314 447672
rect 362370 447616 362375 447672
rect 359812 447614 362375 447616
rect 362309 447611 362375 447614
rect 583520 444668 584960 444908
rect 557533 442914 557599 442917
rect 555956 442912 557599 442914
rect 555956 442856 557538 442912
rect 557594 442856 557599 442912
rect 555956 442854 557599 442856
rect 557533 442851 557599 442854
rect -960 436508 480 436748
rect 361757 436658 361823 436661
rect 359812 436656 361823 436658
rect 359812 436600 361762 436656
rect 361818 436600 361823 436656
rect 359812 436598 361823 436600
rect 361757 436595 361823 436598
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect 362401 425642 362467 425645
rect 359812 425640 362467 425642
rect 359812 425584 362406 425640
rect 362462 425584 362467 425640
rect 359812 425582 362467 425584
rect 362401 425579 362467 425582
rect -960 423602 480 423692
rect 3693 423602 3759 423605
rect -960 423600 3759 423602
rect -960 423544 3698 423600
rect 3754 423544 3759 423600
rect -960 423542 3759 423544
rect -960 423452 480 423542
rect 3693 423539 3759 423542
rect 580809 418298 580875 418301
rect 583520 418298 584960 418388
rect 580809 418296 584960 418298
rect 580809 418240 580814 418296
rect 580870 418240 584960 418296
rect 580809 418238 584960 418240
rect 580809 418235 580875 418238
rect 583520 418148 584960 418238
rect 361573 414626 361639 414629
rect 359812 414624 361639 414626
rect 359812 414568 361578 414624
rect 361634 414568 361639 414624
rect 359812 414566 361639 414568
rect 361573 414563 361639 414566
rect -960 410546 480 410636
rect 3969 410546 4035 410549
rect -960 410544 4035 410546
rect -960 410488 3974 410544
rect 4030 410488 4035 410544
rect -960 410486 4035 410488
rect -960 410396 480 410486
rect 3969 410483 4035 410486
rect 580901 404970 580967 404973
rect 583520 404970 584960 405060
rect 580901 404968 584960 404970
rect 580901 404912 580906 404968
rect 580962 404912 584960 404968
rect 580901 404910 584960 404912
rect 580901 404907 580967 404910
rect 583520 404820 584960 404910
rect 361573 403610 361639 403613
rect 359812 403608 361639 403610
rect 359812 403552 361578 403608
rect 361634 403552 361639 403608
rect 359812 403550 361639 403552
rect 361573 403547 361639 403550
rect -960 397490 480 397580
rect 3877 397490 3943 397493
rect -960 397488 3943 397490
rect -960 397432 3882 397488
rect 3938 397432 3943 397488
rect -960 397430 3943 397432
rect -960 397340 480 397430
rect 3877 397427 3943 397430
rect 361573 392594 361639 392597
rect 359812 392592 361639 392594
rect 359812 392536 361578 392592
rect 361634 392536 361639 392592
rect 359812 392534 361639 392536
rect 361573 392531 361639 392534
rect 583520 391628 584960 391868
rect 459134 391172 459140 391236
rect 459204 391234 459210 391236
rect 472157 391234 472223 391237
rect 459204 391232 472223 391234
rect 459204 391176 472162 391232
rect 472218 391176 472223 391232
rect 459204 391174 472223 391176
rect 459204 391172 459210 391174
rect 472157 391171 472223 391174
rect 472014 388996 472020 389060
rect 472084 389058 472090 389060
rect 472893 389058 472959 389061
rect 474365 389060 474431 389061
rect 474365 389058 474412 389060
rect 472084 389056 472959 389058
rect 472084 389000 472898 389056
rect 472954 389000 472959 389056
rect 472084 388998 472959 389000
rect 474320 389056 474412 389058
rect 474320 389000 474370 389056
rect 474320 388998 474412 389000
rect 472084 388996 472090 388998
rect 472893 388995 472959 388998
rect 474365 388996 474412 388998
rect 474476 388996 474482 389060
rect 474774 388996 474780 389060
rect 474844 389058 474850 389060
rect 475101 389058 475167 389061
rect 474844 389056 475167 389058
rect 474844 389000 475106 389056
rect 475162 389000 475167 389056
rect 474844 388998 475167 389000
rect 474844 388996 474850 388998
rect 474365 388995 474431 388996
rect 475101 388995 475167 388998
rect 476430 388996 476436 389060
rect 476500 389058 476506 389060
rect 476573 389058 476639 389061
rect 476500 389056 476639 389058
rect 476500 389000 476578 389056
rect 476634 389000 476639 389056
rect 476500 388998 476639 389000
rect 476500 388996 476506 388998
rect 476573 388995 476639 388998
rect 478822 388996 478828 389060
rect 478892 389058 478898 389060
rect 479517 389058 479583 389061
rect 478892 389056 479583 389058
rect 478892 389000 479522 389056
rect 479578 389000 479583 389056
rect 478892 388998 479583 389000
rect 478892 388996 478898 388998
rect 479517 388995 479583 388998
rect 473629 388922 473695 388925
rect 474590 388922 474596 388924
rect 473629 388920 474596 388922
rect 473629 388864 473634 388920
rect 473690 388864 474596 388920
rect 473629 388862 474596 388864
rect 473629 388859 473695 388862
rect 474590 388860 474596 388862
rect 474660 388860 474666 388924
rect 449341 385658 449407 385661
rect 487102 385658 487108 385660
rect 449341 385656 487108 385658
rect 449341 385600 449346 385656
rect 449402 385600 487108 385656
rect 449341 385598 487108 385600
rect 449341 385595 449407 385598
rect 487102 385596 487108 385598
rect 487172 385596 487178 385660
rect 512729 384706 512795 384709
rect 509956 384704 512795 384706
rect 509956 384648 512734 384704
rect 512790 384648 512795 384704
rect 509956 384646 512795 384648
rect 512729 384643 512795 384646
rect -960 384284 480 384524
rect 513281 384162 513347 384165
rect 509956 384160 513347 384162
rect 509956 384104 513286 384160
rect 513342 384104 513347 384160
rect 509956 384102 513347 384104
rect 513281 384099 513347 384102
rect 447133 383890 447199 383893
rect 447133 383888 450156 383890
rect 447133 383832 447138 383888
rect 447194 383832 450156 383888
rect 447133 383830 450156 383832
rect 447133 383827 447199 383830
rect 513005 383618 513071 383621
rect 509956 383616 513071 383618
rect 509956 383560 513010 383616
rect 513066 383560 513071 383616
rect 509956 383558 513071 383560
rect 513005 383555 513071 383558
rect 447133 383210 447199 383213
rect 447133 383208 450156 383210
rect 447133 383152 447138 383208
rect 447194 383152 450156 383208
rect 447133 383150 450156 383152
rect 447133 383147 447199 383150
rect 512821 383074 512887 383077
rect 509956 383072 512887 383074
rect 509956 383016 512826 383072
rect 512882 383016 512887 383072
rect 509956 383014 512887 383016
rect 512821 383011 512887 383014
rect 447225 382530 447291 382533
rect 512453 382530 512519 382533
rect 447225 382528 450156 382530
rect 447225 382472 447230 382528
rect 447286 382472 450156 382528
rect 447225 382470 450156 382472
rect 509956 382528 512519 382530
rect 509956 382472 512458 382528
rect 512514 382472 512519 382528
rect 509956 382470 512519 382472
rect 447225 382467 447291 382470
rect 512453 382467 512519 382470
rect 512361 381986 512427 381989
rect 509956 381984 512427 381986
rect 509956 381928 512366 381984
rect 512422 381928 512427 381984
rect 509956 381926 512427 381928
rect 512361 381923 512427 381926
rect 447133 381850 447199 381853
rect 447133 381848 450156 381850
rect 447133 381792 447138 381848
rect 447194 381792 450156 381848
rect 447133 381790 450156 381792
rect 447133 381787 447199 381790
rect 361573 381578 361639 381581
rect 359812 381576 361639 381578
rect 359812 381520 361578 381576
rect 361634 381520 361639 381576
rect 359812 381518 361639 381520
rect 361573 381515 361639 381518
rect 513281 381442 513347 381445
rect 509956 381440 513347 381442
rect 509956 381384 513286 381440
rect 513342 381384 513347 381440
rect 509956 381382 513347 381384
rect 513281 381379 513347 381382
rect 447225 381170 447291 381173
rect 447225 381168 450156 381170
rect 447225 381112 447230 381168
rect 447286 381112 450156 381168
rect 447225 381110 450156 381112
rect 447225 381107 447291 381110
rect 512821 380898 512887 380901
rect 509956 380896 512887 380898
rect 509956 380840 512826 380896
rect 512882 380840 512887 380896
rect 509956 380838 512887 380840
rect 512821 380835 512887 380838
rect 447133 380490 447199 380493
rect 447133 380488 450156 380490
rect 447133 380432 447138 380488
rect 447194 380432 450156 380488
rect 447133 380430 450156 380432
rect 447133 380427 447199 380430
rect 512085 380354 512151 380357
rect 509956 380352 512151 380354
rect 509956 380296 512090 380352
rect 512146 380296 512151 380352
rect 509956 380294 512151 380296
rect 512085 380291 512151 380294
rect 447225 379810 447291 379813
rect 513281 379810 513347 379813
rect 447225 379808 450156 379810
rect 447225 379752 447230 379808
rect 447286 379752 450156 379808
rect 447225 379750 450156 379752
rect 509956 379808 513347 379810
rect 509956 379752 513286 379808
rect 513342 379752 513347 379808
rect 509956 379750 513347 379752
rect 447225 379747 447291 379750
rect 513281 379747 513347 379750
rect 513281 379266 513347 379269
rect 509956 379264 513347 379266
rect 509956 379208 513286 379264
rect 513342 379208 513347 379264
rect 509956 379206 513347 379208
rect 513281 379203 513347 379206
rect 447133 379130 447199 379133
rect 447133 379128 450156 379130
rect 447133 379072 447138 379128
rect 447194 379072 450156 379128
rect 447133 379070 450156 379072
rect 447133 379067 447199 379070
rect 512177 378722 512243 378725
rect 509956 378720 512243 378722
rect 509956 378664 512182 378720
rect 512238 378664 512243 378720
rect 509956 378662 512243 378664
rect 512177 378659 512243 378662
rect 447225 378450 447291 378453
rect 579797 378450 579863 378453
rect 583520 378450 584960 378540
rect 447225 378448 450156 378450
rect 447225 378392 447230 378448
rect 447286 378392 450156 378448
rect 447225 378390 450156 378392
rect 579797 378448 584960 378450
rect 579797 378392 579802 378448
rect 579858 378392 584960 378448
rect 579797 378390 584960 378392
rect 447225 378387 447291 378390
rect 579797 378387 579863 378390
rect 583520 378300 584960 378390
rect 511993 378178 512059 378181
rect 509956 378176 512059 378178
rect 509956 378120 511998 378176
rect 512054 378120 512059 378176
rect 509956 378118 512059 378120
rect 511993 378115 512059 378118
rect 447133 377770 447199 377773
rect 447133 377768 450156 377770
rect 447133 377712 447138 377768
rect 447194 377712 450156 377768
rect 447133 377710 450156 377712
rect 447133 377707 447199 377710
rect 512269 377634 512335 377637
rect 509956 377632 512335 377634
rect 509956 377576 512274 377632
rect 512330 377576 512335 377632
rect 509956 377574 512335 377576
rect 512269 377571 512335 377574
rect 447225 377090 447291 377093
rect 513281 377090 513347 377093
rect 447225 377088 450156 377090
rect 447225 377032 447230 377088
rect 447286 377032 450156 377088
rect 447225 377030 450156 377032
rect 509956 377088 513347 377090
rect 509956 377032 513286 377088
rect 513342 377032 513347 377088
rect 509956 377030 513347 377032
rect 447225 377027 447291 377030
rect 513281 377027 513347 377030
rect 512085 376546 512151 376549
rect 509956 376544 512151 376546
rect 509956 376488 512090 376544
rect 512146 376488 512151 376544
rect 509956 376486 512151 376488
rect 512085 376483 512151 376486
rect 447133 376410 447199 376413
rect 447133 376408 450156 376410
rect 447133 376352 447138 376408
rect 447194 376352 450156 376408
rect 447133 376350 450156 376352
rect 447133 376347 447199 376350
rect 512453 376002 512519 376005
rect 509956 376000 512519 376002
rect 509956 375944 512458 376000
rect 512514 375944 512519 376000
rect 509956 375942 512519 375944
rect 512453 375939 512519 375942
rect 447225 375730 447291 375733
rect 447225 375728 450156 375730
rect 447225 375672 447230 375728
rect 447286 375672 450156 375728
rect 447225 375670 450156 375672
rect 447225 375667 447291 375670
rect 512729 375458 512795 375461
rect 509956 375456 512795 375458
rect 509956 375400 512734 375456
rect 512790 375400 512795 375456
rect 509956 375398 512795 375400
rect 512729 375395 512795 375398
rect 447133 375050 447199 375053
rect 447133 375048 450156 375050
rect 447133 374992 447138 375048
rect 447194 374992 450156 375048
rect 447133 374990 450156 374992
rect 447133 374987 447199 374990
rect 512545 374914 512611 374917
rect 509956 374912 512611 374914
rect 509956 374856 512550 374912
rect 512606 374856 512611 374912
rect 509956 374854 512611 374856
rect 512545 374851 512611 374854
rect 447225 374370 447291 374373
rect 513281 374370 513347 374373
rect 447225 374368 450156 374370
rect 447225 374312 447230 374368
rect 447286 374312 450156 374368
rect 447225 374310 450156 374312
rect 509956 374368 513347 374370
rect 509956 374312 513286 374368
rect 513342 374312 513347 374368
rect 509956 374310 513347 374312
rect 447225 374307 447291 374310
rect 513281 374307 513347 374310
rect 512637 373826 512703 373829
rect 509956 373824 512703 373826
rect 509956 373768 512642 373824
rect 512698 373768 512703 373824
rect 509956 373766 512703 373768
rect 512637 373763 512703 373766
rect 447133 373690 447199 373693
rect 447133 373688 450156 373690
rect 447133 373632 447138 373688
rect 447194 373632 450156 373688
rect 447133 373630 450156 373632
rect 447133 373627 447199 373630
rect 512637 373282 512703 373285
rect 509956 373280 512703 373282
rect 509956 373224 512642 373280
rect 512698 373224 512703 373280
rect 509956 373222 512703 373224
rect 512637 373219 512703 373222
rect 447225 373010 447291 373013
rect 447225 373008 450156 373010
rect 447225 372952 447230 373008
rect 447286 372952 450156 373008
rect 447225 372950 450156 372952
rect 447225 372947 447291 372950
rect 513281 372738 513347 372741
rect 509956 372736 513347 372738
rect 509956 372680 513286 372736
rect 513342 372680 513347 372736
rect 509956 372678 513347 372680
rect 513281 372675 513347 372678
rect 447133 372330 447199 372333
rect 447133 372328 450156 372330
rect 447133 372272 447138 372328
rect 447194 372272 450156 372328
rect 447133 372270 450156 372272
rect 447133 372267 447199 372270
rect 512085 372194 512151 372197
rect 509956 372192 512151 372194
rect 509956 372136 512090 372192
rect 512146 372136 512151 372192
rect 509956 372134 512151 372136
rect 512085 372131 512151 372134
rect 447225 371650 447291 371653
rect 512177 371650 512243 371653
rect 447225 371648 450156 371650
rect 447225 371592 447230 371648
rect 447286 371592 450156 371648
rect 447225 371590 450156 371592
rect 509956 371648 512243 371650
rect 509956 371592 512182 371648
rect 512238 371592 512243 371648
rect 509956 371590 512243 371592
rect 447225 371587 447291 371590
rect 512177 371587 512243 371590
rect -960 371378 480 371468
rect 3969 371378 4035 371381
rect -960 371376 4035 371378
rect -960 371320 3974 371376
rect 4030 371320 4035 371376
rect -960 371318 4035 371320
rect -960 371228 480 371318
rect 3969 371315 4035 371318
rect 512085 371106 512151 371109
rect 509956 371104 512151 371106
rect 509956 371048 512090 371104
rect 512146 371048 512151 371104
rect 509956 371046 512151 371048
rect 512085 371043 512151 371046
rect 447133 370970 447199 370973
rect 447133 370968 450156 370970
rect 447133 370912 447138 370968
rect 447194 370912 450156 370968
rect 447133 370910 450156 370912
rect 447133 370907 447199 370910
rect 361573 370562 361639 370565
rect 513281 370562 513347 370565
rect 359812 370560 361639 370562
rect 359812 370504 361578 370560
rect 361634 370504 361639 370560
rect 359812 370502 361639 370504
rect 509956 370560 513347 370562
rect 509956 370504 513286 370560
rect 513342 370504 513347 370560
rect 509956 370502 513347 370504
rect 361573 370499 361639 370502
rect 513281 370499 513347 370502
rect 447225 370290 447291 370293
rect 447225 370288 450156 370290
rect 447225 370232 447230 370288
rect 447286 370232 450156 370288
rect 447225 370230 450156 370232
rect 447225 370227 447291 370230
rect 512085 370018 512151 370021
rect 509956 370016 512151 370018
rect 509956 369960 512090 370016
rect 512146 369960 512151 370016
rect 509956 369958 512151 369960
rect 512085 369955 512151 369958
rect 447133 369610 447199 369613
rect 447133 369608 450156 369610
rect 447133 369552 447138 369608
rect 447194 369552 450156 369608
rect 447133 369550 450156 369552
rect 447133 369547 447199 369550
rect 512729 369474 512795 369477
rect 509956 369472 512795 369474
rect 509956 369416 512734 369472
rect 512790 369416 512795 369472
rect 509956 369414 512795 369416
rect 512729 369411 512795 369414
rect 447225 368930 447291 368933
rect 512269 368930 512335 368933
rect 447225 368928 450156 368930
rect 447225 368872 447230 368928
rect 447286 368872 450156 368928
rect 447225 368870 450156 368872
rect 509956 368928 512335 368930
rect 509956 368872 512274 368928
rect 512330 368872 512335 368928
rect 509956 368870 512335 368872
rect 447225 368867 447291 368870
rect 512269 368867 512335 368870
rect 513281 368386 513347 368389
rect 509956 368384 513347 368386
rect 509956 368328 513286 368384
rect 513342 368328 513347 368384
rect 509956 368326 513347 368328
rect 513281 368323 513347 368326
rect 447133 368250 447199 368253
rect 447133 368248 450156 368250
rect 447133 368192 447138 368248
rect 447194 368192 450156 368248
rect 447133 368190 450156 368192
rect 447133 368187 447199 368190
rect 511993 367842 512059 367845
rect 509956 367840 512059 367842
rect 509956 367784 511998 367840
rect 512054 367784 512059 367840
rect 509956 367782 512059 367784
rect 511993 367779 512059 367782
rect 447225 367570 447291 367573
rect 447225 367568 450156 367570
rect 447225 367512 447230 367568
rect 447286 367512 450156 367568
rect 447225 367510 450156 367512
rect 447225 367507 447291 367510
rect 513281 367298 513347 367301
rect 509956 367296 513347 367298
rect 509956 367240 513286 367296
rect 513342 367240 513347 367296
rect 509956 367238 513347 367240
rect 513281 367235 513347 367238
rect 447225 366890 447291 366893
rect 447225 366888 450156 366890
rect 447225 366832 447230 366888
rect 447286 366832 450156 366888
rect 447225 366830 450156 366832
rect 447225 366827 447291 366830
rect 513005 366754 513071 366757
rect 509956 366752 513071 366754
rect 509956 366696 513010 366752
rect 513066 366696 513071 366752
rect 509956 366694 513071 366696
rect 513005 366691 513071 366694
rect 447133 366210 447199 366213
rect 513281 366210 513347 366213
rect 447133 366208 450156 366210
rect 447133 366152 447138 366208
rect 447194 366152 450156 366208
rect 447133 366150 450156 366152
rect 509956 366208 513347 366210
rect 509956 366152 513286 366208
rect 513342 366152 513347 366208
rect 509956 366150 513347 366152
rect 447133 366147 447199 366150
rect 513281 366147 513347 366150
rect 511533 365666 511599 365669
rect 509956 365664 511599 365666
rect 509956 365608 511538 365664
rect 511594 365608 511599 365664
rect 509956 365606 511599 365608
rect 511533 365603 511599 365606
rect 447225 365530 447291 365533
rect 447225 365528 450156 365530
rect 447225 365472 447230 365528
rect 447286 365472 450156 365528
rect 447225 365470 450156 365472
rect 447225 365467 447291 365470
rect 512361 365122 512427 365125
rect 509956 365120 512427 365122
rect 509956 365064 512366 365120
rect 512422 365064 512427 365120
rect 509956 365062 512427 365064
rect 512361 365059 512427 365062
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect 447133 364850 447199 364853
rect 447133 364848 450156 364850
rect 447133 364792 447138 364848
rect 447194 364792 450156 364848
rect 447133 364790 450156 364792
rect 447133 364787 447199 364790
rect 510705 364578 510771 364581
rect 509956 364576 510771 364578
rect 509956 364520 510710 364576
rect 510766 364520 510771 364576
rect 509956 364518 510771 364520
rect 510705 364515 510771 364518
rect 447225 364170 447291 364173
rect 447225 364168 450156 364170
rect 447225 364112 447230 364168
rect 447286 364112 450156 364168
rect 447225 364110 450156 364112
rect 447225 364107 447291 364110
rect 511993 364034 512059 364037
rect 509956 364032 512059 364034
rect 509956 363976 511998 364032
rect 512054 363976 512059 364032
rect 509956 363974 512059 363976
rect 511993 363971 512059 363974
rect 447133 363490 447199 363493
rect 513281 363490 513347 363493
rect 447133 363488 450156 363490
rect 447133 363432 447138 363488
rect 447194 363432 450156 363488
rect 447133 363430 450156 363432
rect 509956 363488 513347 363490
rect 509956 363432 513286 363488
rect 513342 363432 513347 363488
rect 509956 363430 513347 363432
rect 447133 363427 447199 363430
rect 513281 363427 513347 363430
rect 447225 362810 447291 362813
rect 447225 362808 450156 362810
rect 447225 362752 447230 362808
rect 447286 362752 450156 362808
rect 447225 362750 450156 362752
rect 447225 362747 447291 362750
rect 509742 362541 509802 362916
rect 509742 362536 509851 362541
rect 509742 362480 509790 362536
rect 509846 362480 509851 362536
rect 509742 362478 509851 362480
rect 509785 362475 509851 362478
rect 510981 362402 511047 362405
rect 509956 362400 511047 362402
rect 509956 362344 510986 362400
rect 511042 362344 511047 362400
rect 509956 362342 511047 362344
rect 510981 362339 511047 362342
rect 447133 362130 447199 362133
rect 447133 362128 450156 362130
rect 447133 362072 447138 362128
rect 447194 362072 450156 362128
rect 447133 362070 450156 362072
rect 447133 362067 447199 362070
rect 512453 361858 512519 361861
rect 509956 361856 512519 361858
rect 509956 361800 512458 361856
rect 512514 361800 512519 361856
rect 509956 361798 512519 361800
rect 512453 361795 512519 361798
rect 447225 361450 447291 361453
rect 447225 361448 450156 361450
rect 447225 361392 447230 361448
rect 447286 361392 450156 361448
rect 447225 361390 450156 361392
rect 447225 361387 447291 361390
rect 511993 361314 512059 361317
rect 509956 361312 512059 361314
rect 509956 361256 511998 361312
rect 512054 361256 512059 361312
rect 509956 361254 512059 361256
rect 511993 361251 512059 361254
rect 447133 360770 447199 360773
rect 447133 360768 450156 360770
rect 447133 360712 447138 360768
rect 447194 360712 450156 360768
rect 447133 360710 450156 360712
rect 447133 360707 447199 360710
rect 509374 360365 509434 360740
rect 509325 360360 509434 360365
rect 509325 360304 509330 360360
rect 509386 360304 509434 360360
rect 509325 360302 509434 360304
rect 509325 360299 509391 360302
rect 513281 360226 513347 360229
rect 509956 360224 513347 360226
rect 509956 360168 513286 360224
rect 513342 360168 513347 360224
rect 509956 360166 513347 360168
rect 513281 360163 513347 360166
rect 447225 360090 447291 360093
rect 447225 360088 450156 360090
rect 447225 360032 447230 360088
rect 447286 360032 450156 360088
rect 447225 360030 450156 360032
rect 447225 360027 447291 360030
rect 512637 359682 512703 359685
rect 509956 359680 512703 359682
rect 509956 359624 512642 359680
rect 512698 359624 512703 359680
rect 509956 359622 512703 359624
rect 512637 359619 512703 359622
rect 362309 359546 362375 359549
rect 359812 359544 362375 359546
rect 359812 359488 362314 359544
rect 362370 359488 362375 359544
rect 359812 359486 362375 359488
rect 362309 359483 362375 359486
rect 447133 359410 447199 359413
rect 447133 359408 450156 359410
rect 447133 359352 447138 359408
rect 447194 359352 450156 359408
rect 447133 359350 450156 359352
rect 447133 359347 447199 359350
rect 509374 358869 509434 359108
rect 450445 358866 450511 358869
rect 450445 358864 450554 358866
rect 450445 358808 450450 358864
rect 450506 358808 450554 358864
rect 450445 358803 450554 358808
rect 509374 358864 509483 358869
rect 509374 358808 509422 358864
rect 509478 358808 509483 358864
rect 509374 358806 509483 358808
rect 509417 358803 509483 358806
rect 450494 358700 450554 358803
rect 511993 358594 512059 358597
rect 509956 358592 512059 358594
rect -960 358458 480 358548
rect 509956 358536 511998 358592
rect 512054 358536 512059 358592
rect 509956 358534 512059 358536
rect 511993 358531 512059 358534
rect 3417 358458 3483 358461
rect -960 358456 3483 358458
rect -960 358400 3422 358456
rect 3478 358400 3483 358456
rect -960 358398 3483 358400
rect -960 358308 480 358398
rect 3417 358395 3483 358398
rect 448973 358050 449039 358053
rect 513189 358050 513255 358053
rect 448973 358048 450156 358050
rect 448973 357992 448978 358048
rect 449034 357992 450156 358048
rect 448973 357990 450156 357992
rect 509956 358048 513255 358050
rect 509956 357992 513194 358048
rect 513250 357992 513255 358048
rect 509956 357990 513255 357992
rect 448973 357987 449039 357990
rect 513189 357987 513255 357990
rect 509509 357642 509575 357645
rect 509509 357640 509618 357642
rect 509509 357584 509514 357640
rect 509570 357584 509618 357640
rect 509509 357579 509618 357584
rect 509558 357476 509618 357579
rect 448421 357370 448487 357373
rect 448421 357368 450156 357370
rect 448421 357312 448426 357368
rect 448482 357312 450156 357368
rect 448421 357310 450156 357312
rect 448421 357307 448487 357310
rect 513281 356962 513347 356965
rect 509956 356960 513347 356962
rect 509956 356904 513286 356960
rect 513342 356904 513347 356960
rect 509956 356902 513347 356904
rect 513281 356899 513347 356902
rect 449433 356690 449499 356693
rect 449433 356688 450156 356690
rect 449433 356632 449438 356688
rect 449494 356632 450156 356688
rect 449433 356630 450156 356632
rect 449433 356627 449499 356630
rect 510889 356418 510955 356421
rect 509956 356416 510955 356418
rect 509956 356360 510894 356416
rect 510950 356360 510955 356416
rect 509956 356358 510955 356360
rect 510889 356355 510955 356358
rect 449801 356010 449867 356013
rect 449801 356008 450156 356010
rect 449801 355952 449806 356008
rect 449862 355952 450156 356008
rect 449801 355950 450156 355952
rect 449801 355947 449867 355950
rect 512269 355874 512335 355877
rect 509956 355872 512335 355874
rect 509956 355816 512274 355872
rect 512330 355816 512335 355872
rect 509956 355814 512335 355816
rect 512269 355811 512335 355814
rect 449525 355330 449591 355333
rect 513281 355330 513347 355333
rect 449525 355328 450156 355330
rect 449525 355272 449530 355328
rect 449586 355272 450156 355328
rect 449525 355270 450156 355272
rect 509956 355328 513347 355330
rect 509956 355272 513286 355328
rect 513342 355272 513347 355328
rect 509956 355270 513347 355272
rect 449525 355267 449591 355270
rect 513281 355267 513347 355270
rect 513281 354786 513347 354789
rect 509956 354784 513347 354786
rect 509956 354728 513286 354784
rect 513342 354728 513347 354784
rect 509956 354726 513347 354728
rect 513281 354723 513347 354726
rect 449617 354650 449683 354653
rect 449617 354648 450156 354650
rect 449617 354592 449622 354648
rect 449678 354592 450156 354648
rect 449617 354590 450156 354592
rect 449617 354587 449683 354590
rect 512453 354242 512519 354245
rect 509956 354240 512519 354242
rect 509956 354184 512458 354240
rect 512514 354184 512519 354240
rect 509956 354182 512519 354184
rect 512453 354179 512519 354182
rect 449709 353970 449775 353973
rect 449709 353968 450156 353970
rect 449709 353912 449714 353968
rect 449770 353912 450156 353968
rect 449709 353910 450156 353912
rect 449709 353907 449775 353910
rect 512821 353698 512887 353701
rect 509956 353696 512887 353698
rect 509956 353640 512826 353696
rect 512882 353640 512887 353696
rect 509956 353638 512887 353640
rect 512821 353635 512887 353638
rect 447685 353290 447751 353293
rect 447685 353288 450156 353290
rect 447685 353232 447690 353288
rect 447746 353232 450156 353288
rect 447685 353230 450156 353232
rect 447685 353227 447751 353230
rect 513005 353154 513071 353157
rect 509956 353152 513071 353154
rect 509956 353096 513010 353152
rect 513066 353096 513071 353152
rect 509956 353094 513071 353096
rect 513005 353091 513071 353094
rect 450261 353018 450327 353021
rect 450261 353016 450370 353018
rect 450261 352960 450266 353016
rect 450322 352960 450370 353016
rect 450261 352955 450370 352960
rect 450310 352580 450370 352955
rect 511073 352610 511139 352613
rect 509956 352608 511139 352610
rect 509956 352552 511078 352608
rect 511134 352552 511139 352608
rect 509956 352550 511139 352552
rect 511073 352547 511139 352550
rect 512453 352066 512519 352069
rect 509956 352064 512519 352066
rect 509956 352008 512458 352064
rect 512514 352008 512519 352064
rect 509956 352006 512519 352008
rect 512453 352003 512519 352006
rect 447133 351930 447199 351933
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 447133 351928 450156 351930
rect 447133 351872 447138 351928
rect 447194 351872 450156 351928
rect 447133 351870 450156 351872
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 447133 351867 447199 351870
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect 513281 351522 513347 351525
rect 509956 351520 513347 351522
rect 509956 351464 513286 351520
rect 513342 351464 513347 351520
rect 509956 351462 513347 351464
rect 513281 351459 513347 351462
rect 448421 351250 448487 351253
rect 448421 351248 450156 351250
rect 448421 351192 448426 351248
rect 448482 351192 450156 351248
rect 448421 351190 450156 351192
rect 448421 351187 448487 351190
rect 512453 350978 512519 350981
rect 509956 350976 512519 350978
rect 509956 350920 512458 350976
rect 512514 350920 512519 350976
rect 509956 350918 512519 350920
rect 512453 350915 512519 350918
rect 447133 350570 447199 350573
rect 447133 350568 450156 350570
rect 447133 350512 447138 350568
rect 447194 350512 450156 350568
rect 447133 350510 450156 350512
rect 447133 350507 447199 350510
rect 512821 350434 512887 350437
rect 509956 350432 512887 350434
rect 509956 350376 512826 350432
rect 512882 350376 512887 350432
rect 509956 350374 512887 350376
rect 512821 350371 512887 350374
rect 449617 349890 449683 349893
rect 512453 349890 512519 349893
rect 449617 349888 450156 349890
rect 449617 349832 449622 349888
rect 449678 349832 450156 349888
rect 449617 349830 450156 349832
rect 509956 349888 512519 349890
rect 509956 349832 512458 349888
rect 512514 349832 512519 349888
rect 509956 349830 512519 349832
rect 449617 349827 449683 349830
rect 512453 349827 512519 349830
rect 512545 349346 512611 349349
rect 509956 349344 512611 349346
rect 509956 349288 512550 349344
rect 512606 349288 512611 349344
rect 509956 349286 512611 349288
rect 512545 349283 512611 349286
rect 447777 349210 447843 349213
rect 447777 349208 450156 349210
rect 447777 349152 447782 349208
rect 447838 349152 450156 349208
rect 447777 349150 450156 349152
rect 447777 349147 447843 349150
rect 450169 348938 450235 348941
rect 450126 348936 450235 348938
rect 450126 348880 450174 348936
rect 450230 348880 450235 348936
rect 450126 348875 450235 348880
rect 361757 348530 361823 348533
rect 359812 348528 361823 348530
rect 359812 348472 361762 348528
rect 361818 348472 361823 348528
rect 450126 348500 450186 348875
rect 513281 348802 513347 348805
rect 509956 348800 513347 348802
rect 509956 348744 513286 348800
rect 513342 348744 513347 348800
rect 509956 348742 513347 348744
rect 513281 348739 513347 348742
rect 359812 348470 361823 348472
rect 361757 348467 361823 348470
rect 450353 348258 450419 348261
rect 513097 348258 513163 348261
rect 450310 348256 450419 348258
rect 450310 348200 450358 348256
rect 450414 348200 450419 348256
rect 450310 348195 450419 348200
rect 509956 348256 513163 348258
rect 509956 348200 513102 348256
rect 513158 348200 513163 348256
rect 509956 348198 513163 348200
rect 513097 348195 513163 348198
rect 450310 347820 450370 348195
rect 511441 347714 511507 347717
rect 509956 347712 511507 347714
rect 509956 347656 511446 347712
rect 511502 347656 511507 347712
rect 509956 347654 511507 347656
rect 511441 347651 511507 347654
rect 447133 347170 447199 347173
rect 513189 347170 513255 347173
rect 447133 347168 450156 347170
rect 447133 347112 447138 347168
rect 447194 347112 450156 347168
rect 447133 347110 450156 347112
rect 509956 347168 513255 347170
rect 509956 347112 513194 347168
rect 513250 347112 513255 347168
rect 509956 347110 513255 347112
rect 447133 347107 447199 347110
rect 513189 347107 513255 347110
rect 449985 346898 450051 346901
rect 449985 346896 450186 346898
rect 449985 346840 449990 346896
rect 450046 346840 450186 346896
rect 449985 346838 450186 346840
rect 449985 346835 450051 346838
rect 450126 346460 450186 346838
rect 512545 346626 512611 346629
rect 509956 346624 512611 346626
rect 509956 346568 512550 346624
rect 512606 346568 512611 346624
rect 509956 346566 512611 346568
rect 512545 346563 512611 346566
rect 449893 346218 449959 346221
rect 449893 346216 450186 346218
rect 449893 346160 449898 346216
rect 449954 346160 450186 346216
rect 449893 346158 450186 346160
rect 449893 346155 449959 346158
rect 450126 345780 450186 346158
rect 511165 346082 511231 346085
rect 509956 346080 511231 346082
rect 509956 346024 511170 346080
rect 511226 346024 511231 346080
rect 509956 346022 511231 346024
rect 511165 346019 511231 346022
rect 513281 345538 513347 345541
rect 509956 345536 513347 345538
rect -960 345402 480 345492
rect 509956 345480 513286 345536
rect 513342 345480 513347 345536
rect 509956 345478 513347 345480
rect 513281 345475 513347 345478
rect 3509 345402 3575 345405
rect -960 345400 3575 345402
rect -960 345344 3514 345400
rect 3570 345344 3575 345400
rect -960 345342 3575 345344
rect -960 345252 480 345342
rect 3509 345339 3575 345342
rect 449801 345130 449867 345133
rect 449801 345128 450156 345130
rect 449801 345072 449806 345128
rect 449862 345072 450156 345128
rect 449801 345070 450156 345072
rect 449801 345067 449867 345070
rect 513281 344994 513347 344997
rect 509956 344992 513347 344994
rect 509956 344936 513286 344992
rect 513342 344936 513347 344992
rect 509956 344934 513347 344936
rect 513281 344931 513347 344934
rect 447777 344450 447843 344453
rect 447777 344448 450156 344450
rect 447777 344392 447782 344448
rect 447838 344392 450156 344448
rect 447777 344390 450156 344392
rect 447777 344387 447843 344390
rect 509558 344045 509618 344420
rect 509558 344040 509667 344045
rect 509558 343984 509606 344040
rect 509662 343984 509667 344040
rect 509558 343982 509667 343984
rect 509601 343979 509667 343982
rect 513281 343906 513347 343909
rect 509956 343904 513347 343906
rect 509956 343848 513286 343904
rect 513342 343848 513347 343904
rect 509956 343846 513347 343848
rect 513281 343843 513347 343846
rect 447317 343770 447383 343773
rect 447317 343768 450156 343770
rect 447317 343712 447322 343768
rect 447378 343712 450156 343768
rect 447317 343710 450156 343712
rect 447317 343707 447383 343710
rect 512453 343362 512519 343365
rect 509956 343360 512519 343362
rect 509956 343304 512458 343360
rect 512514 343304 512519 343360
rect 509956 343302 512519 343304
rect 512453 343299 512519 343302
rect 449709 343090 449775 343093
rect 449709 343088 450156 343090
rect 449709 343032 449714 343088
rect 449770 343032 450156 343088
rect 449709 343030 450156 343032
rect 449709 343027 449775 343030
rect 510654 342818 510660 342820
rect 509956 342758 510660 342818
rect 510654 342756 510660 342758
rect 510724 342756 510730 342820
rect 449065 342410 449131 342413
rect 449065 342408 450156 342410
rect 449065 342352 449070 342408
rect 449126 342352 450156 342408
rect 449065 342350 450156 342352
rect 449065 342347 449131 342350
rect 513281 342274 513347 342277
rect 509956 342272 513347 342274
rect 509956 342216 513286 342272
rect 513342 342216 513347 342272
rect 509956 342214 513347 342216
rect 513281 342211 513347 342214
rect 447133 341730 447199 341733
rect 513281 341730 513347 341733
rect 447133 341728 450156 341730
rect 447133 341672 447138 341728
rect 447194 341672 450156 341728
rect 447133 341670 450156 341672
rect 509956 341728 513347 341730
rect 509956 341672 513286 341728
rect 513342 341672 513347 341728
rect 509956 341670 513347 341672
rect 447133 341667 447199 341670
rect 513281 341667 513347 341670
rect 513097 341186 513163 341189
rect 509956 341184 513163 341186
rect 509956 341128 513102 341184
rect 513158 341128 513163 341184
rect 509956 341126 513163 341128
rect 513097 341123 513163 341126
rect 447225 341050 447291 341053
rect 447225 341048 450156 341050
rect 447225 340992 447230 341048
rect 447286 340992 450156 341048
rect 447225 340990 450156 340992
rect 447225 340987 447291 340990
rect 512637 340642 512703 340645
rect 509956 340640 512703 340642
rect 509956 340584 512642 340640
rect 512698 340584 512703 340640
rect 509956 340582 512703 340584
rect 512637 340579 512703 340582
rect 447133 340370 447199 340373
rect 447133 340368 450156 340370
rect 447133 340312 447138 340368
rect 447194 340312 450156 340368
rect 447133 340310 450156 340312
rect 447133 340307 447199 340310
rect 513281 340098 513347 340101
rect 509956 340096 513347 340098
rect 509956 340040 513286 340096
rect 513342 340040 513347 340096
rect 509956 340038 513347 340040
rect 513281 340035 513347 340038
rect 447225 339690 447291 339693
rect 447225 339688 450156 339690
rect 447225 339632 447230 339688
rect 447286 339632 450156 339688
rect 447225 339630 450156 339632
rect 447225 339627 447291 339630
rect 513281 339554 513347 339557
rect 509956 339552 513347 339554
rect 509956 339496 513286 339552
rect 513342 339496 513347 339552
rect 509956 339494 513347 339496
rect 513281 339491 513347 339494
rect 447225 339010 447291 339013
rect 513005 339010 513071 339013
rect 447225 339008 450156 339010
rect 447225 338952 447230 339008
rect 447286 338952 450156 339008
rect 447225 338950 450156 338952
rect 509956 339008 513071 339010
rect 509956 338952 513010 339008
rect 513066 338952 513071 339008
rect 509956 338950 513071 338952
rect 447225 338947 447291 338950
rect 513005 338947 513071 338950
rect 513281 338466 513347 338469
rect 509956 338464 513347 338466
rect 509956 338408 513286 338464
rect 513342 338408 513347 338464
rect 583520 338452 584960 338692
rect 509956 338406 513347 338408
rect 513281 338403 513347 338406
rect 447133 338330 447199 338333
rect 447133 338328 450156 338330
rect 447133 338272 447138 338328
rect 447194 338272 450156 338328
rect 447133 338270 450156 338272
rect 447133 338267 447199 338270
rect 513005 337922 513071 337925
rect 509956 337920 513071 337922
rect 509956 337864 513010 337920
rect 513066 337864 513071 337920
rect 509956 337862 513071 337864
rect 513005 337859 513071 337862
rect 447225 337650 447291 337653
rect 447225 337648 450156 337650
rect 447225 337592 447230 337648
rect 447286 337592 450156 337648
rect 447225 337590 450156 337592
rect 447225 337587 447291 337590
rect 361757 337514 361823 337517
rect 359812 337512 361823 337514
rect 359812 337456 361762 337512
rect 361818 337456 361823 337512
rect 359812 337454 361823 337456
rect 361757 337451 361823 337454
rect 513097 337378 513163 337381
rect 509956 337376 513163 337378
rect 509956 337320 513102 337376
rect 513158 337320 513163 337376
rect 509956 337318 513163 337320
rect 513097 337315 513163 337318
rect 447133 336970 447199 336973
rect 447133 336968 450156 336970
rect 447133 336912 447138 336968
rect 447194 336912 450156 336968
rect 447133 336910 450156 336912
rect 447133 336907 447199 336910
rect 513281 336834 513347 336837
rect 509956 336832 513347 336834
rect 509956 336776 513286 336832
rect 513342 336776 513347 336832
rect 509956 336774 513347 336776
rect 513281 336771 513347 336774
rect 447225 336290 447291 336293
rect 513281 336290 513347 336293
rect 447225 336288 450156 336290
rect 447225 336232 447230 336288
rect 447286 336232 450156 336288
rect 447225 336230 450156 336232
rect 509956 336288 513347 336290
rect 509956 336232 513286 336288
rect 513342 336232 513347 336288
rect 509956 336230 513347 336232
rect 447225 336227 447291 336230
rect 513281 336227 513347 336230
rect 513281 335746 513347 335749
rect 509956 335744 513347 335746
rect 509956 335688 513286 335744
rect 513342 335688 513347 335744
rect 509956 335686 513347 335688
rect 513281 335683 513347 335686
rect 447317 335610 447383 335613
rect 447317 335608 450156 335610
rect 447317 335552 447322 335608
rect 447378 335552 450156 335608
rect 447317 335550 450156 335552
rect 447317 335547 447383 335550
rect 512821 335202 512887 335205
rect 509956 335200 512887 335202
rect 509956 335144 512826 335200
rect 512882 335144 512887 335200
rect 509956 335142 512887 335144
rect 512821 335139 512887 335142
rect 447317 334930 447383 334933
rect 447317 334928 450156 334930
rect 447317 334872 447322 334928
rect 447378 334872 450156 334928
rect 447317 334870 450156 334872
rect 447317 334867 447383 334870
rect 420729 334794 420795 334797
rect 442441 334794 442507 334797
rect 420729 334792 442507 334794
rect 420729 334736 420734 334792
rect 420790 334736 442446 334792
rect 442502 334736 442507 334792
rect 420729 334734 442507 334736
rect 420729 334731 420795 334734
rect 442441 334731 442507 334734
rect 420085 334658 420151 334661
rect 450537 334658 450603 334661
rect 512453 334658 512519 334661
rect 420085 334656 450603 334658
rect 420085 334600 420090 334656
rect 420146 334600 450542 334656
rect 450598 334600 450603 334656
rect 420085 334598 450603 334600
rect 509956 334656 512519 334658
rect 509956 334600 512458 334656
rect 512514 334600 512519 334656
rect 509956 334598 512519 334600
rect 420085 334595 420151 334598
rect 450537 334595 450603 334598
rect 512453 334595 512519 334598
rect 420729 334522 420795 334525
rect 421046 334522 421052 334524
rect 420729 334520 421052 334522
rect 420729 334464 420734 334520
rect 420790 334464 421052 334520
rect 420729 334462 421052 334464
rect 420729 334459 420795 334462
rect 421046 334460 421052 334462
rect 421116 334460 421122 334524
rect 428089 334522 428155 334525
rect 428406 334522 428412 334524
rect 428089 334520 428412 334522
rect 428089 334464 428094 334520
rect 428150 334464 428412 334520
rect 428089 334462 428412 334464
rect 428089 334459 428155 334462
rect 428406 334460 428412 334462
rect 428476 334460 428482 334524
rect 447225 334250 447291 334253
rect 509693 334250 509759 334253
rect 447225 334248 450156 334250
rect 447225 334192 447230 334248
rect 447286 334192 450156 334248
rect 447225 334190 450156 334192
rect 509693 334248 509802 334250
rect 509693 334192 509698 334248
rect 509754 334192 509802 334248
rect 447225 334187 447291 334190
rect 509693 334187 509802 334192
rect 509742 334084 509802 334187
rect 447317 333570 447383 333573
rect 513281 333570 513347 333573
rect 447317 333568 450156 333570
rect 447317 333512 447322 333568
rect 447378 333512 450156 333568
rect 447317 333510 450156 333512
rect 509956 333568 513347 333570
rect 509956 333512 513286 333568
rect 513342 333512 513347 333568
rect 509956 333510 513347 333512
rect 447317 333507 447383 333510
rect 513281 333507 513347 333510
rect 514886 333026 514892 333028
rect 509956 332966 514892 333026
rect 514886 332964 514892 332966
rect 514956 332964 514962 333028
rect 432597 332890 432663 332893
rect 429916 332888 432663 332890
rect 429916 332832 432602 332888
rect 432658 332832 432663 332888
rect 429916 332830 432663 332832
rect 432597 332827 432663 332830
rect 447225 332890 447291 332893
rect 447225 332888 450156 332890
rect 447225 332832 447230 332888
rect 447286 332832 450156 332888
rect 447225 332830 450156 332832
rect 447225 332827 447291 332830
rect 512821 332482 512887 332485
rect 509956 332480 512887 332482
rect -960 332196 480 332436
rect 509956 332424 512826 332480
rect 512882 332424 512887 332480
rect 509956 332422 512887 332424
rect 512821 332419 512887 332422
rect 447593 332210 447659 332213
rect 447593 332208 450156 332210
rect 447593 332152 447598 332208
rect 447654 332180 450156 332208
rect 447654 332152 450186 332180
rect 447593 332150 450186 332152
rect 447593 332147 447659 332150
rect 449985 331666 450051 331669
rect 450126 331666 450186 332150
rect 513281 331938 513347 331941
rect 509956 331936 513347 331938
rect 509956 331880 513286 331936
rect 513342 331880 513347 331936
rect 509956 331878 513347 331880
rect 513281 331875 513347 331878
rect 449985 331664 450186 331666
rect 449985 331608 449990 331664
rect 450046 331608 450186 331664
rect 449985 331606 450186 331608
rect 449985 331603 450051 331606
rect 447225 331530 447291 331533
rect 509969 331530 510035 331533
rect 447225 331528 450156 331530
rect 447225 331472 447230 331528
rect 447286 331472 450156 331528
rect 447225 331470 450156 331472
rect 509926 331528 510035 331530
rect 509926 331472 509974 331528
rect 510030 331472 510035 331528
rect 447225 331467 447291 331470
rect 509926 331467 510035 331472
rect 509926 331364 509986 331467
rect 447225 330850 447291 330853
rect 514334 330850 514340 330852
rect 447225 330848 450156 330850
rect 447225 330792 447230 330848
rect 447286 330792 450156 330848
rect 447225 330790 450156 330792
rect 509956 330790 514340 330850
rect 447225 330787 447291 330790
rect 514334 330788 514340 330790
rect 514404 330788 514410 330852
rect 514702 330306 514708 330308
rect 509956 330246 514708 330306
rect 514702 330244 514708 330246
rect 514772 330244 514778 330308
rect 447225 330170 447291 330173
rect 447225 330168 450156 330170
rect 447225 330112 447230 330168
rect 447286 330112 450156 330168
rect 447225 330110 450156 330112
rect 447225 330107 447291 330110
rect 447225 329490 447291 329493
rect 447225 329488 450156 329490
rect 447225 329432 447230 329488
rect 447286 329432 450156 329488
rect 447225 329430 450156 329432
rect 447225 329427 447291 329430
rect 509742 329357 509802 329732
rect 509693 329352 509802 329357
rect 509693 329296 509698 329352
rect 509754 329296 509802 329352
rect 509693 329294 509802 329296
rect 509693 329291 509759 329294
rect 432413 329218 432479 329221
rect 517830 329218 517836 329220
rect 429916 329216 432479 329218
rect 429916 329160 432418 329216
rect 432474 329160 432479 329216
rect 429916 329158 432479 329160
rect 509956 329158 517836 329218
rect 432413 329155 432479 329158
rect 517830 329156 517836 329158
rect 517900 329156 517906 329220
rect 447225 328810 447291 328813
rect 447225 328808 450156 328810
rect 447225 328752 447230 328808
rect 447286 328752 450156 328808
rect 447225 328750 450156 328752
rect 447225 328747 447291 328750
rect 512729 328674 512795 328677
rect 509956 328672 512795 328674
rect 509956 328616 512734 328672
rect 512790 328616 512795 328672
rect 509956 328614 512795 328616
rect 512729 328611 512795 328614
rect 447225 328130 447291 328133
rect 448329 328130 448395 328133
rect 514150 328130 514156 328132
rect 447225 328128 450156 328130
rect 447225 328072 447230 328128
rect 447286 328072 448334 328128
rect 448390 328072 450156 328128
rect 447225 328070 450156 328072
rect 509956 328070 514156 328130
rect 447225 328067 447291 328070
rect 448329 328067 448395 328070
rect 514150 328068 514156 328070
rect 514220 328068 514226 328132
rect 510838 327586 510844 327588
rect 509956 327526 510844 327586
rect 510838 327524 510844 327526
rect 510908 327524 510914 327588
rect 448237 327450 448303 327453
rect 448237 327448 450156 327450
rect 448237 327392 448242 327448
rect 448298 327392 450156 327448
rect 448237 327390 450156 327392
rect 448237 327387 448303 327390
rect 448145 326770 448211 326773
rect 448145 326768 450156 326770
rect 448145 326712 448150 326768
rect 448206 326712 450156 326768
rect 448145 326710 450156 326712
rect 448145 326707 448211 326710
rect 509926 326637 509986 327012
rect 509877 326632 509986 326637
rect 509877 326576 509882 326632
rect 509938 326576 509986 326632
rect 509877 326574 509986 326576
rect 509877 326571 509943 326574
rect 362217 326498 362283 326501
rect 511206 326498 511212 326500
rect 359812 326496 362283 326498
rect 359812 326440 362222 326496
rect 362278 326440 362283 326496
rect 359812 326438 362283 326440
rect 509956 326438 511212 326498
rect 362217 326435 362283 326438
rect 511206 326436 511212 326438
rect 511276 326436 511282 326500
rect 447225 326090 447291 326093
rect 447225 326088 450156 326090
rect 447225 326032 447230 326088
rect 447286 326032 450156 326088
rect 447225 326030 450156 326032
rect 447225 326027 447291 326030
rect 511022 325954 511028 325956
rect 509956 325894 511028 325954
rect 511022 325892 511028 325894
rect 511092 325892 511098 325956
rect 432689 325546 432755 325549
rect 429916 325544 432755 325546
rect 429916 325488 432694 325544
rect 432750 325488 432755 325544
rect 429916 325486 432755 325488
rect 432689 325483 432755 325486
rect 448053 325410 448119 325413
rect 512821 325410 512887 325413
rect 448053 325408 450156 325410
rect 448053 325352 448058 325408
rect 448114 325352 450156 325408
rect 448053 325350 450156 325352
rect 509956 325408 512887 325410
rect 509956 325352 512826 325408
rect 512882 325352 512887 325408
rect 509956 325350 512887 325352
rect 448053 325347 448119 325350
rect 512821 325347 512887 325350
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 510286 324866 510292 324868
rect 509956 324806 510292 324866
rect 510286 324804 510292 324806
rect 510356 324804 510362 324868
rect 447961 324730 448027 324733
rect 448237 324730 448303 324733
rect 447961 324728 450156 324730
rect 447961 324672 447966 324728
rect 448022 324672 448242 324728
rect 448298 324672 450156 324728
rect 447961 324670 450156 324672
rect 447961 324667 448027 324670
rect 448237 324667 448303 324670
rect 510153 324322 510219 324325
rect 509956 324320 510219 324322
rect 509956 324264 510158 324320
rect 510214 324264 510219 324320
rect 509956 324262 510219 324264
rect 510153 324259 510219 324262
rect 447317 324050 447383 324053
rect 448329 324050 448395 324053
rect 449341 324050 449407 324053
rect 447317 324048 450156 324050
rect 447317 323992 447322 324048
rect 447378 323992 448334 324048
rect 448390 323992 449346 324048
rect 449402 323992 450156 324048
rect 447317 323990 450156 323992
rect 447317 323987 447383 323990
rect 448329 323987 448395 323990
rect 449341 323987 449407 323990
rect 510470 323778 510476 323780
rect 509956 323718 510476 323778
rect 510470 323716 510476 323718
rect 510540 323716 510546 323780
rect 510613 323234 510679 323237
rect 512913 323234 512979 323237
rect 509956 323232 512979 323234
rect 509956 323176 510618 323232
rect 510674 323176 512918 323232
rect 512974 323176 512979 323232
rect 509956 323174 512979 323176
rect 510613 323171 510679 323174
rect 512913 323171 512979 323174
rect 432873 321874 432939 321877
rect 429916 321872 432939 321874
rect 429916 321816 432878 321872
rect 432934 321816 432939 321872
rect 429916 321814 432939 321816
rect 432873 321811 432939 321814
rect 507761 321874 507827 321877
rect 510286 321874 510292 321876
rect 507761 321872 510292 321874
rect 507761 321816 507766 321872
rect 507822 321816 510292 321872
rect 507761 321814 510292 321816
rect 507761 321811 507827 321814
rect 510286 321812 510292 321814
rect 510356 321812 510362 321876
rect 507117 321738 507183 321741
rect 511022 321738 511028 321740
rect 507117 321736 511028 321738
rect 507117 321680 507122 321736
rect 507178 321680 511028 321736
rect 507117 321678 511028 321680
rect 507117 321675 507183 321678
rect 511022 321676 511028 321678
rect 511092 321676 511098 321740
rect 458265 321466 458331 321469
rect 559414 321466 559420 321468
rect 458265 321464 559420 321466
rect 458265 321408 458270 321464
rect 458326 321408 559420 321464
rect 458265 321406 559420 321408
rect 458265 321403 458331 321406
rect 559414 321404 559420 321406
rect 559484 321404 559490 321468
rect 447726 321268 447732 321332
rect 447796 321330 447802 321332
rect 480897 321330 480963 321333
rect 447796 321328 480963 321330
rect 447796 321272 480902 321328
rect 480958 321272 480963 321328
rect 447796 321270 480963 321272
rect 447796 321268 447802 321270
rect 480897 321267 480963 321270
rect 507669 321330 507735 321333
rect 510838 321330 510844 321332
rect 507669 321328 510844 321330
rect 507669 321272 507674 321328
rect 507730 321272 510844 321328
rect 507669 321270 510844 321272
rect 507669 321267 507735 321270
rect 510838 321268 510844 321270
rect 510908 321268 510914 321332
rect 445477 321194 445543 321197
rect 460749 321194 460815 321197
rect 445477 321192 460815 321194
rect 445477 321136 445482 321192
rect 445538 321136 460754 321192
rect 460810 321136 460815 321192
rect 445477 321134 460815 321136
rect 445477 321131 445543 321134
rect 460749 321131 460815 321134
rect 444230 320996 444236 321060
rect 444300 321058 444306 321060
rect 459921 321058 459987 321061
rect 444300 321056 459987 321058
rect 444300 321000 459926 321056
rect 459982 321000 459987 321056
rect 444300 320998 459987 321000
rect 444300 320996 444306 320998
rect 459921 320995 459987 320998
rect 450486 320860 450492 320924
rect 450556 320922 450562 320924
rect 459645 320922 459711 320925
rect 450556 320920 459711 320922
rect 450556 320864 459650 320920
rect 459706 320864 459711 320920
rect 450556 320862 459711 320864
rect 450556 320860 450562 320862
rect 459645 320859 459711 320862
rect 507301 320922 507367 320925
rect 514334 320922 514340 320924
rect 507301 320920 514340 320922
rect 507301 320864 507306 320920
rect 507362 320864 514340 320920
rect 507301 320862 514340 320864
rect 507301 320859 507367 320862
rect 514334 320860 514340 320862
rect 514404 320860 514410 320924
rect 507485 320786 507551 320789
rect 517830 320786 517836 320788
rect 507485 320784 517836 320786
rect 507485 320728 507490 320784
rect 507546 320728 517836 320784
rect 507485 320726 517836 320728
rect 507485 320723 507551 320726
rect 517830 320724 517836 320726
rect 517900 320724 517906 320788
rect 447910 320044 447916 320108
rect 447980 320106 447986 320108
rect 461301 320106 461367 320109
rect 447980 320104 461367 320106
rect 447980 320048 461306 320104
rect 461362 320048 461367 320104
rect 447980 320046 461367 320048
rect 447980 320044 447986 320046
rect 461301 320043 461367 320046
rect 479241 320106 479307 320109
rect 526294 320106 526300 320108
rect 479241 320104 526300 320106
rect 479241 320048 479246 320104
rect 479302 320048 526300 320104
rect 479241 320046 526300 320048
rect 479241 320043 479307 320046
rect 526294 320044 526300 320046
rect 526364 320044 526370 320108
rect 450670 319908 450676 319972
rect 450740 319970 450746 319972
rect 480621 319970 480687 319973
rect 450740 319968 480687 319970
rect 450740 319912 480626 319968
rect 480682 319912 480687 319968
rect 450740 319910 480687 319912
rect 450740 319908 450746 319910
rect 480621 319907 480687 319910
rect 446254 319772 446260 319836
rect 446324 319834 446330 319836
rect 470961 319834 471027 319837
rect 446324 319832 471027 319834
rect 446324 319776 470966 319832
rect 471022 319776 471027 319832
rect 446324 319774 471027 319776
rect 446324 319772 446330 319774
rect 470961 319771 471027 319774
rect 446765 319698 446831 319701
rect 471237 319698 471303 319701
rect 446765 319696 471303 319698
rect 446765 319640 446770 319696
rect 446826 319640 471242 319696
rect 471298 319640 471303 319696
rect 446765 319638 471303 319640
rect 446765 319635 446831 319638
rect 471237 319635 471303 319638
rect 446438 319500 446444 319564
rect 446508 319562 446514 319564
rect 481449 319562 481515 319565
rect 446508 319560 481515 319562
rect 446508 319504 481454 319560
rect 481510 319504 481515 319560
rect 446508 319502 481515 319504
rect 446508 319500 446514 319502
rect 481449 319499 481515 319502
rect -960 319290 480 319380
rect 3785 319290 3851 319293
rect -960 319288 3851 319290
rect -960 319232 3790 319288
rect 3846 319232 3851 319288
rect -960 319230 3851 319232
rect -960 319140 480 319230
rect 3785 319227 3851 319230
rect 432781 318202 432847 318205
rect 429916 318200 432847 318202
rect 429916 318144 432786 318200
rect 432842 318144 432847 318200
rect 429916 318142 432847 318144
rect 432781 318139 432847 318142
rect 361757 315482 361823 315485
rect 359812 315480 361823 315482
rect 359812 315424 361762 315480
rect 361818 315424 361823 315480
rect 359812 315422 361823 315424
rect 361757 315419 361823 315422
rect 433241 314530 433307 314533
rect 429916 314528 433307 314530
rect 429916 314472 433246 314528
rect 433302 314472 433307 314528
rect 429916 314470 433307 314472
rect 433241 314467 433307 314470
rect 500769 313986 500835 313989
rect 538254 313986 538260 313988
rect 500769 313984 538260 313986
rect 500769 313928 500774 313984
rect 500830 313928 538260 313984
rect 500769 313926 538260 313928
rect 500769 313923 500835 313926
rect 538254 313924 538260 313926
rect 538324 313924 538330 313988
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect 432597 310858 432663 310861
rect 429916 310856 432663 310858
rect 429916 310800 432602 310856
rect 432658 310800 432663 310856
rect 429916 310798 432663 310800
rect 432597 310795 432663 310798
rect 432229 307186 432295 307189
rect 429916 307184 432295 307186
rect 429916 307128 432234 307184
rect 432290 307128 432295 307184
rect 429916 307126 432295 307128
rect 432229 307123 432295 307126
rect -960 306234 480 306324
rect 3693 306234 3759 306237
rect -960 306232 3759 306234
rect -960 306176 3698 306232
rect 3754 306176 3759 306232
rect -960 306174 3759 306176
rect -960 306084 480 306174
rect 3693 306171 3759 306174
rect 384481 306234 384547 306237
rect 510470 306234 510476 306236
rect 384481 306232 510476 306234
rect 384481 306176 384486 306232
rect 384542 306176 510476 306232
rect 384481 306174 510476 306176
rect 384481 306171 384547 306174
rect 510470 306172 510476 306174
rect 510540 306172 510546 306236
rect 384297 306098 384363 306101
rect 510153 306098 510219 306101
rect 384297 306096 510219 306098
rect 384297 306040 384302 306096
rect 384358 306040 510158 306096
rect 510214 306040 510219 306096
rect 384297 306038 510219 306040
rect 384297 306035 384363 306038
rect 510153 306035 510219 306038
rect 384665 305962 384731 305965
rect 510838 305962 510844 305964
rect 384665 305960 510844 305962
rect 384665 305904 384670 305960
rect 384726 305904 510844 305960
rect 384665 305902 510844 305904
rect 384665 305899 384731 305902
rect 510838 305900 510844 305902
rect 510908 305900 510914 305964
rect 381486 305764 381492 305828
rect 381556 305826 381562 305828
rect 510654 305826 510660 305828
rect 381556 305766 510660 305826
rect 381556 305764 381562 305766
rect 510654 305764 510660 305766
rect 510724 305764 510730 305828
rect 370497 305690 370563 305693
rect 512729 305690 512795 305693
rect 370497 305688 512795 305690
rect 370497 305632 370502 305688
rect 370558 305632 512734 305688
rect 512790 305632 512795 305688
rect 370497 305630 512795 305632
rect 370497 305627 370563 305630
rect 512729 305627 512795 305630
rect 361757 304466 361823 304469
rect 359812 304464 361823 304466
rect 359812 304408 361762 304464
rect 361818 304408 361823 304464
rect 359812 304406 361823 304408
rect 361757 304403 361823 304406
rect 382181 303242 382247 303245
rect 509601 303242 509667 303245
rect 382181 303240 509667 303242
rect 382181 303184 382186 303240
rect 382242 303184 509606 303240
rect 509662 303184 509667 303240
rect 382181 303182 509667 303184
rect 382181 303179 382247 303182
rect 509601 303179 509667 303182
rect 381905 303106 381971 303109
rect 511165 303106 511231 303109
rect 381905 303104 511231 303106
rect 381905 303048 381910 303104
rect 381966 303048 511170 303104
rect 511226 303048 511231 303104
rect 381905 303046 511231 303048
rect 381905 303043 381971 303046
rect 511165 303043 511231 303046
rect 376109 302970 376175 302973
rect 514150 302970 514156 302972
rect 376109 302968 514156 302970
rect 376109 302912 376114 302968
rect 376170 302912 514156 302968
rect 376109 302910 514156 302912
rect 376109 302907 376175 302910
rect 514150 302908 514156 302910
rect 514220 302908 514226 302972
rect 361113 302834 361179 302837
rect 512637 302834 512703 302837
rect 361113 302832 512703 302834
rect 361113 302776 361118 302832
rect 361174 302776 512642 302832
rect 512698 302776 512703 302832
rect 361113 302774 512703 302776
rect 361113 302771 361179 302774
rect 512637 302771 512703 302774
rect 370681 300250 370747 300253
rect 509693 300250 509759 300253
rect 370681 300248 509759 300250
rect 370681 300192 370686 300248
rect 370742 300192 509698 300248
rect 509754 300192 509759 300248
rect 370681 300190 509759 300192
rect 370681 300187 370747 300190
rect 509693 300187 509759 300190
rect 368013 300114 368079 300117
rect 514886 300114 514892 300116
rect 368013 300112 514892 300114
rect 368013 300056 368018 300112
rect 368074 300056 514892 300112
rect 368013 300054 514892 300056
rect 368013 300051 368079 300054
rect 514886 300052 514892 300054
rect 514956 300052 514962 300116
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 361757 293450 361823 293453
rect 359812 293448 361823 293450
rect 359812 293392 361762 293448
rect 361818 293392 361823 293448
rect 359812 293390 361823 293392
rect 361757 293387 361823 293390
rect -960 293178 480 293268
rect 3417 293178 3483 293181
rect -960 293176 3483 293178
rect -960 293120 3422 293176
rect 3478 293120 3483 293176
rect -960 293118 3483 293120
rect -960 293028 480 293118
rect 3417 293115 3483 293118
rect 372153 291818 372219 291821
rect 514702 291818 514708 291820
rect 372153 291816 514708 291818
rect 372153 291760 372158 291816
rect 372214 291760 514708 291816
rect 372153 291758 514708 291760
rect 372153 291755 372219 291758
rect 514702 291756 514708 291758
rect 514772 291756 514778 291820
rect 583520 285276 584960 285516
rect 361757 282434 361823 282437
rect 359812 282432 361823 282434
rect 359812 282376 361762 282432
rect 361818 282376 361823 282432
rect 359812 282374 361823 282376
rect 361757 282371 361823 282374
rect -960 279972 480 280212
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect 361757 271418 361823 271421
rect 359812 271416 361823 271418
rect 359812 271360 361762 271416
rect 361818 271360 361823 271416
rect 359812 271358 361823 271360
rect 361757 271355 361823 271358
rect -960 267202 480 267292
rect 3509 267202 3575 267205
rect -960 267200 3575 267202
rect -960 267144 3514 267200
rect 3570 267144 3575 267200
rect -960 267142 3575 267144
rect -960 267052 480 267142
rect 3509 267139 3575 267142
rect 456977 262714 457043 262717
rect 456977 262712 460092 262714
rect 456977 262656 456982 262712
rect 457038 262656 460092 262712
rect 456977 262654 460092 262656
rect 456977 262651 457043 262654
rect 529289 261626 529355 261629
rect 529289 261624 529490 261626
rect 529289 261568 529294 261624
rect 529350 261568 529490 261624
rect 529289 261566 529490 261568
rect 529289 261563 529355 261566
rect 529430 261052 529490 261566
rect 361757 260402 361823 260405
rect 359812 260400 361823 260402
rect 359812 260344 361762 260400
rect 361818 260344 361823 260400
rect 359812 260342 361823 260344
rect 361757 260339 361823 260342
rect 580257 258906 580323 258909
rect 583520 258906 584960 258996
rect 580257 258904 584960 258906
rect 580257 258848 580262 258904
rect 580318 258848 584960 258904
rect 580257 258846 584960 258848
rect 580257 258843 580323 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3601 254146 3667 254149
rect -960 254144 3667 254146
rect -960 254088 3606 254144
rect 3662 254088 3667 254144
rect -960 254086 3667 254088
rect -960 253996 480 254086
rect 3601 254083 3667 254086
rect 361757 249386 361823 249389
rect 359812 249384 361823 249386
rect 359812 249328 361762 249384
rect 361818 249328 361823 249384
rect 359812 249326 361823 249328
rect 361757 249323 361823 249326
rect 458081 248842 458147 248845
rect 458081 248840 460092 248842
rect 458081 248784 458086 248840
rect 458142 248784 460092 248840
rect 458081 248782 460092 248784
rect 458081 248779 458147 248782
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 531313 243674 531379 243677
rect 529828 243672 531379 243674
rect 529828 243616 531318 243672
rect 531374 243616 531379 243672
rect 529828 243614 531379 243616
rect 531313 243611 531379 243614
rect -960 241090 480 241180
rect 3785 241090 3851 241093
rect -960 241088 3851 241090
rect -960 241032 3790 241088
rect 3846 241032 3851 241088
rect -960 241030 3851 241032
rect -960 240940 480 241030
rect 3785 241027 3851 241030
rect 361757 238370 361823 238373
rect 359812 238368 361823 238370
rect 359812 238312 361762 238368
rect 361818 238312 361823 238368
rect 359812 238310 361823 238312
rect 361757 238307 361823 238310
rect 456701 234970 456767 234973
rect 456885 234970 456951 234973
rect 456701 234968 460092 234970
rect 456701 234912 456706 234968
rect 456762 234912 456890 234968
rect 456946 234912 460092 234968
rect 456701 234910 460092 234912
rect 456701 234907 456767 234910
rect 456885 234907 456951 234910
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 361757 227354 361823 227357
rect 359812 227352 361823 227354
rect 359812 227296 361762 227352
rect 361818 227296 361823 227352
rect 359812 227294 361823 227296
rect 361757 227291 361823 227294
rect 530117 226266 530183 226269
rect 529828 226264 530183 226266
rect 529828 226208 530122 226264
rect 530178 226208 530183 226264
rect 529828 226206 530183 226208
rect 530117 226203 530183 226206
rect 457897 221098 457963 221101
rect 459461 221098 459527 221101
rect 457897 221096 460092 221098
rect 457897 221040 457902 221096
rect 457958 221040 459466 221096
rect 459522 221040 460092 221096
rect 457897 221038 460092 221040
rect 457897 221035 457963 221038
rect 459461 221035 459527 221038
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect 361665 216338 361731 216341
rect 359812 216336 361731 216338
rect 359812 216280 361670 216336
rect 361726 216280 361731 216336
rect 359812 216278 361731 216280
rect 361665 216275 361731 216278
rect -960 214978 480 215068
rect 3877 214978 3943 214981
rect -960 214976 3943 214978
rect -960 214920 3882 214976
rect 3938 214920 3943 214976
rect -960 214918 3943 214920
rect -960 214828 480 214918
rect 3877 214915 3943 214918
rect 529933 209266 529999 209269
rect 529798 209264 529999 209266
rect 529798 209208 529938 209264
rect 529994 209208 529999 209264
rect 529798 209206 529999 209208
rect 529798 208828 529858 209206
rect 529933 209203 529999 209206
rect 456701 207226 456767 207229
rect 459369 207226 459435 207229
rect 456701 207224 460092 207226
rect 456701 207168 456706 207224
rect 456762 207168 459374 207224
rect 459430 207168 460092 207224
rect 456701 207166 460092 207168
rect 456701 207163 456767 207166
rect 459369 207163 459435 207166
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect 361757 205322 361823 205325
rect 359812 205320 361823 205322
rect 359812 205264 361762 205320
rect 361818 205264 361823 205320
rect 359812 205262 361823 205264
rect 361757 205259 361823 205262
rect -960 201922 480 202012
rect 3969 201922 4035 201925
rect -960 201920 4035 201922
rect -960 201864 3974 201920
rect 4030 201864 4035 201920
rect -960 201862 4035 201864
rect -960 201772 480 201862
rect 3969 201859 4035 201862
rect 361757 194306 361823 194309
rect 359812 194304 361823 194306
rect 359812 194248 361762 194304
rect 361818 194248 361823 194304
rect 359812 194246 361823 194248
rect 361757 194243 361823 194246
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 4061 188866 4127 188869
rect -960 188864 4127 188866
rect -960 188808 4066 188864
rect 4122 188808 4127 188864
rect -960 188806 4127 188808
rect -960 188716 480 188806
rect 4061 188803 4127 188806
rect 361757 183290 361823 183293
rect 359812 183288 361823 183290
rect 359812 183232 361762 183288
rect 361818 183232 361823 183288
rect 359812 183230 361823 183232
rect 361757 183227 361823 183230
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 361757 172274 361823 172277
rect 359812 172272 361823 172274
rect 359812 172216 361762 172272
rect 361818 172216 361823 172272
rect 359812 172214 361823 172216
rect 361757 172211 361823 172214
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3325 162890 3391 162893
rect -960 162888 3391 162890
rect -960 162832 3330 162888
rect 3386 162832 3391 162888
rect -960 162830 3391 162832
rect -960 162740 480 162830
rect 3325 162827 3391 162830
rect 421046 162692 421052 162756
rect 421116 162754 421122 162756
rect 421741 162754 421807 162757
rect 421116 162752 421807 162754
rect 421116 162696 421746 162752
rect 421802 162696 421807 162752
rect 421116 162694 421807 162696
rect 421116 162692 421122 162694
rect 421741 162691 421807 162694
rect 428406 162692 428412 162756
rect 428476 162754 428482 162756
rect 428641 162754 428707 162757
rect 428476 162752 428707 162754
rect 428476 162696 428646 162752
rect 428702 162696 428707 162752
rect 428476 162694 428707 162696
rect 428476 162692 428482 162694
rect 428641 162691 428707 162694
rect 361757 161258 361823 161261
rect 359812 161256 361823 161258
rect 359812 161200 361762 161256
rect 361818 161200 361823 161256
rect 359812 161198 361823 161200
rect 361757 161195 361823 161198
rect 452561 158402 452627 158405
rect 449758 158400 452627 158402
rect 449758 158344 452566 158400
rect 452622 158344 452627 158400
rect 449758 158342 452627 158344
rect 449758 158304 449818 158342
rect 452561 158339 452627 158342
rect 452377 157314 452443 157317
rect 449758 157312 452443 157314
rect 449758 157256 452382 157312
rect 452438 157256 452443 157312
rect 449758 157254 452443 157256
rect 449758 156944 449818 157254
rect 452377 157251 452443 157254
rect 452377 155818 452443 155821
rect 449758 155816 452443 155818
rect 449758 155760 452382 155816
rect 452438 155760 452443 155816
rect 449758 155758 452443 155760
rect 449758 155584 449818 155758
rect 452377 155755 452443 155758
rect 452377 154322 452443 154325
rect 449758 154320 452443 154322
rect 449758 154264 452382 154320
rect 452438 154264 452443 154320
rect 449758 154262 452443 154264
rect 449758 154224 449818 154262
rect 452377 154259 452443 154262
rect 452469 153098 452535 153101
rect 449758 153096 452535 153098
rect 449758 153040 452474 153096
rect 452530 153040 452535 153096
rect 449758 153038 452535 153040
rect 449758 152864 449818 153038
rect 452469 153035 452535 153038
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect 452285 151738 452351 151741
rect 449758 151736 452351 151738
rect 449758 151680 452290 151736
rect 452346 151680 452351 151736
rect 449758 151678 452351 151680
rect 449758 151504 449818 151678
rect 452285 151675 452351 151678
rect 452101 150378 452167 150381
rect 449758 150376 452167 150378
rect 449758 150320 452106 150376
rect 452162 150320 452167 150376
rect 449758 150318 452167 150320
rect 362585 150242 362651 150245
rect 359812 150240 362651 150242
rect 359812 150184 362590 150240
rect 362646 150184 362651 150240
rect 359812 150182 362651 150184
rect 362585 150179 362651 150182
rect 449758 150144 449818 150318
rect 452101 150315 452167 150318
rect -960 149834 480 149924
rect 3233 149834 3299 149837
rect -960 149832 3299 149834
rect -960 149776 3238 149832
rect 3294 149776 3299 149832
rect -960 149774 3299 149776
rect -960 149684 480 149774
rect 3233 149771 3299 149774
rect 452561 149018 452627 149021
rect 449758 149016 452627 149018
rect 449758 148960 452566 149016
rect 452622 148960 452627 149016
rect 449758 148958 452627 148960
rect 449758 148784 449818 148958
rect 452561 148955 452627 148958
rect 452561 147522 452627 147525
rect 449758 147520 452627 147522
rect 449758 147464 452566 147520
rect 452622 147464 452627 147520
rect 449758 147462 452627 147464
rect 449758 147424 449818 147462
rect 452561 147459 452627 147462
rect 452561 146162 452627 146165
rect 449758 146160 452627 146162
rect 449758 146104 452566 146160
rect 452622 146104 452627 146160
rect 449758 146102 452627 146104
rect 449758 146064 449818 146102
rect 452561 146099 452627 146102
rect 452561 144802 452627 144805
rect 449758 144800 452627 144802
rect 449758 144744 452566 144800
rect 452622 144744 452627 144800
rect 449758 144742 452627 144744
rect 449758 144704 449818 144742
rect 452561 144739 452627 144742
rect 452561 143442 452627 143445
rect 449758 143440 452627 143442
rect 449758 143384 452566 143440
rect 452622 143384 452627 143440
rect 449758 143382 452627 143384
rect 449758 143344 449818 143382
rect 452561 143379 452627 143382
rect 452561 142082 452627 142085
rect 449758 142080 452627 142082
rect 449758 142024 452566 142080
rect 452622 142024 452627 142080
rect 449758 142022 452627 142024
rect 449758 141984 449818 142022
rect 452561 142019 452627 142022
rect 452561 140722 452627 140725
rect 449758 140720 452627 140722
rect 449758 140664 452566 140720
rect 452622 140664 452627 140720
rect 449758 140662 452627 140664
rect 449758 140624 449818 140662
rect 452561 140659 452627 140662
rect 452561 139362 452627 139365
rect 449758 139360 452627 139362
rect 449758 139304 452566 139360
rect 452622 139304 452627 139360
rect 449758 139302 452627 139304
rect 449758 139264 449818 139302
rect 452561 139299 452627 139302
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 361757 139226 361823 139229
rect 359812 139224 361823 139226
rect 359812 139168 361762 139224
rect 361818 139168 361823 139224
rect 583520 139212 584960 139302
rect 359812 139166 361823 139168
rect 361757 139163 361823 139166
rect 452561 137866 452627 137869
rect 449788 137864 452627 137866
rect 449788 137808 452566 137864
rect 452622 137808 452627 137864
rect 449788 137806 452627 137808
rect 452561 137803 452627 137806
rect 539317 137730 539383 137733
rect 539317 137728 539426 137730
rect 539317 137672 539322 137728
rect 539378 137672 539426 137728
rect 539317 137667 539426 137672
rect 539366 137428 539426 137667
rect -960 136778 480 136868
rect 3366 136778 3372 136780
rect -960 136718 3372 136778
rect -960 136628 480 136718
rect 3366 136716 3372 136718
rect 3436 136716 3442 136780
rect 451549 136506 451615 136509
rect 449788 136504 451615 136506
rect 449788 136448 451554 136504
rect 451610 136448 451615 136504
rect 449788 136446 451615 136448
rect 451549 136443 451615 136446
rect 539317 135690 539383 135693
rect 539317 135688 539426 135690
rect 539317 135632 539322 135688
rect 539378 135632 539426 135688
rect 539317 135627 539426 135632
rect 539366 135388 539426 135627
rect 452561 135146 452627 135149
rect 449788 135144 452627 135146
rect 449788 135088 452566 135144
rect 452622 135088 452627 135144
rect 449788 135086 452627 135088
rect 452561 135083 452627 135086
rect 452561 133786 452627 133789
rect 449788 133784 452627 133786
rect 449788 133728 452566 133784
rect 452622 133728 452627 133784
rect 449788 133726 452627 133728
rect 452561 133723 452627 133726
rect 540329 133378 540395 133381
rect 539948 133376 540395 133378
rect 539948 133320 540334 133376
rect 540390 133320 540395 133376
rect 539948 133318 540395 133320
rect 540329 133315 540395 133318
rect 452561 132426 452627 132429
rect 449788 132424 452627 132426
rect 449788 132368 452566 132424
rect 452622 132368 452627 132424
rect 449788 132366 452627 132368
rect 452561 132363 452627 132366
rect 542721 131338 542787 131341
rect 539948 131336 542787 131338
rect 539948 131280 542726 131336
rect 542782 131280 542787 131336
rect 539948 131278 542787 131280
rect 542721 131275 542787 131278
rect 452561 131066 452627 131069
rect 449788 131064 452627 131066
rect 449788 131008 452566 131064
rect 452622 131008 452627 131064
rect 449788 131006 452627 131008
rect 452561 131003 452627 131006
rect 452561 129706 452627 129709
rect 449788 129704 452627 129706
rect 449788 129648 452566 129704
rect 452622 129648 452627 129704
rect 449788 129646 452627 129648
rect 452561 129643 452627 129646
rect 539358 129236 539364 129300
rect 539428 129236 539434 129300
rect 452285 128346 452351 128349
rect 449788 128344 452351 128346
rect 449788 128288 452290 128344
rect 452346 128288 452351 128344
rect 449788 128286 452351 128288
rect 452285 128283 452351 128286
rect 361757 128210 361823 128213
rect 359812 128208 361823 128210
rect 359812 128152 361762 128208
rect 361818 128152 361823 128208
rect 359812 128150 361823 128152
rect 361757 128147 361823 128150
rect 540237 127258 540303 127261
rect 539948 127256 540303 127258
rect 539948 127200 540242 127256
rect 540298 127200 540303 127256
rect 539948 127198 540303 127200
rect 540237 127195 540303 127198
rect 452377 126986 452443 126989
rect 449788 126984 452443 126986
rect 449788 126928 452382 126984
rect 452438 126928 452443 126984
rect 449788 126926 452443 126928
rect 452377 126923 452443 126926
rect 452193 126306 452259 126309
rect 449758 126304 452259 126306
rect 449758 126248 452198 126304
rect 452254 126248 452259 126304
rect 449758 126246 452259 126248
rect 449758 125664 449818 126246
rect 452193 126243 452259 126246
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect 540145 125218 540211 125221
rect 539948 125216 540211 125218
rect 539948 125160 540150 125216
rect 540206 125160 540211 125216
rect 539948 125158 540211 125160
rect 540145 125155 540211 125158
rect 452009 124946 452075 124949
rect 449758 124944 452075 124946
rect 449758 124888 452014 124944
rect 452070 124888 452075 124944
rect 449758 124886 452075 124888
rect 449758 124304 449818 124886
rect 452009 124883 452075 124886
rect -960 123572 480 123812
rect 451917 123586 451983 123589
rect 449758 123584 451983 123586
rect 449758 123528 451922 123584
rect 451978 123528 451983 123584
rect 449758 123526 451983 123528
rect 449758 122944 449818 123526
rect 451917 123523 451983 123526
rect 543089 123178 543155 123181
rect 539948 123176 543155 123178
rect 539948 123120 543094 123176
rect 543150 123120 543155 123176
rect 539948 123118 543155 123120
rect 543089 123115 543155 123118
rect 451917 121546 451983 121549
rect 449788 121544 451983 121546
rect 449788 121488 451922 121544
rect 451978 121488 451983 121544
rect 449788 121486 451983 121488
rect 451917 121483 451983 121486
rect 542445 121138 542511 121141
rect 539948 121136 542511 121138
rect 539948 121080 542450 121136
rect 542506 121080 542511 121136
rect 539948 121078 542511 121080
rect 542445 121075 542511 121078
rect 542997 119098 543063 119101
rect 539948 119096 543063 119098
rect 539948 119040 543002 119096
rect 543058 119040 543063 119096
rect 539948 119038 543063 119040
rect 542997 119035 543063 119038
rect 540053 117330 540119 117333
rect 539918 117328 540119 117330
rect 539918 117272 540058 117328
rect 540114 117272 540119 117328
rect 539918 117270 540119 117272
rect 361757 117194 361823 117197
rect 359812 117192 361823 117194
rect 359812 117136 361762 117192
rect 361818 117136 361823 117192
rect 359812 117134 361823 117136
rect 361757 117131 361823 117134
rect 539918 117028 539978 117270
rect 540053 117267 540119 117270
rect 541525 115018 541591 115021
rect 539948 115016 541591 115018
rect 539948 114960 541530 115016
rect 541586 114960 541591 115016
rect 539948 114958 541591 114960
rect 541525 114955 541591 114958
rect 539918 112845 539978 112948
rect 539918 112840 540027 112845
rect 539918 112784 539966 112840
rect 540022 112784 540027 112840
rect 539918 112782 540027 112784
rect 539961 112779 540027 112782
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect 541157 110938 541223 110941
rect 539948 110936 541223 110938
rect 539948 110880 541162 110936
rect 541218 110880 541223 110936
rect 539948 110878 541223 110880
rect 541157 110875 541223 110878
rect -960 110666 480 110756
rect 3550 110666 3556 110668
rect -960 110606 3556 110666
rect -960 110516 480 110606
rect 3550 110604 3556 110606
rect 3620 110604 3626 110668
rect 539869 109170 539935 109173
rect 539869 109168 539978 109170
rect 539869 109112 539874 109168
rect 539930 109112 539978 109168
rect 539869 109107 539978 109112
rect 539918 108868 539978 109107
rect 541433 106858 541499 106861
rect 539948 106856 541499 106858
rect 539948 106800 541438 106856
rect 541494 106800 541499 106856
rect 539948 106798 541499 106800
rect 541433 106795 541499 106798
rect 361757 106178 361823 106181
rect 359812 106176 361823 106178
rect 359812 106120 361762 106176
rect 361818 106120 361823 106176
rect 359812 106118 361823 106120
rect 361757 106115 361823 106118
rect 541341 104818 541407 104821
rect 539948 104816 541407 104818
rect 539948 104760 541346 104816
rect 541402 104760 541407 104816
rect 539948 104758 541407 104760
rect 541341 104755 541407 104758
rect 541065 102778 541131 102781
rect 539948 102776 541131 102778
rect 539948 102720 541070 102776
rect 541126 102720 541131 102776
rect 539948 102718 541131 102720
rect 541065 102715 541131 102718
rect 539734 100605 539794 100708
rect 539734 100600 539843 100605
rect 539734 100544 539782 100600
rect 539838 100544 539843 100600
rect 539734 100542 539843 100544
rect 539777 100539 539843 100542
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect 539593 99242 539659 99245
rect 539550 99240 539659 99242
rect 539550 99184 539598 99240
rect 539654 99184 539659 99240
rect 539550 99179 539659 99184
rect 539550 98668 539610 99179
rect -960 97610 480 97700
rect 3693 97610 3759 97613
rect -960 97608 3759 97610
rect -960 97552 3698 97608
rect 3754 97552 3759 97608
rect -960 97550 3759 97552
rect -960 97460 480 97550
rect 3693 97547 3759 97550
rect 542905 96658 542971 96661
rect 539948 96656 542971 96658
rect 539948 96600 542910 96656
rect 542966 96600 542971 96656
rect 539948 96598 542971 96600
rect 542905 96595 542971 96598
rect 362677 95162 362743 95165
rect 359812 95160 362743 95162
rect 359812 95104 362682 95160
rect 362738 95104 362743 95160
rect 359812 95102 362743 95104
rect 362677 95099 362743 95102
rect 543181 94618 543247 94621
rect 539948 94616 543247 94618
rect 539948 94560 543186 94616
rect 543242 94560 543247 94616
rect 539948 94558 543247 94560
rect 543181 94555 543247 94558
rect 542813 92578 542879 92581
rect 539948 92576 542879 92578
rect 539948 92520 542818 92576
rect 542874 92520 542879 92576
rect 539948 92518 542879 92520
rect 542813 92515 542879 92518
rect 542629 90538 542695 90541
rect 539948 90536 542695 90538
rect 539948 90480 542634 90536
rect 542690 90480 542695 90536
rect 539948 90478 542695 90480
rect 542629 90475 542695 90478
rect 541249 88498 541315 88501
rect 539948 88496 541315 88498
rect 539948 88440 541254 88496
rect 541310 88440 541315 88496
rect 539948 88438 541315 88440
rect 541249 88435 541315 88438
rect 539685 86866 539751 86869
rect 539685 86864 539794 86866
rect 539685 86808 539690 86864
rect 539746 86808 539794 86864
rect 539685 86803 539794 86808
rect 539734 86428 539794 86803
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 542537 84418 542603 84421
rect 539948 84416 542603 84418
rect 539948 84360 542542 84416
rect 542598 84360 542603 84416
rect 539948 84358 542603 84360
rect 542537 84355 542603 84358
rect 361757 84146 361823 84149
rect 359812 84144 361823 84146
rect 359812 84088 361762 84144
rect 361818 84088 361823 84144
rect 359812 84086 361823 84088
rect 361757 84083 361823 84086
rect 540973 82378 541039 82381
rect 539948 82376 541039 82378
rect 539948 82320 540978 82376
rect 541034 82320 541039 82376
rect 539948 82318 541039 82320
rect 540973 82315 541039 82318
rect 361757 73130 361823 73133
rect 359812 73128 361823 73130
rect 359812 73072 361762 73128
rect 361818 73072 361823 73128
rect 359812 73070 361823 73072
rect 361757 73067 361823 73070
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3141 71634 3207 71637
rect -960 71632 3207 71634
rect -960 71576 3146 71632
rect 3202 71576 3207 71632
rect -960 71574 3207 71576
rect -960 71484 480 71574
rect 3141 71571 3207 71574
rect 462313 67554 462379 67557
rect 462497 67554 462563 67557
rect 460828 67552 462563 67554
rect 460828 67496 462318 67552
rect 462374 67496 462502 67552
rect 462558 67496 462563 67552
rect 460828 67494 462563 67496
rect 462313 67491 462379 67494
rect 462497 67491 462563 67494
rect 361757 62114 361823 62117
rect 359812 62112 361823 62114
rect 359812 62056 361762 62112
rect 361818 62056 361823 62112
rect 359812 62054 361823 62056
rect 361757 62051 361823 62054
rect 3417 59938 3483 59941
rect 22686 59938 22692 59940
rect 3417 59936 22692 59938
rect 3417 59880 3422 59936
rect 3478 59880 22692 59936
rect 3417 59878 22692 59880
rect 3417 59875 3483 59878
rect 22686 59876 22692 59878
rect 22756 59876 22762 59940
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3417 58578 3483 58581
rect -960 58576 3483 58578
rect -960 58520 3422 58576
rect 3478 58520 3483 58576
rect -960 58518 3483 58520
rect -960 58428 480 58518
rect 3417 58515 3483 58518
rect 361757 51098 361823 51101
rect 359812 51096 361823 51098
rect 359812 51040 361762 51096
rect 361818 51040 361823 51096
rect 359812 51038 361823 51040
rect 361757 51035 361823 51038
rect 19333 49602 19399 49605
rect 22134 49602 22140 49604
rect 19333 49600 22140 49602
rect 19333 49544 19338 49600
rect 19394 49544 22140 49600
rect 19333 49542 22140 49544
rect 19333 49539 19399 49542
rect 22134 49540 22140 49542
rect 22204 49540 22210 49604
rect 540605 48922 540671 48925
rect 540605 48920 540714 48922
rect 540605 48864 540610 48920
rect 540666 48864 540714 48920
rect 540605 48859 540714 48864
rect 540654 48348 540714 48859
rect 3366 46956 3372 47020
rect 3436 47018 3442 47020
rect 384849 47018 384915 47021
rect 3436 47016 384915 47018
rect 3436 46960 384854 47016
rect 384910 46960 384915 47016
rect 3436 46958 384915 46960
rect 3436 46956 3442 46958
rect 384849 46955 384915 46958
rect 3550 46820 3556 46884
rect 3620 46882 3626 46884
rect 385769 46882 385835 46885
rect 3620 46880 385835 46882
rect 3620 46824 385774 46880
rect 385830 46824 385835 46880
rect 3620 46822 385835 46824
rect 3620 46820 3626 46822
rect 385769 46819 385835 46822
rect 21357 46746 21423 46749
rect 384757 46746 384823 46749
rect 21357 46744 384823 46746
rect 21357 46688 21362 46744
rect 21418 46688 384762 46744
rect 384818 46688 384823 46744
rect 21357 46686 384823 46688
rect 21357 46683 21423 46686
rect 384757 46683 384823 46686
rect 22686 46548 22692 46612
rect 22756 46610 22762 46612
rect 378593 46610 378659 46613
rect 22756 46608 378659 46610
rect 22756 46552 378598 46608
rect 378654 46552 378659 46608
rect 22756 46550 378659 46552
rect 22756 46548 22762 46550
rect 378593 46547 378659 46550
rect 22134 46412 22140 46476
rect 22204 46474 22210 46476
rect 361389 46474 361455 46477
rect 22204 46472 361455 46474
rect 22204 46416 361394 46472
rect 361450 46416 361455 46472
rect 22204 46414 361455 46416
rect 22204 46412 22210 46414
rect 361389 46411 361455 46414
rect 578877 46338 578943 46341
rect 583520 46338 584960 46428
rect 578877 46336 584960 46338
rect 578877 46280 578882 46336
rect 578938 46280 584960 46336
rect 578877 46278 584960 46280
rect 578877 46275 578943 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3509 45522 3575 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 46933 44842 46999 44845
rect 381486 44842 381492 44844
rect 46933 44840 381492 44842
rect 46933 44784 46938 44840
rect 46994 44784 381492 44840
rect 46933 44782 381492 44784
rect 46933 44779 46999 44782
rect 381486 44780 381492 44782
rect 381556 44780 381562 44844
rect 536833 41034 536899 41037
rect 536833 41032 540132 41034
rect 536833 40976 536838 41032
rect 536894 40976 540132 41032
rect 536833 40974 540132 40976
rect 536833 40971 536899 40974
rect 536833 33690 536899 33693
rect 536833 33688 540132 33690
rect 536833 33632 536838 33688
rect 536894 33632 540132 33688
rect 536833 33630 540132 33632
rect 536833 33627 536899 33630
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 17033 4042 17099 4045
rect 370681 4042 370747 4045
rect 17033 4040 370747 4042
rect 17033 3984 17038 4040
rect 17094 3984 370686 4040
rect 370742 3984 370747 4040
rect 17033 3982 370747 3984
rect 17033 3979 17099 3982
rect 370681 3979 370747 3982
rect 5257 3906 5323 3909
rect 361021 3906 361087 3909
rect 5257 3904 361087 3906
rect 5257 3848 5262 3904
rect 5318 3848 361026 3904
rect 361082 3848 361087 3904
rect 5257 3846 361087 3848
rect 5257 3843 5323 3846
rect 361021 3843 361087 3846
rect 8753 3770 8819 3773
rect 365161 3770 365227 3773
rect 8753 3768 365227 3770
rect 8753 3712 8758 3768
rect 8814 3712 365166 3768
rect 365222 3712 365227 3768
rect 8753 3710 365227 3712
rect 8753 3707 8819 3710
rect 365161 3707 365227 3710
rect 13537 3634 13603 3637
rect 370497 3634 370563 3637
rect 13537 3632 370563 3634
rect 13537 3576 13542 3632
rect 13598 3576 370502 3632
rect 370558 3576 370563 3632
rect 13537 3574 370563 3576
rect 13537 3571 13603 3574
rect 370497 3571 370563 3574
rect 24209 3498 24275 3501
rect 383009 3498 383075 3501
rect 24209 3496 383075 3498
rect 24209 3440 24214 3496
rect 24270 3440 383014 3496
rect 383070 3440 383075 3496
rect 24209 3438 383075 3440
rect 24209 3435 24275 3438
rect 383009 3435 383075 3438
rect 1669 3362 1735 3365
rect 384481 3362 384547 3365
rect 1669 3360 384547 3362
rect 1669 3304 1674 3360
rect 1730 3304 384486 3360
rect 384542 3304 384547 3360
rect 1669 3302 384547 3304
rect 1669 3299 1735 3302
rect 384481 3299 384547 3302
<< via3 >>
rect 450492 700572 450556 700636
rect 444236 700436 444300 700500
rect 447732 700300 447796 700364
rect 526300 699756 526364 699820
rect 559420 699756 559484 699820
rect 450676 683980 450740 684044
rect 446260 683844 446324 683908
rect 446444 683708 446508 683772
rect 3556 683300 3620 683364
rect 3740 683164 3804 683228
rect 3372 682892 3436 682956
rect 447916 682756 447980 682820
rect 3740 671196 3804 671260
rect 458036 665212 458100 665276
rect 457852 662492 457916 662556
rect 459140 630668 459204 630732
rect 3556 619108 3620 619172
rect 3372 606052 3436 606116
rect 474780 599524 474844 599588
rect 476436 598164 476500 598228
rect 478828 542948 478892 543012
rect 458036 522276 458100 522340
rect 457852 521052 457916 521116
rect 474412 520916 474476 520980
rect 472020 519556 472084 519620
rect 474596 519420 474660 519484
rect 487108 453868 487172 453932
rect 459140 391172 459204 391236
rect 472020 388996 472084 389060
rect 474412 389056 474476 389060
rect 474412 389000 474426 389056
rect 474426 389000 474476 389056
rect 474412 388996 474476 389000
rect 474780 388996 474844 389060
rect 476436 388996 476500 389060
rect 478828 388996 478892 389060
rect 474596 388860 474660 388924
rect 487108 385596 487172 385660
rect 510660 342756 510724 342820
rect 421052 334460 421116 334524
rect 428412 334460 428476 334524
rect 514892 332964 514956 333028
rect 514340 330788 514404 330852
rect 514708 330244 514772 330308
rect 517836 329156 517900 329220
rect 514156 328068 514220 328132
rect 510844 327524 510908 327588
rect 511212 326436 511276 326500
rect 511028 325892 511092 325956
rect 510292 324804 510356 324868
rect 510476 323716 510540 323780
rect 510292 321812 510356 321876
rect 511028 321676 511092 321740
rect 559420 321404 559484 321468
rect 447732 321268 447796 321332
rect 510844 321268 510908 321332
rect 444236 320996 444300 321060
rect 450492 320860 450556 320924
rect 514340 320860 514404 320924
rect 517836 320724 517900 320788
rect 447916 320044 447980 320108
rect 526300 320044 526364 320108
rect 450676 319908 450740 319972
rect 446260 319772 446324 319836
rect 446444 319500 446508 319564
rect 538260 313924 538324 313988
rect 510476 306172 510540 306236
rect 510844 305900 510908 305964
rect 381492 305764 381556 305828
rect 510660 305764 510724 305828
rect 514156 302908 514220 302972
rect 514892 300052 514956 300116
rect 514708 291756 514772 291820
rect 421052 162692 421116 162756
rect 428412 162692 428476 162756
rect 3372 136716 3436 136780
rect 539364 129236 539428 129300
rect 3556 110604 3620 110668
rect 22692 59876 22756 59940
rect 22140 49540 22204 49604
rect 3372 46956 3436 47020
rect 3556 46820 3620 46884
rect 22692 46548 22756 46612
rect 22140 46412 22204 46476
rect 381492 44780 381556 44844
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 677494 -8106 711002
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 -8106 677494
rect -8726 677174 -8106 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 -8106 677174
rect -8726 641494 -8106 676938
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 -8106 641494
rect -8726 641174 -8106 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 -8106 641174
rect -8726 605494 -8106 640938
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 -8106 605494
rect -8726 605174 -8106 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 -8106 605174
rect -8726 569494 -8106 604938
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 -8106 569494
rect -8726 569174 -8106 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 -8106 569174
rect -8726 533494 -8106 568938
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 -8106 533494
rect -8726 533174 -8106 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 -8106 533174
rect -8726 497494 -8106 532938
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 -8106 497494
rect -8726 497174 -8106 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 -8106 497174
rect -8726 461494 -8106 496938
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 -8106 461494
rect -8726 461174 -8106 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 -8106 461174
rect -8726 425494 -8106 460938
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 -8106 425494
rect -8726 425174 -8106 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 -8106 425174
rect -8726 389494 -8106 424938
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 -8106 389494
rect -8726 389174 -8106 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 -8106 389174
rect -8726 353494 -8106 388938
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 -8106 353494
rect -8726 353174 -8106 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 -8106 353174
rect -8726 317494 -8106 352938
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 -8106 317494
rect -8726 317174 -8106 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 -8106 317174
rect -8726 281494 -8106 316938
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 -8106 281494
rect -8726 281174 -8106 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 -8106 281174
rect -8726 245494 -8106 280938
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 -8106 245494
rect -8726 245174 -8106 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 -8106 245174
rect -8726 209494 -8106 244938
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 -8106 209494
rect -8726 209174 -8106 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 -8106 209174
rect -8726 173494 -8106 208938
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 -8106 173494
rect -8726 173174 -8106 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 -8106 173174
rect -8726 137494 -8106 172938
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 -8106 137494
rect -8726 137174 -8106 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 -8106 137174
rect -8726 101494 -8106 136938
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 -8106 101494
rect -8726 101174 -8106 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 -8106 101174
rect -8726 65494 -8106 100938
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 -8106 65494
rect -8726 65174 -8106 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 -8106 65174
rect -8726 29494 -8106 64938
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 -8106 29494
rect -8726 29174 -8106 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 -8106 29174
rect -8726 -7066 -8106 28938
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 673774 -7146 710042
rect -7766 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 -7146 673774
rect -7766 673454 -7146 673538
rect -7766 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 -7146 673454
rect -7766 637774 -7146 673218
rect -7766 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 -7146 637774
rect -7766 637454 -7146 637538
rect -7766 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 -7146 637454
rect -7766 601774 -7146 637218
rect -7766 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 -7146 601774
rect -7766 601454 -7146 601538
rect -7766 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 -7146 601454
rect -7766 565774 -7146 601218
rect -7766 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 -7146 565774
rect -7766 565454 -7146 565538
rect -7766 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 -7146 565454
rect -7766 529774 -7146 565218
rect -7766 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 -7146 529774
rect -7766 529454 -7146 529538
rect -7766 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 -7146 529454
rect -7766 493774 -7146 529218
rect -7766 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 -7146 493774
rect -7766 493454 -7146 493538
rect -7766 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 -7146 493454
rect -7766 457774 -7146 493218
rect -7766 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 -7146 457774
rect -7766 457454 -7146 457538
rect -7766 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 -7146 457454
rect -7766 421774 -7146 457218
rect -7766 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 -7146 421774
rect -7766 421454 -7146 421538
rect -7766 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 -7146 421454
rect -7766 385774 -7146 421218
rect -7766 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 -7146 385774
rect -7766 385454 -7146 385538
rect -7766 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 -7146 385454
rect -7766 349774 -7146 385218
rect -7766 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 -7146 349774
rect -7766 349454 -7146 349538
rect -7766 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 -7146 349454
rect -7766 313774 -7146 349218
rect -7766 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 -7146 313774
rect -7766 313454 -7146 313538
rect -7766 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 -7146 313454
rect -7766 277774 -7146 313218
rect -7766 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 -7146 277774
rect -7766 277454 -7146 277538
rect -7766 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 -7146 277454
rect -7766 241774 -7146 277218
rect -7766 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 -7146 241774
rect -7766 241454 -7146 241538
rect -7766 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 -7146 241454
rect -7766 205774 -7146 241218
rect -7766 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 -7146 205774
rect -7766 205454 -7146 205538
rect -7766 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 -7146 205454
rect -7766 169774 -7146 205218
rect -7766 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 -7146 169774
rect -7766 169454 -7146 169538
rect -7766 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 -7146 169454
rect -7766 133774 -7146 169218
rect -7766 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 -7146 133774
rect -7766 133454 -7146 133538
rect -7766 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 -7146 133454
rect -7766 97774 -7146 133218
rect -7766 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 -7146 97774
rect -7766 97454 -7146 97538
rect -7766 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 -7146 97454
rect -7766 61774 -7146 97218
rect -7766 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 -7146 61774
rect -7766 61454 -7146 61538
rect -7766 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 -7146 61454
rect -7766 25774 -7146 61218
rect -7766 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 -7146 25774
rect -7766 25454 -7146 25538
rect -7766 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 -7146 25454
rect -7766 -6106 -7146 25218
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 670054 -6186 709082
rect -6806 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 -6186 670054
rect -6806 669734 -6186 669818
rect -6806 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 -6186 669734
rect -6806 634054 -6186 669498
rect -6806 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 -6186 634054
rect -6806 633734 -6186 633818
rect -6806 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 -6186 633734
rect -6806 598054 -6186 633498
rect -6806 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 -6186 598054
rect -6806 597734 -6186 597818
rect -6806 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 -6186 597734
rect -6806 562054 -6186 597498
rect -6806 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 -6186 562054
rect -6806 561734 -6186 561818
rect -6806 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 -6186 561734
rect -6806 526054 -6186 561498
rect -6806 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 -6186 526054
rect -6806 525734 -6186 525818
rect -6806 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 -6186 525734
rect -6806 490054 -6186 525498
rect -6806 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 -6186 490054
rect -6806 489734 -6186 489818
rect -6806 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 -6186 489734
rect -6806 454054 -6186 489498
rect -6806 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 -6186 454054
rect -6806 453734 -6186 453818
rect -6806 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 -6186 453734
rect -6806 418054 -6186 453498
rect -6806 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 -6186 418054
rect -6806 417734 -6186 417818
rect -6806 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 -6186 417734
rect -6806 382054 -6186 417498
rect -6806 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 -6186 382054
rect -6806 381734 -6186 381818
rect -6806 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 -6186 381734
rect -6806 346054 -6186 381498
rect -6806 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 -6186 346054
rect -6806 345734 -6186 345818
rect -6806 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 -6186 345734
rect -6806 310054 -6186 345498
rect -6806 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 -6186 310054
rect -6806 309734 -6186 309818
rect -6806 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 -6186 309734
rect -6806 274054 -6186 309498
rect -6806 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 -6186 274054
rect -6806 273734 -6186 273818
rect -6806 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 -6186 273734
rect -6806 238054 -6186 273498
rect -6806 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 -6186 238054
rect -6806 237734 -6186 237818
rect -6806 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 -6186 237734
rect -6806 202054 -6186 237498
rect -6806 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 -6186 202054
rect -6806 201734 -6186 201818
rect -6806 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 -6186 201734
rect -6806 166054 -6186 201498
rect -6806 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 -6186 166054
rect -6806 165734 -6186 165818
rect -6806 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 -6186 165734
rect -6806 130054 -6186 165498
rect -6806 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 -6186 130054
rect -6806 129734 -6186 129818
rect -6806 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 -6186 129734
rect -6806 94054 -6186 129498
rect -6806 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 -6186 94054
rect -6806 93734 -6186 93818
rect -6806 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 -6186 93734
rect -6806 58054 -6186 93498
rect -6806 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 -6186 58054
rect -6806 57734 -6186 57818
rect -6806 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 -6186 57734
rect -6806 22054 -6186 57498
rect -6806 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 -6186 22054
rect -6806 21734 -6186 21818
rect -6806 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 -6186 21734
rect -6806 -5146 -6186 21498
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 666334 -5226 708122
rect -5846 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 -5226 666334
rect -5846 666014 -5226 666098
rect -5846 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 -5226 666014
rect -5846 630334 -5226 665778
rect -5846 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 -5226 630334
rect -5846 630014 -5226 630098
rect -5846 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 -5226 630014
rect -5846 594334 -5226 629778
rect -5846 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 -5226 594334
rect -5846 594014 -5226 594098
rect -5846 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 -5226 594014
rect -5846 558334 -5226 593778
rect -5846 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 -5226 558334
rect -5846 558014 -5226 558098
rect -5846 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 -5226 558014
rect -5846 522334 -5226 557778
rect -5846 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 -5226 522334
rect -5846 522014 -5226 522098
rect -5846 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 -5226 522014
rect -5846 486334 -5226 521778
rect -5846 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 -5226 486334
rect -5846 486014 -5226 486098
rect -5846 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 -5226 486014
rect -5846 450334 -5226 485778
rect -5846 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 -5226 450334
rect -5846 450014 -5226 450098
rect -5846 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 -5226 450014
rect -5846 414334 -5226 449778
rect -5846 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 -5226 414334
rect -5846 414014 -5226 414098
rect -5846 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 -5226 414014
rect -5846 378334 -5226 413778
rect -5846 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 -5226 378334
rect -5846 378014 -5226 378098
rect -5846 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 -5226 378014
rect -5846 342334 -5226 377778
rect -5846 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 -5226 342334
rect -5846 342014 -5226 342098
rect -5846 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 -5226 342014
rect -5846 306334 -5226 341778
rect -5846 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 -5226 306334
rect -5846 306014 -5226 306098
rect -5846 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 -5226 306014
rect -5846 270334 -5226 305778
rect -5846 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 -5226 270334
rect -5846 270014 -5226 270098
rect -5846 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 -5226 270014
rect -5846 234334 -5226 269778
rect -5846 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 -5226 234334
rect -5846 234014 -5226 234098
rect -5846 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 -5226 234014
rect -5846 198334 -5226 233778
rect -5846 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 -5226 198334
rect -5846 198014 -5226 198098
rect -5846 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 -5226 198014
rect -5846 162334 -5226 197778
rect -5846 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 -5226 162334
rect -5846 162014 -5226 162098
rect -5846 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 -5226 162014
rect -5846 126334 -5226 161778
rect -5846 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 -5226 126334
rect -5846 126014 -5226 126098
rect -5846 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 -5226 126014
rect -5846 90334 -5226 125778
rect -5846 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 -5226 90334
rect -5846 90014 -5226 90098
rect -5846 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 -5226 90014
rect -5846 54334 -5226 89778
rect -5846 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 -5226 54334
rect -5846 54014 -5226 54098
rect -5846 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 -5226 54014
rect -5846 18334 -5226 53778
rect -5846 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 -5226 18334
rect -5846 18014 -5226 18098
rect -5846 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 -5226 18014
rect -5846 -4186 -5226 17778
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 698614 -4266 707162
rect -4886 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 -4266 698614
rect -4886 698294 -4266 698378
rect -4886 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 -4266 698294
rect -4886 662614 -4266 698058
rect -4886 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 -4266 662614
rect -4886 662294 -4266 662378
rect -4886 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 -4266 662294
rect -4886 626614 -4266 662058
rect -4886 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 -4266 626614
rect -4886 626294 -4266 626378
rect -4886 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 -4266 626294
rect -4886 590614 -4266 626058
rect -4886 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 -4266 590614
rect -4886 590294 -4266 590378
rect -4886 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 -4266 590294
rect -4886 554614 -4266 590058
rect -4886 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 -4266 554614
rect -4886 554294 -4266 554378
rect -4886 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 -4266 554294
rect -4886 518614 -4266 554058
rect -4886 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 -4266 518614
rect -4886 518294 -4266 518378
rect -4886 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 -4266 518294
rect -4886 482614 -4266 518058
rect -4886 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 -4266 482614
rect -4886 482294 -4266 482378
rect -4886 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 -4266 482294
rect -4886 446614 -4266 482058
rect -4886 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 -4266 446614
rect -4886 446294 -4266 446378
rect -4886 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 -4266 446294
rect -4886 410614 -4266 446058
rect -4886 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 -4266 410614
rect -4886 410294 -4266 410378
rect -4886 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 -4266 410294
rect -4886 374614 -4266 410058
rect -4886 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 -4266 374614
rect -4886 374294 -4266 374378
rect -4886 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 -4266 374294
rect -4886 338614 -4266 374058
rect -4886 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 -4266 338614
rect -4886 338294 -4266 338378
rect -4886 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 -4266 338294
rect -4886 302614 -4266 338058
rect -4886 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 -4266 302614
rect -4886 302294 -4266 302378
rect -4886 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 -4266 302294
rect -4886 266614 -4266 302058
rect -4886 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 -4266 266614
rect -4886 266294 -4266 266378
rect -4886 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 -4266 266294
rect -4886 230614 -4266 266058
rect -4886 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 -4266 230614
rect -4886 230294 -4266 230378
rect -4886 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 -4266 230294
rect -4886 194614 -4266 230058
rect -4886 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 -4266 194614
rect -4886 194294 -4266 194378
rect -4886 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 -4266 194294
rect -4886 158614 -4266 194058
rect -4886 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 -4266 158614
rect -4886 158294 -4266 158378
rect -4886 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 -4266 158294
rect -4886 122614 -4266 158058
rect -4886 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 -4266 122614
rect -4886 122294 -4266 122378
rect -4886 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 -4266 122294
rect -4886 86614 -4266 122058
rect -4886 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 -4266 86614
rect -4886 86294 -4266 86378
rect -4886 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 -4266 86294
rect -4886 50614 -4266 86058
rect -4886 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 -4266 50614
rect -4886 50294 -4266 50378
rect -4886 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 -4266 50294
rect -4886 14614 -4266 50058
rect -4886 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 -4266 14614
rect -4886 14294 -4266 14378
rect -4886 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 -4266 14294
rect -4886 -3226 -4266 14058
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 694894 -3306 706202
rect -3926 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 -3306 694894
rect -3926 694574 -3306 694658
rect -3926 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 -3306 694574
rect -3926 658894 -3306 694338
rect -3926 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 -3306 658894
rect -3926 658574 -3306 658658
rect -3926 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 -3306 658574
rect -3926 622894 -3306 658338
rect -3926 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 -3306 622894
rect -3926 622574 -3306 622658
rect -3926 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 -3306 622574
rect -3926 586894 -3306 622338
rect -3926 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 -3306 586894
rect -3926 586574 -3306 586658
rect -3926 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 -3306 586574
rect -3926 550894 -3306 586338
rect -3926 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 -3306 550894
rect -3926 550574 -3306 550658
rect -3926 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 -3306 550574
rect -3926 514894 -3306 550338
rect -3926 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 -3306 514894
rect -3926 514574 -3306 514658
rect -3926 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 -3306 514574
rect -3926 478894 -3306 514338
rect -3926 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 -3306 478894
rect -3926 478574 -3306 478658
rect -3926 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 -3306 478574
rect -3926 442894 -3306 478338
rect -3926 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 -3306 442894
rect -3926 442574 -3306 442658
rect -3926 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 -3306 442574
rect -3926 406894 -3306 442338
rect -3926 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 -3306 406894
rect -3926 406574 -3306 406658
rect -3926 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 -3306 406574
rect -3926 370894 -3306 406338
rect -3926 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 -3306 370894
rect -3926 370574 -3306 370658
rect -3926 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 -3306 370574
rect -3926 334894 -3306 370338
rect -3926 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 -3306 334894
rect -3926 334574 -3306 334658
rect -3926 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 -3306 334574
rect -3926 298894 -3306 334338
rect -3926 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 -3306 298894
rect -3926 298574 -3306 298658
rect -3926 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 -3306 298574
rect -3926 262894 -3306 298338
rect -3926 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 -3306 262894
rect -3926 262574 -3306 262658
rect -3926 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 -3306 262574
rect -3926 226894 -3306 262338
rect -3926 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 -3306 226894
rect -3926 226574 -3306 226658
rect -3926 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 -3306 226574
rect -3926 190894 -3306 226338
rect -3926 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 -3306 190894
rect -3926 190574 -3306 190658
rect -3926 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 -3306 190574
rect -3926 154894 -3306 190338
rect -3926 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 -3306 154894
rect -3926 154574 -3306 154658
rect -3926 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 -3306 154574
rect -3926 118894 -3306 154338
rect -3926 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 -3306 118894
rect -3926 118574 -3306 118658
rect -3926 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 -3306 118574
rect -3926 82894 -3306 118338
rect -3926 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 -3306 82894
rect -3926 82574 -3306 82658
rect -3926 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 -3306 82574
rect -3926 46894 -3306 82338
rect -3926 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 -3306 46894
rect -3926 46574 -3306 46658
rect -3926 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 -3306 46574
rect -3926 10894 -3306 46338
rect -3926 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 -3306 10894
rect -3926 10574 -3306 10658
rect -3926 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 -3306 10574
rect -3926 -2266 -3306 10338
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691174 -2346 705242
rect -2966 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 -2346 691174
rect -2966 690854 -2346 690938
rect -2966 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 -2346 690854
rect -2966 655174 -2346 690618
rect -2966 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 -2346 655174
rect -2966 654854 -2346 654938
rect -2966 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 -2346 654854
rect -2966 619174 -2346 654618
rect -2966 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 -2346 619174
rect -2966 618854 -2346 618938
rect -2966 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 -2346 618854
rect -2966 583174 -2346 618618
rect -2966 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 -2346 583174
rect -2966 582854 -2346 582938
rect -2966 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 -2346 582854
rect -2966 547174 -2346 582618
rect -2966 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 -2346 547174
rect -2966 546854 -2346 546938
rect -2966 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 -2346 546854
rect -2966 511174 -2346 546618
rect -2966 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 -2346 511174
rect -2966 510854 -2346 510938
rect -2966 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 -2346 510854
rect -2966 475174 -2346 510618
rect -2966 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 -2346 475174
rect -2966 474854 -2346 474938
rect -2966 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 -2346 474854
rect -2966 439174 -2346 474618
rect -2966 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 -2346 439174
rect -2966 438854 -2346 438938
rect -2966 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 -2346 438854
rect -2966 403174 -2346 438618
rect -2966 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 -2346 403174
rect -2966 402854 -2346 402938
rect -2966 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 -2346 402854
rect -2966 367174 -2346 402618
rect -2966 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 -2346 367174
rect -2966 366854 -2346 366938
rect -2966 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 -2346 366854
rect -2966 331174 -2346 366618
rect -2966 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 -2346 331174
rect -2966 330854 -2346 330938
rect -2966 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 -2346 330854
rect -2966 295174 -2346 330618
rect -2966 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 -2346 295174
rect -2966 294854 -2346 294938
rect -2966 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 -2346 294854
rect -2966 259174 -2346 294618
rect -2966 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 -2346 259174
rect -2966 258854 -2346 258938
rect -2966 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 -2346 258854
rect -2966 223174 -2346 258618
rect -2966 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 -2346 223174
rect -2966 222854 -2346 222938
rect -2966 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 -2346 222854
rect -2966 187174 -2346 222618
rect -2966 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 -2346 187174
rect -2966 186854 -2346 186938
rect -2966 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 -2346 186854
rect -2966 151174 -2346 186618
rect -2966 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 -2346 151174
rect -2966 150854 -2346 150938
rect -2966 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 -2346 150854
rect -2966 115174 -2346 150618
rect -2966 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 -2346 115174
rect -2966 114854 -2346 114938
rect -2966 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 -2346 114854
rect -2966 79174 -2346 114618
rect -2966 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 -2346 79174
rect -2966 78854 -2346 78938
rect -2966 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 -2346 78854
rect -2966 43174 -2346 78618
rect -2966 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 -2346 43174
rect -2966 42854 -2346 42938
rect -2966 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 -2346 42854
rect -2966 7174 -2346 42618
rect -2966 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 -2346 7174
rect -2966 6854 -2346 6938
rect -2966 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 -2346 6854
rect -2966 -1306 -2346 6618
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 5514 705798 6134 711590
rect 5514 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 6134 705798
rect 5514 705478 6134 705562
rect 5514 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 6134 705478
rect 5514 691174 6134 705242
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 3555 683364 3621 683365
rect 3555 683300 3556 683364
rect 3620 683300 3621 683364
rect 3555 683299 3621 683300
rect 3371 682956 3437 682957
rect 3371 682892 3372 682956
rect 3436 682892 3437 682956
rect 3371 682891 3437 682892
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 3374 606117 3434 682891
rect 3558 619173 3618 683299
rect 3739 683228 3805 683229
rect 3739 683164 3740 683228
rect 3804 683164 3805 683228
rect 3739 683163 3805 683164
rect 3742 671261 3802 683163
rect 3739 671260 3805 671261
rect 3739 671196 3740 671260
rect 3804 671196 3805 671260
rect 3739 671195 3805 671196
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 3555 619172 3621 619173
rect 3555 619108 3556 619172
rect 3620 619108 3621 619172
rect 3555 619107 3621 619108
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 3371 606116 3437 606117
rect 3371 606052 3372 606116
rect 3436 606052 3437 606116
rect 3371 606051 3437 606052
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 3371 136780 3437 136781
rect 3371 136716 3372 136780
rect 3436 136716 3437 136780
rect 3371 136715 3437 136716
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 3374 47021 3434 136715
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 3555 110668 3621 110669
rect 3555 110604 3556 110668
rect 3620 110604 3621 110668
rect 3555 110603 3621 110604
rect 3371 47020 3437 47021
rect 3371 46956 3372 47020
rect 3436 46956 3437 47020
rect 3371 46955 3437 46956
rect 3558 46885 3618 110603
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 3555 46884 3621 46885
rect 3555 46820 3556 46884
rect 3620 46820 3621 46884
rect 3555 46819 3621 46820
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect 5514 -1306 6134 6618
rect 5514 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 6134 -1306
rect 5514 -1626 6134 -1542
rect 5514 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 6134 -1626
rect 5514 -7654 6134 -1862
rect 9234 706758 9854 711590
rect 9234 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 9854 706758
rect 9234 706438 9854 706522
rect 9234 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 9854 706438
rect 9234 694894 9854 706202
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect 9234 -2266 9854 10338
rect 9234 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 9854 -2266
rect 9234 -2586 9854 -2502
rect 9234 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 9854 -2586
rect 9234 -7654 9854 -2822
rect 12954 707718 13574 711590
rect 12954 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 13574 707718
rect 12954 707398 13574 707482
rect 12954 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 13574 707398
rect 12954 698614 13574 707162
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect 12954 -3226 13574 14058
rect 12954 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 13574 -3226
rect 12954 -3546 13574 -3462
rect 12954 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 13574 -3546
rect 12954 -7654 13574 -3782
rect 16674 708678 17294 711590
rect 16674 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 17294 708678
rect 16674 708358 17294 708442
rect 16674 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 17294 708358
rect 16674 666334 17294 708122
rect 16674 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 17294 666334
rect 16674 666014 17294 666098
rect 16674 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 17294 666014
rect 16674 630334 17294 665778
rect 16674 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 17294 630334
rect 16674 630014 17294 630098
rect 16674 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 17294 630014
rect 16674 594334 17294 629778
rect 16674 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 17294 594334
rect 16674 594014 17294 594098
rect 16674 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 17294 594014
rect 16674 558334 17294 593778
rect 16674 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 17294 558334
rect 16674 558014 17294 558098
rect 16674 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 17294 558014
rect 16674 522334 17294 557778
rect 16674 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 17294 522334
rect 16674 522014 17294 522098
rect 16674 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 17294 522014
rect 16674 486334 17294 521778
rect 16674 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 17294 486334
rect 16674 486014 17294 486098
rect 16674 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 17294 486014
rect 16674 450334 17294 485778
rect 16674 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 17294 450334
rect 16674 450014 17294 450098
rect 16674 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 17294 450014
rect 16674 414334 17294 449778
rect 16674 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 17294 414334
rect 16674 414014 17294 414098
rect 16674 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 17294 414014
rect 16674 378334 17294 413778
rect 16674 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 17294 378334
rect 16674 378014 17294 378098
rect 16674 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 17294 378014
rect 16674 342334 17294 377778
rect 16674 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 17294 342334
rect 16674 342014 17294 342098
rect 16674 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 17294 342014
rect 16674 306334 17294 341778
rect 16674 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 17294 306334
rect 16674 306014 17294 306098
rect 16674 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 17294 306014
rect 16674 270334 17294 305778
rect 16674 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 17294 270334
rect 16674 270014 17294 270098
rect 16674 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 17294 270014
rect 16674 234334 17294 269778
rect 16674 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 17294 234334
rect 16674 234014 17294 234098
rect 16674 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 17294 234014
rect 16674 198334 17294 233778
rect 16674 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 17294 198334
rect 16674 198014 17294 198098
rect 16674 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 17294 198014
rect 16674 162334 17294 197778
rect 16674 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 17294 162334
rect 16674 162014 17294 162098
rect 16674 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 17294 162014
rect 16674 126334 17294 161778
rect 16674 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 17294 126334
rect 16674 126014 17294 126098
rect 16674 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 17294 126014
rect 16674 90334 17294 125778
rect 16674 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 17294 90334
rect 16674 90014 17294 90098
rect 16674 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 17294 90014
rect 16674 54334 17294 89778
rect 16674 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 17294 54334
rect 16674 54014 17294 54098
rect 16674 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 17294 54014
rect 16674 18334 17294 53778
rect 16674 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 17294 18334
rect 16674 18014 17294 18098
rect 16674 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 17294 18014
rect 16674 -4186 17294 17778
rect 16674 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 17294 -4186
rect 16674 -4506 17294 -4422
rect 16674 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 17294 -4506
rect 16674 -7654 17294 -4742
rect 20394 709638 21014 711590
rect 20394 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 21014 709638
rect 20394 709318 21014 709402
rect 20394 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 21014 709318
rect 20394 670054 21014 709082
rect 20394 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 21014 670054
rect 20394 669734 21014 669818
rect 20394 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 21014 669734
rect 20394 634054 21014 669498
rect 27834 711558 28454 711590
rect 27834 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 28454 711558
rect 27834 711238 28454 711322
rect 27834 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 28454 711238
rect 27834 677494 28454 711002
rect 27834 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 28454 677494
rect 27834 677174 28454 677258
rect 27834 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 28454 677174
rect 24208 651454 24528 651486
rect 24208 651218 24250 651454
rect 24486 651218 24528 651454
rect 24208 651134 24528 651218
rect 24208 650898 24250 651134
rect 24486 650898 24528 651134
rect 24208 650866 24528 650898
rect 20394 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 21014 634054
rect 20394 633734 21014 633818
rect 20394 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 21014 633734
rect 20394 598054 21014 633498
rect 27834 641494 28454 676938
rect 27834 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 28454 641494
rect 27834 641174 28454 641258
rect 27834 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 28454 641174
rect 24208 615454 24528 615486
rect 24208 615218 24250 615454
rect 24486 615218 24528 615454
rect 24208 615134 24528 615218
rect 24208 614898 24250 615134
rect 24486 614898 24528 615134
rect 24208 614866 24528 614898
rect 20394 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 21014 598054
rect 20394 597734 21014 597818
rect 20394 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 21014 597734
rect 20394 562054 21014 597498
rect 27834 605494 28454 640938
rect 27834 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 28454 605494
rect 27834 605174 28454 605258
rect 27834 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 28454 605174
rect 24208 579454 24528 579486
rect 24208 579218 24250 579454
rect 24486 579218 24528 579454
rect 24208 579134 24528 579218
rect 24208 578898 24250 579134
rect 24486 578898 24528 579134
rect 24208 578866 24528 578898
rect 20394 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 21014 562054
rect 20394 561734 21014 561818
rect 20394 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 21014 561734
rect 20394 526054 21014 561498
rect 27834 569494 28454 604938
rect 27834 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 28454 569494
rect 27834 569174 28454 569258
rect 27834 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 28454 569174
rect 24208 543454 24528 543486
rect 24208 543218 24250 543454
rect 24486 543218 24528 543454
rect 24208 543134 24528 543218
rect 24208 542898 24250 543134
rect 24486 542898 24528 543134
rect 24208 542866 24528 542898
rect 20394 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 21014 526054
rect 20394 525734 21014 525818
rect 20394 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 21014 525734
rect 20394 490054 21014 525498
rect 27834 533494 28454 568938
rect 27834 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 28454 533494
rect 27834 533174 28454 533258
rect 27834 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 28454 533174
rect 24208 507454 24528 507486
rect 24208 507218 24250 507454
rect 24486 507218 24528 507454
rect 24208 507134 24528 507218
rect 24208 506898 24250 507134
rect 24486 506898 24528 507134
rect 24208 506866 24528 506898
rect 20394 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 21014 490054
rect 20394 489734 21014 489818
rect 20394 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 21014 489734
rect 20394 454054 21014 489498
rect 27834 497494 28454 532938
rect 27834 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 28454 497494
rect 27834 497174 28454 497258
rect 27834 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 28454 497174
rect 24208 471454 24528 471486
rect 24208 471218 24250 471454
rect 24486 471218 24528 471454
rect 24208 471134 24528 471218
rect 24208 470898 24250 471134
rect 24486 470898 24528 471134
rect 24208 470866 24528 470898
rect 20394 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 21014 454054
rect 20394 453734 21014 453818
rect 20394 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 21014 453734
rect 20394 418054 21014 453498
rect 27834 461494 28454 496938
rect 27834 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 28454 461494
rect 27834 461174 28454 461258
rect 27834 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 28454 461174
rect 24208 435454 24528 435486
rect 24208 435218 24250 435454
rect 24486 435218 24528 435454
rect 24208 435134 24528 435218
rect 24208 434898 24250 435134
rect 24486 434898 24528 435134
rect 24208 434866 24528 434898
rect 20394 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 21014 418054
rect 20394 417734 21014 417818
rect 20394 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 21014 417734
rect 20394 382054 21014 417498
rect 27834 425494 28454 460938
rect 27834 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 28454 425494
rect 27834 425174 28454 425258
rect 27834 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 28454 425174
rect 24208 399454 24528 399486
rect 24208 399218 24250 399454
rect 24486 399218 24528 399454
rect 24208 399134 24528 399218
rect 24208 398898 24250 399134
rect 24486 398898 24528 399134
rect 24208 398866 24528 398898
rect 20394 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 21014 382054
rect 20394 381734 21014 381818
rect 20394 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 21014 381734
rect 20394 346054 21014 381498
rect 27834 389494 28454 424938
rect 27834 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 28454 389494
rect 27834 389174 28454 389258
rect 27834 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 28454 389174
rect 24208 363454 24528 363486
rect 24208 363218 24250 363454
rect 24486 363218 24528 363454
rect 24208 363134 24528 363218
rect 24208 362898 24250 363134
rect 24486 362898 24528 363134
rect 24208 362866 24528 362898
rect 20394 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 21014 346054
rect 20394 345734 21014 345818
rect 20394 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 21014 345734
rect 20394 310054 21014 345498
rect 27834 353494 28454 388938
rect 27834 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 28454 353494
rect 27834 353174 28454 353258
rect 27834 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 28454 353174
rect 24208 327454 24528 327486
rect 24208 327218 24250 327454
rect 24486 327218 24528 327454
rect 24208 327134 24528 327218
rect 24208 326898 24250 327134
rect 24486 326898 24528 327134
rect 24208 326866 24528 326898
rect 20394 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 21014 310054
rect 20394 309734 21014 309818
rect 20394 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 21014 309734
rect 20394 274054 21014 309498
rect 27834 317494 28454 352938
rect 27834 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 28454 317494
rect 27834 317174 28454 317258
rect 27834 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 28454 317174
rect 24208 291454 24528 291486
rect 24208 291218 24250 291454
rect 24486 291218 24528 291454
rect 24208 291134 24528 291218
rect 24208 290898 24250 291134
rect 24486 290898 24528 291134
rect 24208 290866 24528 290898
rect 20394 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 21014 274054
rect 20394 273734 21014 273818
rect 20394 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 21014 273734
rect 20394 238054 21014 273498
rect 27834 281494 28454 316938
rect 27834 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 28454 281494
rect 27834 281174 28454 281258
rect 27834 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 28454 281174
rect 24208 255454 24528 255486
rect 24208 255218 24250 255454
rect 24486 255218 24528 255454
rect 24208 255134 24528 255218
rect 24208 254898 24250 255134
rect 24486 254898 24528 255134
rect 24208 254866 24528 254898
rect 20394 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 21014 238054
rect 20394 237734 21014 237818
rect 20394 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 21014 237734
rect 20394 202054 21014 237498
rect 27834 245494 28454 280938
rect 27834 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 28454 245494
rect 27834 245174 28454 245258
rect 27834 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 28454 245174
rect 24208 219454 24528 219486
rect 24208 219218 24250 219454
rect 24486 219218 24528 219454
rect 24208 219134 24528 219218
rect 24208 218898 24250 219134
rect 24486 218898 24528 219134
rect 24208 218866 24528 218898
rect 20394 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 21014 202054
rect 20394 201734 21014 201818
rect 20394 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 21014 201734
rect 20394 166054 21014 201498
rect 27834 209494 28454 244938
rect 27834 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 28454 209494
rect 27834 209174 28454 209258
rect 27834 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 28454 209174
rect 24208 183454 24528 183486
rect 24208 183218 24250 183454
rect 24486 183218 24528 183454
rect 24208 183134 24528 183218
rect 24208 182898 24250 183134
rect 24486 182898 24528 183134
rect 24208 182866 24528 182898
rect 20394 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 21014 166054
rect 20394 165734 21014 165818
rect 20394 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 21014 165734
rect 20394 130054 21014 165498
rect 27834 173494 28454 208938
rect 27834 173258 27866 173494
rect 28102 173258 28186 173494
rect 28422 173258 28454 173494
rect 27834 173174 28454 173258
rect 27834 172938 27866 173174
rect 28102 172938 28186 173174
rect 28422 172938 28454 173174
rect 24208 147454 24528 147486
rect 24208 147218 24250 147454
rect 24486 147218 24528 147454
rect 24208 147134 24528 147218
rect 24208 146898 24250 147134
rect 24486 146898 24528 147134
rect 24208 146866 24528 146898
rect 20394 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 21014 130054
rect 20394 129734 21014 129818
rect 20394 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 21014 129734
rect 20394 94054 21014 129498
rect 27834 137494 28454 172938
rect 27834 137258 27866 137494
rect 28102 137258 28186 137494
rect 28422 137258 28454 137494
rect 27834 137174 28454 137258
rect 27834 136938 27866 137174
rect 28102 136938 28186 137174
rect 28422 136938 28454 137174
rect 24208 111454 24528 111486
rect 24208 111218 24250 111454
rect 24486 111218 24528 111454
rect 24208 111134 24528 111218
rect 24208 110898 24250 111134
rect 24486 110898 24528 111134
rect 24208 110866 24528 110898
rect 20394 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 21014 94054
rect 20394 93734 21014 93818
rect 20394 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 21014 93734
rect 20394 58054 21014 93498
rect 27834 101494 28454 136938
rect 27834 101258 27866 101494
rect 28102 101258 28186 101494
rect 28422 101258 28454 101494
rect 27834 101174 28454 101258
rect 27834 100938 27866 101174
rect 28102 100938 28186 101174
rect 28422 100938 28454 101174
rect 24208 75454 24528 75486
rect 24208 75218 24250 75454
rect 24486 75218 24528 75454
rect 24208 75134 24528 75218
rect 24208 74898 24250 75134
rect 24486 74898 24528 75134
rect 24208 74866 24528 74898
rect 27834 65494 28454 100938
rect 27834 65258 27866 65494
rect 28102 65258 28186 65494
rect 28422 65258 28454 65494
rect 27834 65174 28454 65258
rect 27834 64938 27866 65174
rect 28102 64938 28186 65174
rect 28422 64938 28454 65174
rect 22691 59940 22757 59941
rect 22691 59876 22692 59940
rect 22756 59876 22757 59940
rect 22691 59875 22757 59876
rect 20394 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 21014 58054
rect 20394 57734 21014 57818
rect 20394 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 21014 57734
rect 20394 22054 21014 57498
rect 22139 49604 22205 49605
rect 22139 49540 22140 49604
rect 22204 49540 22205 49604
rect 22139 49539 22205 49540
rect 22142 46477 22202 49539
rect 22694 46613 22754 59875
rect 22691 46612 22757 46613
rect 22691 46548 22692 46612
rect 22756 46548 22757 46612
rect 22691 46547 22757 46548
rect 22139 46476 22205 46477
rect 22139 46412 22140 46476
rect 22204 46412 22205 46476
rect 22139 46411 22205 46412
rect 20394 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 21014 22054
rect 20394 21734 21014 21818
rect 20394 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 21014 21734
rect 20394 -5146 21014 21498
rect 20394 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 21014 -5146
rect 20394 -5466 21014 -5382
rect 20394 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 21014 -5466
rect 20394 -7654 21014 -5702
rect 24114 25774 24734 45068
rect 24114 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 24734 25774
rect 24114 25454 24734 25538
rect 24114 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 24734 25454
rect 24114 -6106 24734 25218
rect 24114 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 24734 -6106
rect 24114 -6426 24734 -6342
rect 24114 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 24734 -6426
rect 24114 -7654 24734 -6662
rect 27834 29494 28454 64938
rect 27834 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 28454 29494
rect 27834 29174 28454 29258
rect 27834 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 28454 29174
rect 27834 -7066 28454 28938
rect 27834 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 28454 -7066
rect 27834 -7386 28454 -7302
rect 27834 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 28454 -7386
rect 27834 -7654 28454 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 41514 705798 42134 711590
rect 41514 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 42134 705798
rect 41514 705478 42134 705562
rect 41514 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 42134 705478
rect 41514 691174 42134 705242
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 39568 655174 39888 655206
rect 39568 654938 39610 655174
rect 39846 654938 39888 655174
rect 39568 654854 39888 654938
rect 39568 654618 39610 654854
rect 39846 654618 39888 654854
rect 39568 654586 39888 654618
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 39568 619174 39888 619206
rect 39568 618938 39610 619174
rect 39846 618938 39888 619174
rect 39568 618854 39888 618938
rect 39568 618618 39610 618854
rect 39846 618618 39888 618854
rect 39568 618586 39888 618618
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 39568 583174 39888 583206
rect 39568 582938 39610 583174
rect 39846 582938 39888 583174
rect 39568 582854 39888 582938
rect 39568 582618 39610 582854
rect 39846 582618 39888 582854
rect 39568 582586 39888 582618
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 39568 547174 39888 547206
rect 39568 546938 39610 547174
rect 39846 546938 39888 547174
rect 39568 546854 39888 546938
rect 39568 546618 39610 546854
rect 39846 546618 39888 546854
rect 39568 546586 39888 546618
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 39568 511174 39888 511206
rect 39568 510938 39610 511174
rect 39846 510938 39888 511174
rect 39568 510854 39888 510938
rect 39568 510618 39610 510854
rect 39846 510618 39888 510854
rect 39568 510586 39888 510618
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 39568 475174 39888 475206
rect 39568 474938 39610 475174
rect 39846 474938 39888 475174
rect 39568 474854 39888 474938
rect 39568 474618 39610 474854
rect 39846 474618 39888 474854
rect 39568 474586 39888 474618
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 39568 439174 39888 439206
rect 39568 438938 39610 439174
rect 39846 438938 39888 439174
rect 39568 438854 39888 438938
rect 39568 438618 39610 438854
rect 39846 438618 39888 438854
rect 39568 438586 39888 438618
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 39568 403174 39888 403206
rect 39568 402938 39610 403174
rect 39846 402938 39888 403174
rect 39568 402854 39888 402938
rect 39568 402618 39610 402854
rect 39846 402618 39888 402854
rect 39568 402586 39888 402618
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 39568 367174 39888 367206
rect 39568 366938 39610 367174
rect 39846 366938 39888 367174
rect 39568 366854 39888 366938
rect 39568 366618 39610 366854
rect 39846 366618 39888 366854
rect 39568 366586 39888 366618
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 39568 331174 39888 331206
rect 39568 330938 39610 331174
rect 39846 330938 39888 331174
rect 39568 330854 39888 330938
rect 39568 330618 39610 330854
rect 39846 330618 39888 330854
rect 39568 330586 39888 330618
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 39568 295174 39888 295206
rect 39568 294938 39610 295174
rect 39846 294938 39888 295174
rect 39568 294854 39888 294938
rect 39568 294618 39610 294854
rect 39846 294618 39888 294854
rect 39568 294586 39888 294618
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 39568 259174 39888 259206
rect 39568 258938 39610 259174
rect 39846 258938 39888 259174
rect 39568 258854 39888 258938
rect 39568 258618 39610 258854
rect 39846 258618 39888 258854
rect 39568 258586 39888 258618
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 39568 223174 39888 223206
rect 39568 222938 39610 223174
rect 39846 222938 39888 223174
rect 39568 222854 39888 222938
rect 39568 222618 39610 222854
rect 39846 222618 39888 222854
rect 39568 222586 39888 222618
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 39568 187174 39888 187206
rect 39568 186938 39610 187174
rect 39846 186938 39888 187174
rect 39568 186854 39888 186938
rect 39568 186618 39610 186854
rect 39846 186618 39888 186854
rect 39568 186586 39888 186618
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 39568 151174 39888 151206
rect 39568 150938 39610 151174
rect 39846 150938 39888 151174
rect 39568 150854 39888 150938
rect 39568 150618 39610 150854
rect 39846 150618 39888 150854
rect 39568 150586 39888 150618
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 39568 115174 39888 115206
rect 39568 114938 39610 115174
rect 39846 114938 39888 115174
rect 39568 114854 39888 114938
rect 39568 114618 39610 114854
rect 39846 114618 39888 114854
rect 39568 114586 39888 114618
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 39568 79174 39888 79206
rect 39568 78938 39610 79174
rect 39846 78938 39888 79174
rect 39568 78854 39888 78938
rect 39568 78618 39610 78854
rect 39846 78618 39888 78854
rect 39568 78586 39888 78618
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -1306 42134 6618
rect 41514 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 42134 -1306
rect 41514 -1626 42134 -1542
rect 41514 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 42134 -1626
rect 41514 -7654 42134 -1862
rect 45234 706758 45854 711590
rect 45234 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 45854 706758
rect 45234 706438 45854 706522
rect 45234 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 45854 706438
rect 45234 694894 45854 706202
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -2266 45854 10338
rect 45234 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 45854 -2266
rect 45234 -2586 45854 -2502
rect 45234 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 45854 -2586
rect 45234 -7654 45854 -2822
rect 48954 707718 49574 711590
rect 48954 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 49574 707718
rect 48954 707398 49574 707482
rect 48954 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 49574 707398
rect 48954 698614 49574 707162
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 680513 74414 686898
rect 77514 705798 78134 711590
rect 77514 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 78134 705798
rect 77514 705478 78134 705562
rect 77514 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 78134 705478
rect 77514 691174 78134 705242
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 680513 78134 690618
rect 81234 706758 81854 711590
rect 81234 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 81854 706758
rect 81234 706438 81854 706522
rect 81234 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 81854 706438
rect 81234 694894 81854 706202
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 680513 81854 694338
rect 84954 707718 85574 711590
rect 84954 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 85574 707718
rect 84954 707398 85574 707482
rect 84954 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 85574 707398
rect 84954 698614 85574 707162
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 680513 85574 698058
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 680513 110414 686898
rect 113514 705798 114134 711590
rect 113514 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 114134 705798
rect 113514 705478 114134 705562
rect 113514 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 114134 705478
rect 113514 691174 114134 705242
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 680513 114134 690618
rect 117234 706758 117854 711590
rect 117234 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 117854 706758
rect 117234 706438 117854 706522
rect 117234 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 117854 706438
rect 117234 694894 117854 706202
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 680513 117854 694338
rect 120954 707718 121574 711590
rect 120954 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 121574 707718
rect 120954 707398 121574 707482
rect 120954 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 121574 707398
rect 120954 698614 121574 707162
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 680513 121574 698058
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 680513 146414 686898
rect 149514 705798 150134 711590
rect 149514 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 150134 705798
rect 149514 705478 150134 705562
rect 149514 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 150134 705478
rect 149514 691174 150134 705242
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 680513 150134 690618
rect 153234 706758 153854 711590
rect 153234 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 153854 706758
rect 153234 706438 153854 706522
rect 153234 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 153854 706438
rect 153234 694894 153854 706202
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 680513 153854 694338
rect 156954 707718 157574 711590
rect 156954 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 157574 707718
rect 156954 707398 157574 707482
rect 156954 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 157574 707398
rect 156954 698614 157574 707162
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 680513 157574 698058
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 680513 182414 686898
rect 185514 705798 186134 711590
rect 185514 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 186134 705798
rect 185514 705478 186134 705562
rect 185514 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 186134 705478
rect 185514 691174 186134 705242
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 680513 186134 690618
rect 189234 706758 189854 711590
rect 189234 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 189854 706758
rect 189234 706438 189854 706522
rect 189234 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 189854 706438
rect 189234 694894 189854 706202
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 680513 189854 694338
rect 192954 707718 193574 711590
rect 192954 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 193574 707718
rect 192954 707398 193574 707482
rect 192954 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 193574 707398
rect 192954 698614 193574 707162
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 684676 193574 698058
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 680513 218414 686898
rect 221514 705798 222134 711590
rect 221514 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 222134 705798
rect 221514 705478 222134 705562
rect 221514 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 222134 705478
rect 221514 691174 222134 705242
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 680513 222134 690618
rect 225234 706758 225854 711590
rect 225234 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 225854 706758
rect 225234 706438 225854 706522
rect 225234 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 225854 706438
rect 225234 694894 225854 706202
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 680513 225854 694338
rect 228954 707718 229574 711590
rect 228954 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 229574 707718
rect 228954 707398 229574 707482
rect 228954 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 229574 707398
rect 228954 698614 229574 707162
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 680513 229574 698058
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 680513 254414 686898
rect 257514 705798 258134 711590
rect 257514 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 258134 705798
rect 257514 705478 258134 705562
rect 257514 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 258134 705478
rect 257514 691174 258134 705242
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 680513 258134 690618
rect 261234 706758 261854 711590
rect 261234 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 261854 706758
rect 261234 706438 261854 706522
rect 261234 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 261854 706438
rect 261234 694894 261854 706202
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 680513 261854 694338
rect 264954 707718 265574 711590
rect 264954 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 265574 707718
rect 264954 707398 265574 707482
rect 264954 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 265574 707398
rect 264954 698614 265574 707162
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 680513 265574 698058
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 680513 290414 686898
rect 293514 705798 294134 711590
rect 293514 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 294134 705798
rect 293514 705478 294134 705562
rect 293514 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 294134 705478
rect 293514 691174 294134 705242
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 680513 294134 690618
rect 297234 706758 297854 711590
rect 297234 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 297854 706758
rect 297234 706438 297854 706522
rect 297234 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 297854 706438
rect 297234 694894 297854 706202
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 680513 297854 694338
rect 300954 707718 301574 711590
rect 300954 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 301574 707718
rect 300954 707398 301574 707482
rect 300954 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 301574 707398
rect 300954 698614 301574 707162
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 684676 301574 698058
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 680513 326414 686898
rect 329514 705798 330134 711590
rect 329514 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 330134 705798
rect 329514 705478 330134 705562
rect 329514 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 330134 705478
rect 329514 691174 330134 705242
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 680513 330134 690618
rect 333234 706758 333854 711590
rect 333234 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 333854 706758
rect 333234 706438 333854 706522
rect 333234 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 333854 706438
rect 333234 694894 333854 706202
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 680513 333854 694338
rect 336954 707718 337574 711590
rect 336954 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 337574 707718
rect 336954 707398 337574 707482
rect 336954 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 337574 707398
rect 336954 698614 337574 707162
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 680513 337574 698058
rect 344394 709638 345014 711590
rect 344394 709402 344426 709638
rect 344662 709402 344746 709638
rect 344982 709402 345014 709638
rect 344394 709318 345014 709402
rect 344394 709082 344426 709318
rect 344662 709082 344746 709318
rect 344982 709082 345014 709318
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 344394 670054 345014 709082
rect 344394 669818 344426 670054
rect 344662 669818 344746 670054
rect 344982 669818 345014 670054
rect 344394 669734 345014 669818
rect 344394 669498 344426 669734
rect 344662 669498 344746 669734
rect 344982 669498 345014 669734
rect 70288 655174 70608 655206
rect 70288 654938 70330 655174
rect 70566 654938 70608 655174
rect 70288 654854 70608 654938
rect 70288 654618 70330 654854
rect 70566 654618 70608 654854
rect 70288 654586 70608 654618
rect 101008 655174 101328 655206
rect 101008 654938 101050 655174
rect 101286 654938 101328 655174
rect 101008 654854 101328 654938
rect 101008 654618 101050 654854
rect 101286 654618 101328 654854
rect 101008 654586 101328 654618
rect 131728 655174 132048 655206
rect 131728 654938 131770 655174
rect 132006 654938 132048 655174
rect 131728 654854 132048 654938
rect 131728 654618 131770 654854
rect 132006 654618 132048 654854
rect 131728 654586 132048 654618
rect 162448 655174 162768 655206
rect 162448 654938 162490 655174
rect 162726 654938 162768 655174
rect 162448 654854 162768 654938
rect 162448 654618 162490 654854
rect 162726 654618 162768 654854
rect 162448 654586 162768 654618
rect 193168 655174 193488 655206
rect 193168 654938 193210 655174
rect 193446 654938 193488 655174
rect 193168 654854 193488 654938
rect 193168 654618 193210 654854
rect 193446 654618 193488 654854
rect 193168 654586 193488 654618
rect 223888 655174 224208 655206
rect 223888 654938 223930 655174
rect 224166 654938 224208 655174
rect 223888 654854 224208 654938
rect 223888 654618 223930 654854
rect 224166 654618 224208 654854
rect 223888 654586 224208 654618
rect 254608 655174 254928 655206
rect 254608 654938 254650 655174
rect 254886 654938 254928 655174
rect 254608 654854 254928 654938
rect 254608 654618 254650 654854
rect 254886 654618 254928 654854
rect 254608 654586 254928 654618
rect 285328 655174 285648 655206
rect 285328 654938 285370 655174
rect 285606 654938 285648 655174
rect 285328 654854 285648 654938
rect 285328 654618 285370 654854
rect 285606 654618 285648 654854
rect 285328 654586 285648 654618
rect 316048 655174 316368 655206
rect 316048 654938 316090 655174
rect 316326 654938 316368 655174
rect 316048 654854 316368 654938
rect 316048 654618 316090 654854
rect 316326 654618 316368 654854
rect 316048 654586 316368 654618
rect 54928 651454 55248 651486
rect 54928 651218 54970 651454
rect 55206 651218 55248 651454
rect 54928 651134 55248 651218
rect 54928 650898 54970 651134
rect 55206 650898 55248 651134
rect 54928 650866 55248 650898
rect 85648 651454 85968 651486
rect 85648 651218 85690 651454
rect 85926 651218 85968 651454
rect 85648 651134 85968 651218
rect 85648 650898 85690 651134
rect 85926 650898 85968 651134
rect 85648 650866 85968 650898
rect 116368 651454 116688 651486
rect 116368 651218 116410 651454
rect 116646 651218 116688 651454
rect 116368 651134 116688 651218
rect 116368 650898 116410 651134
rect 116646 650898 116688 651134
rect 116368 650866 116688 650898
rect 147088 651454 147408 651486
rect 147088 651218 147130 651454
rect 147366 651218 147408 651454
rect 147088 651134 147408 651218
rect 147088 650898 147130 651134
rect 147366 650898 147408 651134
rect 147088 650866 147408 650898
rect 177808 651454 178128 651486
rect 177808 651218 177850 651454
rect 178086 651218 178128 651454
rect 177808 651134 178128 651218
rect 177808 650898 177850 651134
rect 178086 650898 178128 651134
rect 177808 650866 178128 650898
rect 208528 651454 208848 651486
rect 208528 651218 208570 651454
rect 208806 651218 208848 651454
rect 208528 651134 208848 651218
rect 208528 650898 208570 651134
rect 208806 650898 208848 651134
rect 208528 650866 208848 650898
rect 239248 651454 239568 651486
rect 239248 651218 239290 651454
rect 239526 651218 239568 651454
rect 239248 651134 239568 651218
rect 239248 650898 239290 651134
rect 239526 650898 239568 651134
rect 239248 650866 239568 650898
rect 269968 651454 270288 651486
rect 269968 651218 270010 651454
rect 270246 651218 270288 651454
rect 269968 651134 270288 651218
rect 269968 650898 270010 651134
rect 270246 650898 270288 651134
rect 269968 650866 270288 650898
rect 300688 651454 301008 651486
rect 300688 651218 300730 651454
rect 300966 651218 301008 651454
rect 300688 651134 301008 651218
rect 300688 650898 300730 651134
rect 300966 650898 301008 651134
rect 300688 650866 301008 650898
rect 331408 651454 331728 651486
rect 331408 651218 331450 651454
rect 331686 651218 331728 651454
rect 331408 651134 331728 651218
rect 331408 650898 331450 651134
rect 331686 650898 331728 651134
rect 331408 650866 331728 650898
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 344394 634054 345014 669498
rect 348114 710598 348734 711590
rect 348114 710362 348146 710598
rect 348382 710362 348466 710598
rect 348702 710362 348734 710598
rect 348114 710278 348734 710362
rect 348114 710042 348146 710278
rect 348382 710042 348466 710278
rect 348702 710042 348734 710278
rect 348114 673774 348734 710042
rect 348114 673538 348146 673774
rect 348382 673538 348466 673774
rect 348702 673538 348734 673774
rect 348114 673454 348734 673538
rect 348114 673218 348146 673454
rect 348382 673218 348466 673454
rect 348702 673218 348734 673454
rect 346768 655174 347088 655206
rect 346768 654938 346810 655174
rect 347046 654938 347088 655174
rect 346768 654854 347088 654938
rect 346768 654618 346810 654854
rect 347046 654618 347088 654854
rect 346768 654586 347088 654618
rect 344394 633818 344426 634054
rect 344662 633818 344746 634054
rect 344982 633818 345014 634054
rect 344394 633734 345014 633818
rect 344394 633498 344426 633734
rect 344662 633498 344746 633734
rect 344982 633498 345014 633734
rect 70288 619174 70608 619206
rect 70288 618938 70330 619174
rect 70566 618938 70608 619174
rect 70288 618854 70608 618938
rect 70288 618618 70330 618854
rect 70566 618618 70608 618854
rect 70288 618586 70608 618618
rect 101008 619174 101328 619206
rect 101008 618938 101050 619174
rect 101286 618938 101328 619174
rect 101008 618854 101328 618938
rect 101008 618618 101050 618854
rect 101286 618618 101328 618854
rect 101008 618586 101328 618618
rect 131728 619174 132048 619206
rect 131728 618938 131770 619174
rect 132006 618938 132048 619174
rect 131728 618854 132048 618938
rect 131728 618618 131770 618854
rect 132006 618618 132048 618854
rect 131728 618586 132048 618618
rect 162448 619174 162768 619206
rect 162448 618938 162490 619174
rect 162726 618938 162768 619174
rect 162448 618854 162768 618938
rect 162448 618618 162490 618854
rect 162726 618618 162768 618854
rect 162448 618586 162768 618618
rect 193168 619174 193488 619206
rect 193168 618938 193210 619174
rect 193446 618938 193488 619174
rect 193168 618854 193488 618938
rect 193168 618618 193210 618854
rect 193446 618618 193488 618854
rect 193168 618586 193488 618618
rect 223888 619174 224208 619206
rect 223888 618938 223930 619174
rect 224166 618938 224208 619174
rect 223888 618854 224208 618938
rect 223888 618618 223930 618854
rect 224166 618618 224208 618854
rect 223888 618586 224208 618618
rect 254608 619174 254928 619206
rect 254608 618938 254650 619174
rect 254886 618938 254928 619174
rect 254608 618854 254928 618938
rect 254608 618618 254650 618854
rect 254886 618618 254928 618854
rect 254608 618586 254928 618618
rect 285328 619174 285648 619206
rect 285328 618938 285370 619174
rect 285606 618938 285648 619174
rect 285328 618854 285648 618938
rect 285328 618618 285370 618854
rect 285606 618618 285648 618854
rect 285328 618586 285648 618618
rect 316048 619174 316368 619206
rect 316048 618938 316090 619174
rect 316326 618938 316368 619174
rect 316048 618854 316368 618938
rect 316048 618618 316090 618854
rect 316326 618618 316368 618854
rect 316048 618586 316368 618618
rect 54928 615454 55248 615486
rect 54928 615218 54970 615454
rect 55206 615218 55248 615454
rect 54928 615134 55248 615218
rect 54928 614898 54970 615134
rect 55206 614898 55248 615134
rect 54928 614866 55248 614898
rect 85648 615454 85968 615486
rect 85648 615218 85690 615454
rect 85926 615218 85968 615454
rect 85648 615134 85968 615218
rect 85648 614898 85690 615134
rect 85926 614898 85968 615134
rect 85648 614866 85968 614898
rect 116368 615454 116688 615486
rect 116368 615218 116410 615454
rect 116646 615218 116688 615454
rect 116368 615134 116688 615218
rect 116368 614898 116410 615134
rect 116646 614898 116688 615134
rect 116368 614866 116688 614898
rect 147088 615454 147408 615486
rect 147088 615218 147130 615454
rect 147366 615218 147408 615454
rect 147088 615134 147408 615218
rect 147088 614898 147130 615134
rect 147366 614898 147408 615134
rect 147088 614866 147408 614898
rect 177808 615454 178128 615486
rect 177808 615218 177850 615454
rect 178086 615218 178128 615454
rect 177808 615134 178128 615218
rect 177808 614898 177850 615134
rect 178086 614898 178128 615134
rect 177808 614866 178128 614898
rect 208528 615454 208848 615486
rect 208528 615218 208570 615454
rect 208806 615218 208848 615454
rect 208528 615134 208848 615218
rect 208528 614898 208570 615134
rect 208806 614898 208848 615134
rect 208528 614866 208848 614898
rect 239248 615454 239568 615486
rect 239248 615218 239290 615454
rect 239526 615218 239568 615454
rect 239248 615134 239568 615218
rect 239248 614898 239290 615134
rect 239526 614898 239568 615134
rect 239248 614866 239568 614898
rect 269968 615454 270288 615486
rect 269968 615218 270010 615454
rect 270246 615218 270288 615454
rect 269968 615134 270288 615218
rect 269968 614898 270010 615134
rect 270246 614898 270288 615134
rect 269968 614866 270288 614898
rect 300688 615454 301008 615486
rect 300688 615218 300730 615454
rect 300966 615218 301008 615454
rect 300688 615134 301008 615218
rect 300688 614898 300730 615134
rect 300966 614898 301008 615134
rect 300688 614866 301008 614898
rect 331408 615454 331728 615486
rect 331408 615218 331450 615454
rect 331686 615218 331728 615454
rect 331408 615134 331728 615218
rect 331408 614898 331450 615134
rect 331686 614898 331728 615134
rect 331408 614866 331728 614898
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 344394 598054 345014 633498
rect 348114 637774 348734 673218
rect 348114 637538 348146 637774
rect 348382 637538 348466 637774
rect 348702 637538 348734 637774
rect 348114 637454 348734 637538
rect 348114 637218 348146 637454
rect 348382 637218 348466 637454
rect 348702 637218 348734 637454
rect 346768 619174 347088 619206
rect 346768 618938 346810 619174
rect 347046 618938 347088 619174
rect 346768 618854 347088 618938
rect 346768 618618 346810 618854
rect 347046 618618 347088 618854
rect 346768 618586 347088 618618
rect 344394 597818 344426 598054
rect 344662 597818 344746 598054
rect 344982 597818 345014 598054
rect 344394 597734 345014 597818
rect 344394 597498 344426 597734
rect 344662 597498 344746 597734
rect 344982 597498 345014 597734
rect 70288 583174 70608 583206
rect 70288 582938 70330 583174
rect 70566 582938 70608 583174
rect 70288 582854 70608 582938
rect 70288 582618 70330 582854
rect 70566 582618 70608 582854
rect 70288 582586 70608 582618
rect 101008 583174 101328 583206
rect 101008 582938 101050 583174
rect 101286 582938 101328 583174
rect 101008 582854 101328 582938
rect 101008 582618 101050 582854
rect 101286 582618 101328 582854
rect 101008 582586 101328 582618
rect 131728 583174 132048 583206
rect 131728 582938 131770 583174
rect 132006 582938 132048 583174
rect 131728 582854 132048 582938
rect 131728 582618 131770 582854
rect 132006 582618 132048 582854
rect 131728 582586 132048 582618
rect 162448 583174 162768 583206
rect 162448 582938 162490 583174
rect 162726 582938 162768 583174
rect 162448 582854 162768 582938
rect 162448 582618 162490 582854
rect 162726 582618 162768 582854
rect 162448 582586 162768 582618
rect 193168 583174 193488 583206
rect 193168 582938 193210 583174
rect 193446 582938 193488 583174
rect 193168 582854 193488 582938
rect 193168 582618 193210 582854
rect 193446 582618 193488 582854
rect 193168 582586 193488 582618
rect 223888 583174 224208 583206
rect 223888 582938 223930 583174
rect 224166 582938 224208 583174
rect 223888 582854 224208 582938
rect 223888 582618 223930 582854
rect 224166 582618 224208 582854
rect 223888 582586 224208 582618
rect 254608 583174 254928 583206
rect 254608 582938 254650 583174
rect 254886 582938 254928 583174
rect 254608 582854 254928 582938
rect 254608 582618 254650 582854
rect 254886 582618 254928 582854
rect 254608 582586 254928 582618
rect 285328 583174 285648 583206
rect 285328 582938 285370 583174
rect 285606 582938 285648 583174
rect 285328 582854 285648 582938
rect 285328 582618 285370 582854
rect 285606 582618 285648 582854
rect 285328 582586 285648 582618
rect 316048 583174 316368 583206
rect 316048 582938 316090 583174
rect 316326 582938 316368 583174
rect 316048 582854 316368 582938
rect 316048 582618 316090 582854
rect 316326 582618 316368 582854
rect 316048 582586 316368 582618
rect 54928 579454 55248 579486
rect 54928 579218 54970 579454
rect 55206 579218 55248 579454
rect 54928 579134 55248 579218
rect 54928 578898 54970 579134
rect 55206 578898 55248 579134
rect 54928 578866 55248 578898
rect 85648 579454 85968 579486
rect 85648 579218 85690 579454
rect 85926 579218 85968 579454
rect 85648 579134 85968 579218
rect 85648 578898 85690 579134
rect 85926 578898 85968 579134
rect 85648 578866 85968 578898
rect 116368 579454 116688 579486
rect 116368 579218 116410 579454
rect 116646 579218 116688 579454
rect 116368 579134 116688 579218
rect 116368 578898 116410 579134
rect 116646 578898 116688 579134
rect 116368 578866 116688 578898
rect 147088 579454 147408 579486
rect 147088 579218 147130 579454
rect 147366 579218 147408 579454
rect 147088 579134 147408 579218
rect 147088 578898 147130 579134
rect 147366 578898 147408 579134
rect 147088 578866 147408 578898
rect 177808 579454 178128 579486
rect 177808 579218 177850 579454
rect 178086 579218 178128 579454
rect 177808 579134 178128 579218
rect 177808 578898 177850 579134
rect 178086 578898 178128 579134
rect 177808 578866 178128 578898
rect 208528 579454 208848 579486
rect 208528 579218 208570 579454
rect 208806 579218 208848 579454
rect 208528 579134 208848 579218
rect 208528 578898 208570 579134
rect 208806 578898 208848 579134
rect 208528 578866 208848 578898
rect 239248 579454 239568 579486
rect 239248 579218 239290 579454
rect 239526 579218 239568 579454
rect 239248 579134 239568 579218
rect 239248 578898 239290 579134
rect 239526 578898 239568 579134
rect 239248 578866 239568 578898
rect 269968 579454 270288 579486
rect 269968 579218 270010 579454
rect 270246 579218 270288 579454
rect 269968 579134 270288 579218
rect 269968 578898 270010 579134
rect 270246 578898 270288 579134
rect 269968 578866 270288 578898
rect 300688 579454 301008 579486
rect 300688 579218 300730 579454
rect 300966 579218 301008 579454
rect 300688 579134 301008 579218
rect 300688 578898 300730 579134
rect 300966 578898 301008 579134
rect 300688 578866 301008 578898
rect 331408 579454 331728 579486
rect 331408 579218 331450 579454
rect 331686 579218 331728 579454
rect 331408 579134 331728 579218
rect 331408 578898 331450 579134
rect 331686 578898 331728 579134
rect 331408 578866 331728 578898
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 344394 562054 345014 597498
rect 348114 601774 348734 637218
rect 348114 601538 348146 601774
rect 348382 601538 348466 601774
rect 348702 601538 348734 601774
rect 348114 601454 348734 601538
rect 348114 601218 348146 601454
rect 348382 601218 348466 601454
rect 348702 601218 348734 601454
rect 346768 583174 347088 583206
rect 346768 582938 346810 583174
rect 347046 582938 347088 583174
rect 346768 582854 347088 582938
rect 346768 582618 346810 582854
rect 347046 582618 347088 582854
rect 346768 582586 347088 582618
rect 344394 561818 344426 562054
rect 344662 561818 344746 562054
rect 344982 561818 345014 562054
rect 344394 561734 345014 561818
rect 344394 561498 344426 561734
rect 344662 561498 344746 561734
rect 344982 561498 345014 561734
rect 70288 547174 70608 547206
rect 70288 546938 70330 547174
rect 70566 546938 70608 547174
rect 70288 546854 70608 546938
rect 70288 546618 70330 546854
rect 70566 546618 70608 546854
rect 70288 546586 70608 546618
rect 101008 547174 101328 547206
rect 101008 546938 101050 547174
rect 101286 546938 101328 547174
rect 101008 546854 101328 546938
rect 101008 546618 101050 546854
rect 101286 546618 101328 546854
rect 101008 546586 101328 546618
rect 131728 547174 132048 547206
rect 131728 546938 131770 547174
rect 132006 546938 132048 547174
rect 131728 546854 132048 546938
rect 131728 546618 131770 546854
rect 132006 546618 132048 546854
rect 131728 546586 132048 546618
rect 162448 547174 162768 547206
rect 162448 546938 162490 547174
rect 162726 546938 162768 547174
rect 162448 546854 162768 546938
rect 162448 546618 162490 546854
rect 162726 546618 162768 546854
rect 162448 546586 162768 546618
rect 193168 547174 193488 547206
rect 193168 546938 193210 547174
rect 193446 546938 193488 547174
rect 193168 546854 193488 546938
rect 193168 546618 193210 546854
rect 193446 546618 193488 546854
rect 193168 546586 193488 546618
rect 223888 547174 224208 547206
rect 223888 546938 223930 547174
rect 224166 546938 224208 547174
rect 223888 546854 224208 546938
rect 223888 546618 223930 546854
rect 224166 546618 224208 546854
rect 223888 546586 224208 546618
rect 254608 547174 254928 547206
rect 254608 546938 254650 547174
rect 254886 546938 254928 547174
rect 254608 546854 254928 546938
rect 254608 546618 254650 546854
rect 254886 546618 254928 546854
rect 254608 546586 254928 546618
rect 285328 547174 285648 547206
rect 285328 546938 285370 547174
rect 285606 546938 285648 547174
rect 285328 546854 285648 546938
rect 285328 546618 285370 546854
rect 285606 546618 285648 546854
rect 285328 546586 285648 546618
rect 316048 547174 316368 547206
rect 316048 546938 316090 547174
rect 316326 546938 316368 547174
rect 316048 546854 316368 546938
rect 316048 546618 316090 546854
rect 316326 546618 316368 546854
rect 316048 546586 316368 546618
rect 54928 543454 55248 543486
rect 54928 543218 54970 543454
rect 55206 543218 55248 543454
rect 54928 543134 55248 543218
rect 54928 542898 54970 543134
rect 55206 542898 55248 543134
rect 54928 542866 55248 542898
rect 85648 543454 85968 543486
rect 85648 543218 85690 543454
rect 85926 543218 85968 543454
rect 85648 543134 85968 543218
rect 85648 542898 85690 543134
rect 85926 542898 85968 543134
rect 85648 542866 85968 542898
rect 116368 543454 116688 543486
rect 116368 543218 116410 543454
rect 116646 543218 116688 543454
rect 116368 543134 116688 543218
rect 116368 542898 116410 543134
rect 116646 542898 116688 543134
rect 116368 542866 116688 542898
rect 147088 543454 147408 543486
rect 147088 543218 147130 543454
rect 147366 543218 147408 543454
rect 147088 543134 147408 543218
rect 147088 542898 147130 543134
rect 147366 542898 147408 543134
rect 147088 542866 147408 542898
rect 177808 543454 178128 543486
rect 177808 543218 177850 543454
rect 178086 543218 178128 543454
rect 177808 543134 178128 543218
rect 177808 542898 177850 543134
rect 178086 542898 178128 543134
rect 177808 542866 178128 542898
rect 208528 543454 208848 543486
rect 208528 543218 208570 543454
rect 208806 543218 208848 543454
rect 208528 543134 208848 543218
rect 208528 542898 208570 543134
rect 208806 542898 208848 543134
rect 208528 542866 208848 542898
rect 239248 543454 239568 543486
rect 239248 543218 239290 543454
rect 239526 543218 239568 543454
rect 239248 543134 239568 543218
rect 239248 542898 239290 543134
rect 239526 542898 239568 543134
rect 239248 542866 239568 542898
rect 269968 543454 270288 543486
rect 269968 543218 270010 543454
rect 270246 543218 270288 543454
rect 269968 543134 270288 543218
rect 269968 542898 270010 543134
rect 270246 542898 270288 543134
rect 269968 542866 270288 542898
rect 300688 543454 301008 543486
rect 300688 543218 300730 543454
rect 300966 543218 301008 543454
rect 300688 543134 301008 543218
rect 300688 542898 300730 543134
rect 300966 542898 301008 543134
rect 300688 542866 301008 542898
rect 331408 543454 331728 543486
rect 331408 543218 331450 543454
rect 331686 543218 331728 543454
rect 331408 543134 331728 543218
rect 331408 542898 331450 543134
rect 331686 542898 331728 543134
rect 331408 542866 331728 542898
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 344394 526054 345014 561498
rect 348114 565774 348734 601218
rect 348114 565538 348146 565774
rect 348382 565538 348466 565774
rect 348702 565538 348734 565774
rect 348114 565454 348734 565538
rect 348114 565218 348146 565454
rect 348382 565218 348466 565454
rect 348702 565218 348734 565454
rect 346768 547174 347088 547206
rect 346768 546938 346810 547174
rect 347046 546938 347088 547174
rect 346768 546854 347088 546938
rect 346768 546618 346810 546854
rect 347046 546618 347088 546854
rect 346768 546586 347088 546618
rect 344394 525818 344426 526054
rect 344662 525818 344746 526054
rect 344982 525818 345014 526054
rect 344394 525734 345014 525818
rect 344394 525498 344426 525734
rect 344662 525498 344746 525734
rect 344982 525498 345014 525734
rect 70288 511174 70608 511206
rect 70288 510938 70330 511174
rect 70566 510938 70608 511174
rect 70288 510854 70608 510938
rect 70288 510618 70330 510854
rect 70566 510618 70608 510854
rect 70288 510586 70608 510618
rect 101008 511174 101328 511206
rect 101008 510938 101050 511174
rect 101286 510938 101328 511174
rect 101008 510854 101328 510938
rect 101008 510618 101050 510854
rect 101286 510618 101328 510854
rect 101008 510586 101328 510618
rect 131728 511174 132048 511206
rect 131728 510938 131770 511174
rect 132006 510938 132048 511174
rect 131728 510854 132048 510938
rect 131728 510618 131770 510854
rect 132006 510618 132048 510854
rect 131728 510586 132048 510618
rect 162448 511174 162768 511206
rect 162448 510938 162490 511174
rect 162726 510938 162768 511174
rect 162448 510854 162768 510938
rect 162448 510618 162490 510854
rect 162726 510618 162768 510854
rect 162448 510586 162768 510618
rect 193168 511174 193488 511206
rect 193168 510938 193210 511174
rect 193446 510938 193488 511174
rect 193168 510854 193488 510938
rect 193168 510618 193210 510854
rect 193446 510618 193488 510854
rect 193168 510586 193488 510618
rect 223888 511174 224208 511206
rect 223888 510938 223930 511174
rect 224166 510938 224208 511174
rect 223888 510854 224208 510938
rect 223888 510618 223930 510854
rect 224166 510618 224208 510854
rect 223888 510586 224208 510618
rect 254608 511174 254928 511206
rect 254608 510938 254650 511174
rect 254886 510938 254928 511174
rect 254608 510854 254928 510938
rect 254608 510618 254650 510854
rect 254886 510618 254928 510854
rect 254608 510586 254928 510618
rect 285328 511174 285648 511206
rect 285328 510938 285370 511174
rect 285606 510938 285648 511174
rect 285328 510854 285648 510938
rect 285328 510618 285370 510854
rect 285606 510618 285648 510854
rect 285328 510586 285648 510618
rect 316048 511174 316368 511206
rect 316048 510938 316090 511174
rect 316326 510938 316368 511174
rect 316048 510854 316368 510938
rect 316048 510618 316090 510854
rect 316326 510618 316368 510854
rect 316048 510586 316368 510618
rect 54928 507454 55248 507486
rect 54928 507218 54970 507454
rect 55206 507218 55248 507454
rect 54928 507134 55248 507218
rect 54928 506898 54970 507134
rect 55206 506898 55248 507134
rect 54928 506866 55248 506898
rect 85648 507454 85968 507486
rect 85648 507218 85690 507454
rect 85926 507218 85968 507454
rect 85648 507134 85968 507218
rect 85648 506898 85690 507134
rect 85926 506898 85968 507134
rect 85648 506866 85968 506898
rect 116368 507454 116688 507486
rect 116368 507218 116410 507454
rect 116646 507218 116688 507454
rect 116368 507134 116688 507218
rect 116368 506898 116410 507134
rect 116646 506898 116688 507134
rect 116368 506866 116688 506898
rect 147088 507454 147408 507486
rect 147088 507218 147130 507454
rect 147366 507218 147408 507454
rect 147088 507134 147408 507218
rect 147088 506898 147130 507134
rect 147366 506898 147408 507134
rect 147088 506866 147408 506898
rect 177808 507454 178128 507486
rect 177808 507218 177850 507454
rect 178086 507218 178128 507454
rect 177808 507134 178128 507218
rect 177808 506898 177850 507134
rect 178086 506898 178128 507134
rect 177808 506866 178128 506898
rect 208528 507454 208848 507486
rect 208528 507218 208570 507454
rect 208806 507218 208848 507454
rect 208528 507134 208848 507218
rect 208528 506898 208570 507134
rect 208806 506898 208848 507134
rect 208528 506866 208848 506898
rect 239248 507454 239568 507486
rect 239248 507218 239290 507454
rect 239526 507218 239568 507454
rect 239248 507134 239568 507218
rect 239248 506898 239290 507134
rect 239526 506898 239568 507134
rect 239248 506866 239568 506898
rect 269968 507454 270288 507486
rect 269968 507218 270010 507454
rect 270246 507218 270288 507454
rect 269968 507134 270288 507218
rect 269968 506898 270010 507134
rect 270246 506898 270288 507134
rect 269968 506866 270288 506898
rect 300688 507454 301008 507486
rect 300688 507218 300730 507454
rect 300966 507218 301008 507454
rect 300688 507134 301008 507218
rect 300688 506898 300730 507134
rect 300966 506898 301008 507134
rect 300688 506866 301008 506898
rect 331408 507454 331728 507486
rect 331408 507218 331450 507454
rect 331686 507218 331728 507454
rect 331408 507134 331728 507218
rect 331408 506898 331450 507134
rect 331686 506898 331728 507134
rect 331408 506866 331728 506898
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 344394 490054 345014 525498
rect 348114 529774 348734 565218
rect 348114 529538 348146 529774
rect 348382 529538 348466 529774
rect 348702 529538 348734 529774
rect 348114 529454 348734 529538
rect 348114 529218 348146 529454
rect 348382 529218 348466 529454
rect 348702 529218 348734 529454
rect 346768 511174 347088 511206
rect 346768 510938 346810 511174
rect 347046 510938 347088 511174
rect 346768 510854 347088 510938
rect 346768 510618 346810 510854
rect 347046 510618 347088 510854
rect 346768 510586 347088 510618
rect 344394 489818 344426 490054
rect 344662 489818 344746 490054
rect 344982 489818 345014 490054
rect 344394 489734 345014 489818
rect 344394 489498 344426 489734
rect 344662 489498 344746 489734
rect 344982 489498 345014 489734
rect 70288 475174 70608 475206
rect 70288 474938 70330 475174
rect 70566 474938 70608 475174
rect 70288 474854 70608 474938
rect 70288 474618 70330 474854
rect 70566 474618 70608 474854
rect 70288 474586 70608 474618
rect 101008 475174 101328 475206
rect 101008 474938 101050 475174
rect 101286 474938 101328 475174
rect 101008 474854 101328 474938
rect 101008 474618 101050 474854
rect 101286 474618 101328 474854
rect 101008 474586 101328 474618
rect 131728 475174 132048 475206
rect 131728 474938 131770 475174
rect 132006 474938 132048 475174
rect 131728 474854 132048 474938
rect 131728 474618 131770 474854
rect 132006 474618 132048 474854
rect 131728 474586 132048 474618
rect 162448 475174 162768 475206
rect 162448 474938 162490 475174
rect 162726 474938 162768 475174
rect 162448 474854 162768 474938
rect 162448 474618 162490 474854
rect 162726 474618 162768 474854
rect 162448 474586 162768 474618
rect 193168 475174 193488 475206
rect 193168 474938 193210 475174
rect 193446 474938 193488 475174
rect 193168 474854 193488 474938
rect 193168 474618 193210 474854
rect 193446 474618 193488 474854
rect 193168 474586 193488 474618
rect 223888 475174 224208 475206
rect 223888 474938 223930 475174
rect 224166 474938 224208 475174
rect 223888 474854 224208 474938
rect 223888 474618 223930 474854
rect 224166 474618 224208 474854
rect 223888 474586 224208 474618
rect 254608 475174 254928 475206
rect 254608 474938 254650 475174
rect 254886 474938 254928 475174
rect 254608 474854 254928 474938
rect 254608 474618 254650 474854
rect 254886 474618 254928 474854
rect 254608 474586 254928 474618
rect 285328 475174 285648 475206
rect 285328 474938 285370 475174
rect 285606 474938 285648 475174
rect 285328 474854 285648 474938
rect 285328 474618 285370 474854
rect 285606 474618 285648 474854
rect 285328 474586 285648 474618
rect 316048 475174 316368 475206
rect 316048 474938 316090 475174
rect 316326 474938 316368 475174
rect 316048 474854 316368 474938
rect 316048 474618 316090 474854
rect 316326 474618 316368 474854
rect 316048 474586 316368 474618
rect 54928 471454 55248 471486
rect 54928 471218 54970 471454
rect 55206 471218 55248 471454
rect 54928 471134 55248 471218
rect 54928 470898 54970 471134
rect 55206 470898 55248 471134
rect 54928 470866 55248 470898
rect 85648 471454 85968 471486
rect 85648 471218 85690 471454
rect 85926 471218 85968 471454
rect 85648 471134 85968 471218
rect 85648 470898 85690 471134
rect 85926 470898 85968 471134
rect 85648 470866 85968 470898
rect 116368 471454 116688 471486
rect 116368 471218 116410 471454
rect 116646 471218 116688 471454
rect 116368 471134 116688 471218
rect 116368 470898 116410 471134
rect 116646 470898 116688 471134
rect 116368 470866 116688 470898
rect 147088 471454 147408 471486
rect 147088 471218 147130 471454
rect 147366 471218 147408 471454
rect 147088 471134 147408 471218
rect 147088 470898 147130 471134
rect 147366 470898 147408 471134
rect 147088 470866 147408 470898
rect 177808 471454 178128 471486
rect 177808 471218 177850 471454
rect 178086 471218 178128 471454
rect 177808 471134 178128 471218
rect 177808 470898 177850 471134
rect 178086 470898 178128 471134
rect 177808 470866 178128 470898
rect 208528 471454 208848 471486
rect 208528 471218 208570 471454
rect 208806 471218 208848 471454
rect 208528 471134 208848 471218
rect 208528 470898 208570 471134
rect 208806 470898 208848 471134
rect 208528 470866 208848 470898
rect 239248 471454 239568 471486
rect 239248 471218 239290 471454
rect 239526 471218 239568 471454
rect 239248 471134 239568 471218
rect 239248 470898 239290 471134
rect 239526 470898 239568 471134
rect 239248 470866 239568 470898
rect 269968 471454 270288 471486
rect 269968 471218 270010 471454
rect 270246 471218 270288 471454
rect 269968 471134 270288 471218
rect 269968 470898 270010 471134
rect 270246 470898 270288 471134
rect 269968 470866 270288 470898
rect 300688 471454 301008 471486
rect 300688 471218 300730 471454
rect 300966 471218 301008 471454
rect 300688 471134 301008 471218
rect 300688 470898 300730 471134
rect 300966 470898 301008 471134
rect 300688 470866 301008 470898
rect 331408 471454 331728 471486
rect 331408 471218 331450 471454
rect 331686 471218 331728 471454
rect 331408 471134 331728 471218
rect 331408 470898 331450 471134
rect 331686 470898 331728 471134
rect 331408 470866 331728 470898
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 344394 454054 345014 489498
rect 348114 493774 348734 529218
rect 348114 493538 348146 493774
rect 348382 493538 348466 493774
rect 348702 493538 348734 493774
rect 348114 493454 348734 493538
rect 348114 493218 348146 493454
rect 348382 493218 348466 493454
rect 348702 493218 348734 493454
rect 346768 475174 347088 475206
rect 346768 474938 346810 475174
rect 347046 474938 347088 475174
rect 346768 474854 347088 474938
rect 346768 474618 346810 474854
rect 347046 474618 347088 474854
rect 346768 474586 347088 474618
rect 344394 453818 344426 454054
rect 344662 453818 344746 454054
rect 344982 453818 345014 454054
rect 344394 453734 345014 453818
rect 344394 453498 344426 453734
rect 344662 453498 344746 453734
rect 344982 453498 345014 453734
rect 70288 439174 70608 439206
rect 70288 438938 70330 439174
rect 70566 438938 70608 439174
rect 70288 438854 70608 438938
rect 70288 438618 70330 438854
rect 70566 438618 70608 438854
rect 70288 438586 70608 438618
rect 101008 439174 101328 439206
rect 101008 438938 101050 439174
rect 101286 438938 101328 439174
rect 101008 438854 101328 438938
rect 101008 438618 101050 438854
rect 101286 438618 101328 438854
rect 101008 438586 101328 438618
rect 131728 439174 132048 439206
rect 131728 438938 131770 439174
rect 132006 438938 132048 439174
rect 131728 438854 132048 438938
rect 131728 438618 131770 438854
rect 132006 438618 132048 438854
rect 131728 438586 132048 438618
rect 162448 439174 162768 439206
rect 162448 438938 162490 439174
rect 162726 438938 162768 439174
rect 162448 438854 162768 438938
rect 162448 438618 162490 438854
rect 162726 438618 162768 438854
rect 162448 438586 162768 438618
rect 193168 439174 193488 439206
rect 193168 438938 193210 439174
rect 193446 438938 193488 439174
rect 193168 438854 193488 438938
rect 193168 438618 193210 438854
rect 193446 438618 193488 438854
rect 193168 438586 193488 438618
rect 223888 439174 224208 439206
rect 223888 438938 223930 439174
rect 224166 438938 224208 439174
rect 223888 438854 224208 438938
rect 223888 438618 223930 438854
rect 224166 438618 224208 438854
rect 223888 438586 224208 438618
rect 254608 439174 254928 439206
rect 254608 438938 254650 439174
rect 254886 438938 254928 439174
rect 254608 438854 254928 438938
rect 254608 438618 254650 438854
rect 254886 438618 254928 438854
rect 254608 438586 254928 438618
rect 285328 439174 285648 439206
rect 285328 438938 285370 439174
rect 285606 438938 285648 439174
rect 285328 438854 285648 438938
rect 285328 438618 285370 438854
rect 285606 438618 285648 438854
rect 285328 438586 285648 438618
rect 316048 439174 316368 439206
rect 316048 438938 316090 439174
rect 316326 438938 316368 439174
rect 316048 438854 316368 438938
rect 316048 438618 316090 438854
rect 316326 438618 316368 438854
rect 316048 438586 316368 438618
rect 54928 435454 55248 435486
rect 54928 435218 54970 435454
rect 55206 435218 55248 435454
rect 54928 435134 55248 435218
rect 54928 434898 54970 435134
rect 55206 434898 55248 435134
rect 54928 434866 55248 434898
rect 85648 435454 85968 435486
rect 85648 435218 85690 435454
rect 85926 435218 85968 435454
rect 85648 435134 85968 435218
rect 85648 434898 85690 435134
rect 85926 434898 85968 435134
rect 85648 434866 85968 434898
rect 116368 435454 116688 435486
rect 116368 435218 116410 435454
rect 116646 435218 116688 435454
rect 116368 435134 116688 435218
rect 116368 434898 116410 435134
rect 116646 434898 116688 435134
rect 116368 434866 116688 434898
rect 147088 435454 147408 435486
rect 147088 435218 147130 435454
rect 147366 435218 147408 435454
rect 147088 435134 147408 435218
rect 147088 434898 147130 435134
rect 147366 434898 147408 435134
rect 147088 434866 147408 434898
rect 177808 435454 178128 435486
rect 177808 435218 177850 435454
rect 178086 435218 178128 435454
rect 177808 435134 178128 435218
rect 177808 434898 177850 435134
rect 178086 434898 178128 435134
rect 177808 434866 178128 434898
rect 208528 435454 208848 435486
rect 208528 435218 208570 435454
rect 208806 435218 208848 435454
rect 208528 435134 208848 435218
rect 208528 434898 208570 435134
rect 208806 434898 208848 435134
rect 208528 434866 208848 434898
rect 239248 435454 239568 435486
rect 239248 435218 239290 435454
rect 239526 435218 239568 435454
rect 239248 435134 239568 435218
rect 239248 434898 239290 435134
rect 239526 434898 239568 435134
rect 239248 434866 239568 434898
rect 269968 435454 270288 435486
rect 269968 435218 270010 435454
rect 270246 435218 270288 435454
rect 269968 435134 270288 435218
rect 269968 434898 270010 435134
rect 270246 434898 270288 435134
rect 269968 434866 270288 434898
rect 300688 435454 301008 435486
rect 300688 435218 300730 435454
rect 300966 435218 301008 435454
rect 300688 435134 301008 435218
rect 300688 434898 300730 435134
rect 300966 434898 301008 435134
rect 300688 434866 301008 434898
rect 331408 435454 331728 435486
rect 331408 435218 331450 435454
rect 331686 435218 331728 435454
rect 331408 435134 331728 435218
rect 331408 434898 331450 435134
rect 331686 434898 331728 435134
rect 331408 434866 331728 434898
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 344394 418054 345014 453498
rect 348114 457774 348734 493218
rect 348114 457538 348146 457774
rect 348382 457538 348466 457774
rect 348702 457538 348734 457774
rect 348114 457454 348734 457538
rect 348114 457218 348146 457454
rect 348382 457218 348466 457454
rect 348702 457218 348734 457454
rect 346768 439174 347088 439206
rect 346768 438938 346810 439174
rect 347046 438938 347088 439174
rect 346768 438854 347088 438938
rect 346768 438618 346810 438854
rect 347046 438618 347088 438854
rect 346768 438586 347088 438618
rect 344394 417818 344426 418054
rect 344662 417818 344746 418054
rect 344982 417818 345014 418054
rect 344394 417734 345014 417818
rect 344394 417498 344426 417734
rect 344662 417498 344746 417734
rect 344982 417498 345014 417734
rect 70288 403174 70608 403206
rect 70288 402938 70330 403174
rect 70566 402938 70608 403174
rect 70288 402854 70608 402938
rect 70288 402618 70330 402854
rect 70566 402618 70608 402854
rect 70288 402586 70608 402618
rect 101008 403174 101328 403206
rect 101008 402938 101050 403174
rect 101286 402938 101328 403174
rect 101008 402854 101328 402938
rect 101008 402618 101050 402854
rect 101286 402618 101328 402854
rect 101008 402586 101328 402618
rect 131728 403174 132048 403206
rect 131728 402938 131770 403174
rect 132006 402938 132048 403174
rect 131728 402854 132048 402938
rect 131728 402618 131770 402854
rect 132006 402618 132048 402854
rect 131728 402586 132048 402618
rect 162448 403174 162768 403206
rect 162448 402938 162490 403174
rect 162726 402938 162768 403174
rect 162448 402854 162768 402938
rect 162448 402618 162490 402854
rect 162726 402618 162768 402854
rect 162448 402586 162768 402618
rect 193168 403174 193488 403206
rect 193168 402938 193210 403174
rect 193446 402938 193488 403174
rect 193168 402854 193488 402938
rect 193168 402618 193210 402854
rect 193446 402618 193488 402854
rect 193168 402586 193488 402618
rect 223888 403174 224208 403206
rect 223888 402938 223930 403174
rect 224166 402938 224208 403174
rect 223888 402854 224208 402938
rect 223888 402618 223930 402854
rect 224166 402618 224208 402854
rect 223888 402586 224208 402618
rect 254608 403174 254928 403206
rect 254608 402938 254650 403174
rect 254886 402938 254928 403174
rect 254608 402854 254928 402938
rect 254608 402618 254650 402854
rect 254886 402618 254928 402854
rect 254608 402586 254928 402618
rect 285328 403174 285648 403206
rect 285328 402938 285370 403174
rect 285606 402938 285648 403174
rect 285328 402854 285648 402938
rect 285328 402618 285370 402854
rect 285606 402618 285648 402854
rect 285328 402586 285648 402618
rect 316048 403174 316368 403206
rect 316048 402938 316090 403174
rect 316326 402938 316368 403174
rect 316048 402854 316368 402938
rect 316048 402618 316090 402854
rect 316326 402618 316368 402854
rect 316048 402586 316368 402618
rect 54928 399454 55248 399486
rect 54928 399218 54970 399454
rect 55206 399218 55248 399454
rect 54928 399134 55248 399218
rect 54928 398898 54970 399134
rect 55206 398898 55248 399134
rect 54928 398866 55248 398898
rect 85648 399454 85968 399486
rect 85648 399218 85690 399454
rect 85926 399218 85968 399454
rect 85648 399134 85968 399218
rect 85648 398898 85690 399134
rect 85926 398898 85968 399134
rect 85648 398866 85968 398898
rect 116368 399454 116688 399486
rect 116368 399218 116410 399454
rect 116646 399218 116688 399454
rect 116368 399134 116688 399218
rect 116368 398898 116410 399134
rect 116646 398898 116688 399134
rect 116368 398866 116688 398898
rect 147088 399454 147408 399486
rect 147088 399218 147130 399454
rect 147366 399218 147408 399454
rect 147088 399134 147408 399218
rect 147088 398898 147130 399134
rect 147366 398898 147408 399134
rect 147088 398866 147408 398898
rect 177808 399454 178128 399486
rect 177808 399218 177850 399454
rect 178086 399218 178128 399454
rect 177808 399134 178128 399218
rect 177808 398898 177850 399134
rect 178086 398898 178128 399134
rect 177808 398866 178128 398898
rect 208528 399454 208848 399486
rect 208528 399218 208570 399454
rect 208806 399218 208848 399454
rect 208528 399134 208848 399218
rect 208528 398898 208570 399134
rect 208806 398898 208848 399134
rect 208528 398866 208848 398898
rect 239248 399454 239568 399486
rect 239248 399218 239290 399454
rect 239526 399218 239568 399454
rect 239248 399134 239568 399218
rect 239248 398898 239290 399134
rect 239526 398898 239568 399134
rect 239248 398866 239568 398898
rect 269968 399454 270288 399486
rect 269968 399218 270010 399454
rect 270246 399218 270288 399454
rect 269968 399134 270288 399218
rect 269968 398898 270010 399134
rect 270246 398898 270288 399134
rect 269968 398866 270288 398898
rect 300688 399454 301008 399486
rect 300688 399218 300730 399454
rect 300966 399218 301008 399454
rect 300688 399134 301008 399218
rect 300688 398898 300730 399134
rect 300966 398898 301008 399134
rect 300688 398866 301008 398898
rect 331408 399454 331728 399486
rect 331408 399218 331450 399454
rect 331686 399218 331728 399454
rect 331408 399134 331728 399218
rect 331408 398898 331450 399134
rect 331686 398898 331728 399134
rect 331408 398866 331728 398898
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 344394 382054 345014 417498
rect 348114 421774 348734 457218
rect 348114 421538 348146 421774
rect 348382 421538 348466 421774
rect 348702 421538 348734 421774
rect 348114 421454 348734 421538
rect 348114 421218 348146 421454
rect 348382 421218 348466 421454
rect 348702 421218 348734 421454
rect 346768 403174 347088 403206
rect 346768 402938 346810 403174
rect 347046 402938 347088 403174
rect 346768 402854 347088 402938
rect 346768 402618 346810 402854
rect 347046 402618 347088 402854
rect 346768 402586 347088 402618
rect 344394 381818 344426 382054
rect 344662 381818 344746 382054
rect 344982 381818 345014 382054
rect 344394 381734 345014 381818
rect 344394 381498 344426 381734
rect 344662 381498 344746 381734
rect 344982 381498 345014 381734
rect 70288 367174 70608 367206
rect 70288 366938 70330 367174
rect 70566 366938 70608 367174
rect 70288 366854 70608 366938
rect 70288 366618 70330 366854
rect 70566 366618 70608 366854
rect 70288 366586 70608 366618
rect 101008 367174 101328 367206
rect 101008 366938 101050 367174
rect 101286 366938 101328 367174
rect 101008 366854 101328 366938
rect 101008 366618 101050 366854
rect 101286 366618 101328 366854
rect 101008 366586 101328 366618
rect 131728 367174 132048 367206
rect 131728 366938 131770 367174
rect 132006 366938 132048 367174
rect 131728 366854 132048 366938
rect 131728 366618 131770 366854
rect 132006 366618 132048 366854
rect 131728 366586 132048 366618
rect 162448 367174 162768 367206
rect 162448 366938 162490 367174
rect 162726 366938 162768 367174
rect 162448 366854 162768 366938
rect 162448 366618 162490 366854
rect 162726 366618 162768 366854
rect 162448 366586 162768 366618
rect 193168 367174 193488 367206
rect 193168 366938 193210 367174
rect 193446 366938 193488 367174
rect 193168 366854 193488 366938
rect 193168 366618 193210 366854
rect 193446 366618 193488 366854
rect 193168 366586 193488 366618
rect 223888 367174 224208 367206
rect 223888 366938 223930 367174
rect 224166 366938 224208 367174
rect 223888 366854 224208 366938
rect 223888 366618 223930 366854
rect 224166 366618 224208 366854
rect 223888 366586 224208 366618
rect 254608 367174 254928 367206
rect 254608 366938 254650 367174
rect 254886 366938 254928 367174
rect 254608 366854 254928 366938
rect 254608 366618 254650 366854
rect 254886 366618 254928 366854
rect 254608 366586 254928 366618
rect 285328 367174 285648 367206
rect 285328 366938 285370 367174
rect 285606 366938 285648 367174
rect 285328 366854 285648 366938
rect 285328 366618 285370 366854
rect 285606 366618 285648 366854
rect 285328 366586 285648 366618
rect 316048 367174 316368 367206
rect 316048 366938 316090 367174
rect 316326 366938 316368 367174
rect 316048 366854 316368 366938
rect 316048 366618 316090 366854
rect 316326 366618 316368 366854
rect 316048 366586 316368 366618
rect 54928 363454 55248 363486
rect 54928 363218 54970 363454
rect 55206 363218 55248 363454
rect 54928 363134 55248 363218
rect 54928 362898 54970 363134
rect 55206 362898 55248 363134
rect 54928 362866 55248 362898
rect 85648 363454 85968 363486
rect 85648 363218 85690 363454
rect 85926 363218 85968 363454
rect 85648 363134 85968 363218
rect 85648 362898 85690 363134
rect 85926 362898 85968 363134
rect 85648 362866 85968 362898
rect 116368 363454 116688 363486
rect 116368 363218 116410 363454
rect 116646 363218 116688 363454
rect 116368 363134 116688 363218
rect 116368 362898 116410 363134
rect 116646 362898 116688 363134
rect 116368 362866 116688 362898
rect 147088 363454 147408 363486
rect 147088 363218 147130 363454
rect 147366 363218 147408 363454
rect 147088 363134 147408 363218
rect 147088 362898 147130 363134
rect 147366 362898 147408 363134
rect 147088 362866 147408 362898
rect 177808 363454 178128 363486
rect 177808 363218 177850 363454
rect 178086 363218 178128 363454
rect 177808 363134 178128 363218
rect 177808 362898 177850 363134
rect 178086 362898 178128 363134
rect 177808 362866 178128 362898
rect 208528 363454 208848 363486
rect 208528 363218 208570 363454
rect 208806 363218 208848 363454
rect 208528 363134 208848 363218
rect 208528 362898 208570 363134
rect 208806 362898 208848 363134
rect 208528 362866 208848 362898
rect 239248 363454 239568 363486
rect 239248 363218 239290 363454
rect 239526 363218 239568 363454
rect 239248 363134 239568 363218
rect 239248 362898 239290 363134
rect 239526 362898 239568 363134
rect 239248 362866 239568 362898
rect 269968 363454 270288 363486
rect 269968 363218 270010 363454
rect 270246 363218 270288 363454
rect 269968 363134 270288 363218
rect 269968 362898 270010 363134
rect 270246 362898 270288 363134
rect 269968 362866 270288 362898
rect 300688 363454 301008 363486
rect 300688 363218 300730 363454
rect 300966 363218 301008 363454
rect 300688 363134 301008 363218
rect 300688 362898 300730 363134
rect 300966 362898 301008 363134
rect 300688 362866 301008 362898
rect 331408 363454 331728 363486
rect 331408 363218 331450 363454
rect 331686 363218 331728 363454
rect 331408 363134 331728 363218
rect 331408 362898 331450 363134
rect 331686 362898 331728 363134
rect 331408 362866 331728 362898
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 344394 346054 345014 381498
rect 348114 385774 348734 421218
rect 348114 385538 348146 385774
rect 348382 385538 348466 385774
rect 348702 385538 348734 385774
rect 348114 385454 348734 385538
rect 348114 385218 348146 385454
rect 348382 385218 348466 385454
rect 348702 385218 348734 385454
rect 346768 367174 347088 367206
rect 346768 366938 346810 367174
rect 347046 366938 347088 367174
rect 346768 366854 347088 366938
rect 346768 366618 346810 366854
rect 347046 366618 347088 366854
rect 346768 366586 347088 366618
rect 344394 345818 344426 346054
rect 344662 345818 344746 346054
rect 344982 345818 345014 346054
rect 344394 345734 345014 345818
rect 344394 345498 344426 345734
rect 344662 345498 344746 345734
rect 344982 345498 345014 345734
rect 70288 331174 70608 331206
rect 70288 330938 70330 331174
rect 70566 330938 70608 331174
rect 70288 330854 70608 330938
rect 70288 330618 70330 330854
rect 70566 330618 70608 330854
rect 70288 330586 70608 330618
rect 101008 331174 101328 331206
rect 101008 330938 101050 331174
rect 101286 330938 101328 331174
rect 101008 330854 101328 330938
rect 101008 330618 101050 330854
rect 101286 330618 101328 330854
rect 101008 330586 101328 330618
rect 131728 331174 132048 331206
rect 131728 330938 131770 331174
rect 132006 330938 132048 331174
rect 131728 330854 132048 330938
rect 131728 330618 131770 330854
rect 132006 330618 132048 330854
rect 131728 330586 132048 330618
rect 162448 331174 162768 331206
rect 162448 330938 162490 331174
rect 162726 330938 162768 331174
rect 162448 330854 162768 330938
rect 162448 330618 162490 330854
rect 162726 330618 162768 330854
rect 162448 330586 162768 330618
rect 193168 331174 193488 331206
rect 193168 330938 193210 331174
rect 193446 330938 193488 331174
rect 193168 330854 193488 330938
rect 193168 330618 193210 330854
rect 193446 330618 193488 330854
rect 193168 330586 193488 330618
rect 223888 331174 224208 331206
rect 223888 330938 223930 331174
rect 224166 330938 224208 331174
rect 223888 330854 224208 330938
rect 223888 330618 223930 330854
rect 224166 330618 224208 330854
rect 223888 330586 224208 330618
rect 254608 331174 254928 331206
rect 254608 330938 254650 331174
rect 254886 330938 254928 331174
rect 254608 330854 254928 330938
rect 254608 330618 254650 330854
rect 254886 330618 254928 330854
rect 254608 330586 254928 330618
rect 285328 331174 285648 331206
rect 285328 330938 285370 331174
rect 285606 330938 285648 331174
rect 285328 330854 285648 330938
rect 285328 330618 285370 330854
rect 285606 330618 285648 330854
rect 285328 330586 285648 330618
rect 316048 331174 316368 331206
rect 316048 330938 316090 331174
rect 316326 330938 316368 331174
rect 316048 330854 316368 330938
rect 316048 330618 316090 330854
rect 316326 330618 316368 330854
rect 316048 330586 316368 330618
rect 54928 327454 55248 327486
rect 54928 327218 54970 327454
rect 55206 327218 55248 327454
rect 54928 327134 55248 327218
rect 54928 326898 54970 327134
rect 55206 326898 55248 327134
rect 54928 326866 55248 326898
rect 85648 327454 85968 327486
rect 85648 327218 85690 327454
rect 85926 327218 85968 327454
rect 85648 327134 85968 327218
rect 85648 326898 85690 327134
rect 85926 326898 85968 327134
rect 85648 326866 85968 326898
rect 116368 327454 116688 327486
rect 116368 327218 116410 327454
rect 116646 327218 116688 327454
rect 116368 327134 116688 327218
rect 116368 326898 116410 327134
rect 116646 326898 116688 327134
rect 116368 326866 116688 326898
rect 147088 327454 147408 327486
rect 147088 327218 147130 327454
rect 147366 327218 147408 327454
rect 147088 327134 147408 327218
rect 147088 326898 147130 327134
rect 147366 326898 147408 327134
rect 147088 326866 147408 326898
rect 177808 327454 178128 327486
rect 177808 327218 177850 327454
rect 178086 327218 178128 327454
rect 177808 327134 178128 327218
rect 177808 326898 177850 327134
rect 178086 326898 178128 327134
rect 177808 326866 178128 326898
rect 208528 327454 208848 327486
rect 208528 327218 208570 327454
rect 208806 327218 208848 327454
rect 208528 327134 208848 327218
rect 208528 326898 208570 327134
rect 208806 326898 208848 327134
rect 208528 326866 208848 326898
rect 239248 327454 239568 327486
rect 239248 327218 239290 327454
rect 239526 327218 239568 327454
rect 239248 327134 239568 327218
rect 239248 326898 239290 327134
rect 239526 326898 239568 327134
rect 239248 326866 239568 326898
rect 269968 327454 270288 327486
rect 269968 327218 270010 327454
rect 270246 327218 270288 327454
rect 269968 327134 270288 327218
rect 269968 326898 270010 327134
rect 270246 326898 270288 327134
rect 269968 326866 270288 326898
rect 300688 327454 301008 327486
rect 300688 327218 300730 327454
rect 300966 327218 301008 327454
rect 300688 327134 301008 327218
rect 300688 326898 300730 327134
rect 300966 326898 301008 327134
rect 300688 326866 301008 326898
rect 331408 327454 331728 327486
rect 331408 327218 331450 327454
rect 331686 327218 331728 327454
rect 331408 327134 331728 327218
rect 331408 326898 331450 327134
rect 331686 326898 331728 327134
rect 331408 326866 331728 326898
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 344394 310054 345014 345498
rect 348114 349774 348734 385218
rect 348114 349538 348146 349774
rect 348382 349538 348466 349774
rect 348702 349538 348734 349774
rect 348114 349454 348734 349538
rect 348114 349218 348146 349454
rect 348382 349218 348466 349454
rect 348702 349218 348734 349454
rect 346768 331174 347088 331206
rect 346768 330938 346810 331174
rect 347046 330938 347088 331174
rect 346768 330854 347088 330938
rect 346768 330618 346810 330854
rect 347046 330618 347088 330854
rect 346768 330586 347088 330618
rect 344394 309818 344426 310054
rect 344662 309818 344746 310054
rect 344982 309818 345014 310054
rect 344394 309734 345014 309818
rect 344394 309498 344426 309734
rect 344662 309498 344746 309734
rect 344982 309498 345014 309734
rect 70288 295174 70608 295206
rect 70288 294938 70330 295174
rect 70566 294938 70608 295174
rect 70288 294854 70608 294938
rect 70288 294618 70330 294854
rect 70566 294618 70608 294854
rect 70288 294586 70608 294618
rect 101008 295174 101328 295206
rect 101008 294938 101050 295174
rect 101286 294938 101328 295174
rect 101008 294854 101328 294938
rect 101008 294618 101050 294854
rect 101286 294618 101328 294854
rect 101008 294586 101328 294618
rect 131728 295174 132048 295206
rect 131728 294938 131770 295174
rect 132006 294938 132048 295174
rect 131728 294854 132048 294938
rect 131728 294618 131770 294854
rect 132006 294618 132048 294854
rect 131728 294586 132048 294618
rect 162448 295174 162768 295206
rect 162448 294938 162490 295174
rect 162726 294938 162768 295174
rect 162448 294854 162768 294938
rect 162448 294618 162490 294854
rect 162726 294618 162768 294854
rect 162448 294586 162768 294618
rect 193168 295174 193488 295206
rect 193168 294938 193210 295174
rect 193446 294938 193488 295174
rect 193168 294854 193488 294938
rect 193168 294618 193210 294854
rect 193446 294618 193488 294854
rect 193168 294586 193488 294618
rect 223888 295174 224208 295206
rect 223888 294938 223930 295174
rect 224166 294938 224208 295174
rect 223888 294854 224208 294938
rect 223888 294618 223930 294854
rect 224166 294618 224208 294854
rect 223888 294586 224208 294618
rect 254608 295174 254928 295206
rect 254608 294938 254650 295174
rect 254886 294938 254928 295174
rect 254608 294854 254928 294938
rect 254608 294618 254650 294854
rect 254886 294618 254928 294854
rect 254608 294586 254928 294618
rect 285328 295174 285648 295206
rect 285328 294938 285370 295174
rect 285606 294938 285648 295174
rect 285328 294854 285648 294938
rect 285328 294618 285370 294854
rect 285606 294618 285648 294854
rect 285328 294586 285648 294618
rect 316048 295174 316368 295206
rect 316048 294938 316090 295174
rect 316326 294938 316368 295174
rect 316048 294854 316368 294938
rect 316048 294618 316090 294854
rect 316326 294618 316368 294854
rect 316048 294586 316368 294618
rect 54928 291454 55248 291486
rect 54928 291218 54970 291454
rect 55206 291218 55248 291454
rect 54928 291134 55248 291218
rect 54928 290898 54970 291134
rect 55206 290898 55248 291134
rect 54928 290866 55248 290898
rect 85648 291454 85968 291486
rect 85648 291218 85690 291454
rect 85926 291218 85968 291454
rect 85648 291134 85968 291218
rect 85648 290898 85690 291134
rect 85926 290898 85968 291134
rect 85648 290866 85968 290898
rect 116368 291454 116688 291486
rect 116368 291218 116410 291454
rect 116646 291218 116688 291454
rect 116368 291134 116688 291218
rect 116368 290898 116410 291134
rect 116646 290898 116688 291134
rect 116368 290866 116688 290898
rect 147088 291454 147408 291486
rect 147088 291218 147130 291454
rect 147366 291218 147408 291454
rect 147088 291134 147408 291218
rect 147088 290898 147130 291134
rect 147366 290898 147408 291134
rect 147088 290866 147408 290898
rect 177808 291454 178128 291486
rect 177808 291218 177850 291454
rect 178086 291218 178128 291454
rect 177808 291134 178128 291218
rect 177808 290898 177850 291134
rect 178086 290898 178128 291134
rect 177808 290866 178128 290898
rect 208528 291454 208848 291486
rect 208528 291218 208570 291454
rect 208806 291218 208848 291454
rect 208528 291134 208848 291218
rect 208528 290898 208570 291134
rect 208806 290898 208848 291134
rect 208528 290866 208848 290898
rect 239248 291454 239568 291486
rect 239248 291218 239290 291454
rect 239526 291218 239568 291454
rect 239248 291134 239568 291218
rect 239248 290898 239290 291134
rect 239526 290898 239568 291134
rect 239248 290866 239568 290898
rect 269968 291454 270288 291486
rect 269968 291218 270010 291454
rect 270246 291218 270288 291454
rect 269968 291134 270288 291218
rect 269968 290898 270010 291134
rect 270246 290898 270288 291134
rect 269968 290866 270288 290898
rect 300688 291454 301008 291486
rect 300688 291218 300730 291454
rect 300966 291218 301008 291454
rect 300688 291134 301008 291218
rect 300688 290898 300730 291134
rect 300966 290898 301008 291134
rect 300688 290866 301008 290898
rect 331408 291454 331728 291486
rect 331408 291218 331450 291454
rect 331686 291218 331728 291454
rect 331408 291134 331728 291218
rect 331408 290898 331450 291134
rect 331686 290898 331728 291134
rect 331408 290866 331728 290898
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 344394 274054 345014 309498
rect 348114 313774 348734 349218
rect 348114 313538 348146 313774
rect 348382 313538 348466 313774
rect 348702 313538 348734 313774
rect 348114 313454 348734 313538
rect 348114 313218 348146 313454
rect 348382 313218 348466 313454
rect 348702 313218 348734 313454
rect 346768 295174 347088 295206
rect 346768 294938 346810 295174
rect 347046 294938 347088 295174
rect 346768 294854 347088 294938
rect 346768 294618 346810 294854
rect 347046 294618 347088 294854
rect 346768 294586 347088 294618
rect 344394 273818 344426 274054
rect 344662 273818 344746 274054
rect 344982 273818 345014 274054
rect 344394 273734 345014 273818
rect 344394 273498 344426 273734
rect 344662 273498 344746 273734
rect 344982 273498 345014 273734
rect 70288 259174 70608 259206
rect 70288 258938 70330 259174
rect 70566 258938 70608 259174
rect 70288 258854 70608 258938
rect 70288 258618 70330 258854
rect 70566 258618 70608 258854
rect 70288 258586 70608 258618
rect 101008 259174 101328 259206
rect 101008 258938 101050 259174
rect 101286 258938 101328 259174
rect 101008 258854 101328 258938
rect 101008 258618 101050 258854
rect 101286 258618 101328 258854
rect 101008 258586 101328 258618
rect 131728 259174 132048 259206
rect 131728 258938 131770 259174
rect 132006 258938 132048 259174
rect 131728 258854 132048 258938
rect 131728 258618 131770 258854
rect 132006 258618 132048 258854
rect 131728 258586 132048 258618
rect 162448 259174 162768 259206
rect 162448 258938 162490 259174
rect 162726 258938 162768 259174
rect 162448 258854 162768 258938
rect 162448 258618 162490 258854
rect 162726 258618 162768 258854
rect 162448 258586 162768 258618
rect 193168 259174 193488 259206
rect 193168 258938 193210 259174
rect 193446 258938 193488 259174
rect 193168 258854 193488 258938
rect 193168 258618 193210 258854
rect 193446 258618 193488 258854
rect 193168 258586 193488 258618
rect 223888 259174 224208 259206
rect 223888 258938 223930 259174
rect 224166 258938 224208 259174
rect 223888 258854 224208 258938
rect 223888 258618 223930 258854
rect 224166 258618 224208 258854
rect 223888 258586 224208 258618
rect 254608 259174 254928 259206
rect 254608 258938 254650 259174
rect 254886 258938 254928 259174
rect 254608 258854 254928 258938
rect 254608 258618 254650 258854
rect 254886 258618 254928 258854
rect 254608 258586 254928 258618
rect 285328 259174 285648 259206
rect 285328 258938 285370 259174
rect 285606 258938 285648 259174
rect 285328 258854 285648 258938
rect 285328 258618 285370 258854
rect 285606 258618 285648 258854
rect 285328 258586 285648 258618
rect 316048 259174 316368 259206
rect 316048 258938 316090 259174
rect 316326 258938 316368 259174
rect 316048 258854 316368 258938
rect 316048 258618 316090 258854
rect 316326 258618 316368 258854
rect 316048 258586 316368 258618
rect 54928 255454 55248 255486
rect 54928 255218 54970 255454
rect 55206 255218 55248 255454
rect 54928 255134 55248 255218
rect 54928 254898 54970 255134
rect 55206 254898 55248 255134
rect 54928 254866 55248 254898
rect 85648 255454 85968 255486
rect 85648 255218 85690 255454
rect 85926 255218 85968 255454
rect 85648 255134 85968 255218
rect 85648 254898 85690 255134
rect 85926 254898 85968 255134
rect 85648 254866 85968 254898
rect 116368 255454 116688 255486
rect 116368 255218 116410 255454
rect 116646 255218 116688 255454
rect 116368 255134 116688 255218
rect 116368 254898 116410 255134
rect 116646 254898 116688 255134
rect 116368 254866 116688 254898
rect 147088 255454 147408 255486
rect 147088 255218 147130 255454
rect 147366 255218 147408 255454
rect 147088 255134 147408 255218
rect 147088 254898 147130 255134
rect 147366 254898 147408 255134
rect 147088 254866 147408 254898
rect 177808 255454 178128 255486
rect 177808 255218 177850 255454
rect 178086 255218 178128 255454
rect 177808 255134 178128 255218
rect 177808 254898 177850 255134
rect 178086 254898 178128 255134
rect 177808 254866 178128 254898
rect 208528 255454 208848 255486
rect 208528 255218 208570 255454
rect 208806 255218 208848 255454
rect 208528 255134 208848 255218
rect 208528 254898 208570 255134
rect 208806 254898 208848 255134
rect 208528 254866 208848 254898
rect 239248 255454 239568 255486
rect 239248 255218 239290 255454
rect 239526 255218 239568 255454
rect 239248 255134 239568 255218
rect 239248 254898 239290 255134
rect 239526 254898 239568 255134
rect 239248 254866 239568 254898
rect 269968 255454 270288 255486
rect 269968 255218 270010 255454
rect 270246 255218 270288 255454
rect 269968 255134 270288 255218
rect 269968 254898 270010 255134
rect 270246 254898 270288 255134
rect 269968 254866 270288 254898
rect 300688 255454 301008 255486
rect 300688 255218 300730 255454
rect 300966 255218 301008 255454
rect 300688 255134 301008 255218
rect 300688 254898 300730 255134
rect 300966 254898 301008 255134
rect 300688 254866 301008 254898
rect 331408 255454 331728 255486
rect 331408 255218 331450 255454
rect 331686 255218 331728 255454
rect 331408 255134 331728 255218
rect 331408 254898 331450 255134
rect 331686 254898 331728 255134
rect 331408 254866 331728 254898
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 344394 238054 345014 273498
rect 348114 277774 348734 313218
rect 348114 277538 348146 277774
rect 348382 277538 348466 277774
rect 348702 277538 348734 277774
rect 348114 277454 348734 277538
rect 348114 277218 348146 277454
rect 348382 277218 348466 277454
rect 348702 277218 348734 277454
rect 346768 259174 347088 259206
rect 346768 258938 346810 259174
rect 347046 258938 347088 259174
rect 346768 258854 347088 258938
rect 346768 258618 346810 258854
rect 347046 258618 347088 258854
rect 346768 258586 347088 258618
rect 344394 237818 344426 238054
rect 344662 237818 344746 238054
rect 344982 237818 345014 238054
rect 344394 237734 345014 237818
rect 344394 237498 344426 237734
rect 344662 237498 344746 237734
rect 344982 237498 345014 237734
rect 70288 223174 70608 223206
rect 70288 222938 70330 223174
rect 70566 222938 70608 223174
rect 70288 222854 70608 222938
rect 70288 222618 70330 222854
rect 70566 222618 70608 222854
rect 70288 222586 70608 222618
rect 101008 223174 101328 223206
rect 101008 222938 101050 223174
rect 101286 222938 101328 223174
rect 101008 222854 101328 222938
rect 101008 222618 101050 222854
rect 101286 222618 101328 222854
rect 101008 222586 101328 222618
rect 131728 223174 132048 223206
rect 131728 222938 131770 223174
rect 132006 222938 132048 223174
rect 131728 222854 132048 222938
rect 131728 222618 131770 222854
rect 132006 222618 132048 222854
rect 131728 222586 132048 222618
rect 162448 223174 162768 223206
rect 162448 222938 162490 223174
rect 162726 222938 162768 223174
rect 162448 222854 162768 222938
rect 162448 222618 162490 222854
rect 162726 222618 162768 222854
rect 162448 222586 162768 222618
rect 193168 223174 193488 223206
rect 193168 222938 193210 223174
rect 193446 222938 193488 223174
rect 193168 222854 193488 222938
rect 193168 222618 193210 222854
rect 193446 222618 193488 222854
rect 193168 222586 193488 222618
rect 223888 223174 224208 223206
rect 223888 222938 223930 223174
rect 224166 222938 224208 223174
rect 223888 222854 224208 222938
rect 223888 222618 223930 222854
rect 224166 222618 224208 222854
rect 223888 222586 224208 222618
rect 254608 223174 254928 223206
rect 254608 222938 254650 223174
rect 254886 222938 254928 223174
rect 254608 222854 254928 222938
rect 254608 222618 254650 222854
rect 254886 222618 254928 222854
rect 254608 222586 254928 222618
rect 285328 223174 285648 223206
rect 285328 222938 285370 223174
rect 285606 222938 285648 223174
rect 285328 222854 285648 222938
rect 285328 222618 285370 222854
rect 285606 222618 285648 222854
rect 285328 222586 285648 222618
rect 316048 223174 316368 223206
rect 316048 222938 316090 223174
rect 316326 222938 316368 223174
rect 316048 222854 316368 222938
rect 316048 222618 316090 222854
rect 316326 222618 316368 222854
rect 316048 222586 316368 222618
rect 54928 219454 55248 219486
rect 54928 219218 54970 219454
rect 55206 219218 55248 219454
rect 54928 219134 55248 219218
rect 54928 218898 54970 219134
rect 55206 218898 55248 219134
rect 54928 218866 55248 218898
rect 85648 219454 85968 219486
rect 85648 219218 85690 219454
rect 85926 219218 85968 219454
rect 85648 219134 85968 219218
rect 85648 218898 85690 219134
rect 85926 218898 85968 219134
rect 85648 218866 85968 218898
rect 116368 219454 116688 219486
rect 116368 219218 116410 219454
rect 116646 219218 116688 219454
rect 116368 219134 116688 219218
rect 116368 218898 116410 219134
rect 116646 218898 116688 219134
rect 116368 218866 116688 218898
rect 147088 219454 147408 219486
rect 147088 219218 147130 219454
rect 147366 219218 147408 219454
rect 147088 219134 147408 219218
rect 147088 218898 147130 219134
rect 147366 218898 147408 219134
rect 147088 218866 147408 218898
rect 177808 219454 178128 219486
rect 177808 219218 177850 219454
rect 178086 219218 178128 219454
rect 177808 219134 178128 219218
rect 177808 218898 177850 219134
rect 178086 218898 178128 219134
rect 177808 218866 178128 218898
rect 208528 219454 208848 219486
rect 208528 219218 208570 219454
rect 208806 219218 208848 219454
rect 208528 219134 208848 219218
rect 208528 218898 208570 219134
rect 208806 218898 208848 219134
rect 208528 218866 208848 218898
rect 239248 219454 239568 219486
rect 239248 219218 239290 219454
rect 239526 219218 239568 219454
rect 239248 219134 239568 219218
rect 239248 218898 239290 219134
rect 239526 218898 239568 219134
rect 239248 218866 239568 218898
rect 269968 219454 270288 219486
rect 269968 219218 270010 219454
rect 270246 219218 270288 219454
rect 269968 219134 270288 219218
rect 269968 218898 270010 219134
rect 270246 218898 270288 219134
rect 269968 218866 270288 218898
rect 300688 219454 301008 219486
rect 300688 219218 300730 219454
rect 300966 219218 301008 219454
rect 300688 219134 301008 219218
rect 300688 218898 300730 219134
rect 300966 218898 301008 219134
rect 300688 218866 301008 218898
rect 331408 219454 331728 219486
rect 331408 219218 331450 219454
rect 331686 219218 331728 219454
rect 331408 219134 331728 219218
rect 331408 218898 331450 219134
rect 331686 218898 331728 219134
rect 331408 218866 331728 218898
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 344394 202054 345014 237498
rect 348114 241774 348734 277218
rect 348114 241538 348146 241774
rect 348382 241538 348466 241774
rect 348702 241538 348734 241774
rect 348114 241454 348734 241538
rect 348114 241218 348146 241454
rect 348382 241218 348466 241454
rect 348702 241218 348734 241454
rect 346768 223174 347088 223206
rect 346768 222938 346810 223174
rect 347046 222938 347088 223174
rect 346768 222854 347088 222938
rect 346768 222618 346810 222854
rect 347046 222618 347088 222854
rect 346768 222586 347088 222618
rect 344394 201818 344426 202054
rect 344662 201818 344746 202054
rect 344982 201818 345014 202054
rect 344394 201734 345014 201818
rect 344394 201498 344426 201734
rect 344662 201498 344746 201734
rect 344982 201498 345014 201734
rect 70288 187174 70608 187206
rect 70288 186938 70330 187174
rect 70566 186938 70608 187174
rect 70288 186854 70608 186938
rect 70288 186618 70330 186854
rect 70566 186618 70608 186854
rect 70288 186586 70608 186618
rect 101008 187174 101328 187206
rect 101008 186938 101050 187174
rect 101286 186938 101328 187174
rect 101008 186854 101328 186938
rect 101008 186618 101050 186854
rect 101286 186618 101328 186854
rect 101008 186586 101328 186618
rect 131728 187174 132048 187206
rect 131728 186938 131770 187174
rect 132006 186938 132048 187174
rect 131728 186854 132048 186938
rect 131728 186618 131770 186854
rect 132006 186618 132048 186854
rect 131728 186586 132048 186618
rect 162448 187174 162768 187206
rect 162448 186938 162490 187174
rect 162726 186938 162768 187174
rect 162448 186854 162768 186938
rect 162448 186618 162490 186854
rect 162726 186618 162768 186854
rect 162448 186586 162768 186618
rect 193168 187174 193488 187206
rect 193168 186938 193210 187174
rect 193446 186938 193488 187174
rect 193168 186854 193488 186938
rect 193168 186618 193210 186854
rect 193446 186618 193488 186854
rect 193168 186586 193488 186618
rect 223888 187174 224208 187206
rect 223888 186938 223930 187174
rect 224166 186938 224208 187174
rect 223888 186854 224208 186938
rect 223888 186618 223930 186854
rect 224166 186618 224208 186854
rect 223888 186586 224208 186618
rect 254608 187174 254928 187206
rect 254608 186938 254650 187174
rect 254886 186938 254928 187174
rect 254608 186854 254928 186938
rect 254608 186618 254650 186854
rect 254886 186618 254928 186854
rect 254608 186586 254928 186618
rect 285328 187174 285648 187206
rect 285328 186938 285370 187174
rect 285606 186938 285648 187174
rect 285328 186854 285648 186938
rect 285328 186618 285370 186854
rect 285606 186618 285648 186854
rect 285328 186586 285648 186618
rect 316048 187174 316368 187206
rect 316048 186938 316090 187174
rect 316326 186938 316368 187174
rect 316048 186854 316368 186938
rect 316048 186618 316090 186854
rect 316326 186618 316368 186854
rect 316048 186586 316368 186618
rect 54928 183454 55248 183486
rect 54928 183218 54970 183454
rect 55206 183218 55248 183454
rect 54928 183134 55248 183218
rect 54928 182898 54970 183134
rect 55206 182898 55248 183134
rect 54928 182866 55248 182898
rect 85648 183454 85968 183486
rect 85648 183218 85690 183454
rect 85926 183218 85968 183454
rect 85648 183134 85968 183218
rect 85648 182898 85690 183134
rect 85926 182898 85968 183134
rect 85648 182866 85968 182898
rect 116368 183454 116688 183486
rect 116368 183218 116410 183454
rect 116646 183218 116688 183454
rect 116368 183134 116688 183218
rect 116368 182898 116410 183134
rect 116646 182898 116688 183134
rect 116368 182866 116688 182898
rect 147088 183454 147408 183486
rect 147088 183218 147130 183454
rect 147366 183218 147408 183454
rect 147088 183134 147408 183218
rect 147088 182898 147130 183134
rect 147366 182898 147408 183134
rect 147088 182866 147408 182898
rect 177808 183454 178128 183486
rect 177808 183218 177850 183454
rect 178086 183218 178128 183454
rect 177808 183134 178128 183218
rect 177808 182898 177850 183134
rect 178086 182898 178128 183134
rect 177808 182866 178128 182898
rect 208528 183454 208848 183486
rect 208528 183218 208570 183454
rect 208806 183218 208848 183454
rect 208528 183134 208848 183218
rect 208528 182898 208570 183134
rect 208806 182898 208848 183134
rect 208528 182866 208848 182898
rect 239248 183454 239568 183486
rect 239248 183218 239290 183454
rect 239526 183218 239568 183454
rect 239248 183134 239568 183218
rect 239248 182898 239290 183134
rect 239526 182898 239568 183134
rect 239248 182866 239568 182898
rect 269968 183454 270288 183486
rect 269968 183218 270010 183454
rect 270246 183218 270288 183454
rect 269968 183134 270288 183218
rect 269968 182898 270010 183134
rect 270246 182898 270288 183134
rect 269968 182866 270288 182898
rect 300688 183454 301008 183486
rect 300688 183218 300730 183454
rect 300966 183218 301008 183454
rect 300688 183134 301008 183218
rect 300688 182898 300730 183134
rect 300966 182898 301008 183134
rect 300688 182866 301008 182898
rect 331408 183454 331728 183486
rect 331408 183218 331450 183454
rect 331686 183218 331728 183454
rect 331408 183134 331728 183218
rect 331408 182898 331450 183134
rect 331686 182898 331728 183134
rect 331408 182866 331728 182898
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 344394 166054 345014 201498
rect 348114 205774 348734 241218
rect 348114 205538 348146 205774
rect 348382 205538 348466 205774
rect 348702 205538 348734 205774
rect 348114 205454 348734 205538
rect 348114 205218 348146 205454
rect 348382 205218 348466 205454
rect 348702 205218 348734 205454
rect 346768 187174 347088 187206
rect 346768 186938 346810 187174
rect 347046 186938 347088 187174
rect 346768 186854 347088 186938
rect 346768 186618 346810 186854
rect 347046 186618 347088 186854
rect 346768 186586 347088 186618
rect 344394 165818 344426 166054
rect 344662 165818 344746 166054
rect 344982 165818 345014 166054
rect 344394 165734 345014 165818
rect 344394 165498 344426 165734
rect 344662 165498 344746 165734
rect 344982 165498 345014 165734
rect 70288 151174 70608 151206
rect 70288 150938 70330 151174
rect 70566 150938 70608 151174
rect 70288 150854 70608 150938
rect 70288 150618 70330 150854
rect 70566 150618 70608 150854
rect 70288 150586 70608 150618
rect 101008 151174 101328 151206
rect 101008 150938 101050 151174
rect 101286 150938 101328 151174
rect 101008 150854 101328 150938
rect 101008 150618 101050 150854
rect 101286 150618 101328 150854
rect 101008 150586 101328 150618
rect 131728 151174 132048 151206
rect 131728 150938 131770 151174
rect 132006 150938 132048 151174
rect 131728 150854 132048 150938
rect 131728 150618 131770 150854
rect 132006 150618 132048 150854
rect 131728 150586 132048 150618
rect 162448 151174 162768 151206
rect 162448 150938 162490 151174
rect 162726 150938 162768 151174
rect 162448 150854 162768 150938
rect 162448 150618 162490 150854
rect 162726 150618 162768 150854
rect 162448 150586 162768 150618
rect 193168 151174 193488 151206
rect 193168 150938 193210 151174
rect 193446 150938 193488 151174
rect 193168 150854 193488 150938
rect 193168 150618 193210 150854
rect 193446 150618 193488 150854
rect 193168 150586 193488 150618
rect 223888 151174 224208 151206
rect 223888 150938 223930 151174
rect 224166 150938 224208 151174
rect 223888 150854 224208 150938
rect 223888 150618 223930 150854
rect 224166 150618 224208 150854
rect 223888 150586 224208 150618
rect 254608 151174 254928 151206
rect 254608 150938 254650 151174
rect 254886 150938 254928 151174
rect 254608 150854 254928 150938
rect 254608 150618 254650 150854
rect 254886 150618 254928 150854
rect 254608 150586 254928 150618
rect 285328 151174 285648 151206
rect 285328 150938 285370 151174
rect 285606 150938 285648 151174
rect 285328 150854 285648 150938
rect 285328 150618 285370 150854
rect 285606 150618 285648 150854
rect 285328 150586 285648 150618
rect 316048 151174 316368 151206
rect 316048 150938 316090 151174
rect 316326 150938 316368 151174
rect 316048 150854 316368 150938
rect 316048 150618 316090 150854
rect 316326 150618 316368 150854
rect 316048 150586 316368 150618
rect 54928 147454 55248 147486
rect 54928 147218 54970 147454
rect 55206 147218 55248 147454
rect 54928 147134 55248 147218
rect 54928 146898 54970 147134
rect 55206 146898 55248 147134
rect 54928 146866 55248 146898
rect 85648 147454 85968 147486
rect 85648 147218 85690 147454
rect 85926 147218 85968 147454
rect 85648 147134 85968 147218
rect 85648 146898 85690 147134
rect 85926 146898 85968 147134
rect 85648 146866 85968 146898
rect 116368 147454 116688 147486
rect 116368 147218 116410 147454
rect 116646 147218 116688 147454
rect 116368 147134 116688 147218
rect 116368 146898 116410 147134
rect 116646 146898 116688 147134
rect 116368 146866 116688 146898
rect 147088 147454 147408 147486
rect 147088 147218 147130 147454
rect 147366 147218 147408 147454
rect 147088 147134 147408 147218
rect 147088 146898 147130 147134
rect 147366 146898 147408 147134
rect 147088 146866 147408 146898
rect 177808 147454 178128 147486
rect 177808 147218 177850 147454
rect 178086 147218 178128 147454
rect 177808 147134 178128 147218
rect 177808 146898 177850 147134
rect 178086 146898 178128 147134
rect 177808 146866 178128 146898
rect 208528 147454 208848 147486
rect 208528 147218 208570 147454
rect 208806 147218 208848 147454
rect 208528 147134 208848 147218
rect 208528 146898 208570 147134
rect 208806 146898 208848 147134
rect 208528 146866 208848 146898
rect 239248 147454 239568 147486
rect 239248 147218 239290 147454
rect 239526 147218 239568 147454
rect 239248 147134 239568 147218
rect 239248 146898 239290 147134
rect 239526 146898 239568 147134
rect 239248 146866 239568 146898
rect 269968 147454 270288 147486
rect 269968 147218 270010 147454
rect 270246 147218 270288 147454
rect 269968 147134 270288 147218
rect 269968 146898 270010 147134
rect 270246 146898 270288 147134
rect 269968 146866 270288 146898
rect 300688 147454 301008 147486
rect 300688 147218 300730 147454
rect 300966 147218 301008 147454
rect 300688 147134 301008 147218
rect 300688 146898 300730 147134
rect 300966 146898 301008 147134
rect 300688 146866 301008 146898
rect 331408 147454 331728 147486
rect 331408 147218 331450 147454
rect 331686 147218 331728 147454
rect 331408 147134 331728 147218
rect 331408 146898 331450 147134
rect 331686 146898 331728 147134
rect 331408 146866 331728 146898
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 344394 130054 345014 165498
rect 348114 169774 348734 205218
rect 348114 169538 348146 169774
rect 348382 169538 348466 169774
rect 348702 169538 348734 169774
rect 348114 169454 348734 169538
rect 348114 169218 348146 169454
rect 348382 169218 348466 169454
rect 348702 169218 348734 169454
rect 346768 151174 347088 151206
rect 346768 150938 346810 151174
rect 347046 150938 347088 151174
rect 346768 150854 347088 150938
rect 346768 150618 346810 150854
rect 347046 150618 347088 150854
rect 346768 150586 347088 150618
rect 344394 129818 344426 130054
rect 344662 129818 344746 130054
rect 344982 129818 345014 130054
rect 344394 129734 345014 129818
rect 344394 129498 344426 129734
rect 344662 129498 344746 129734
rect 344982 129498 345014 129734
rect 70288 115174 70608 115206
rect 70288 114938 70330 115174
rect 70566 114938 70608 115174
rect 70288 114854 70608 114938
rect 70288 114618 70330 114854
rect 70566 114618 70608 114854
rect 70288 114586 70608 114618
rect 101008 115174 101328 115206
rect 101008 114938 101050 115174
rect 101286 114938 101328 115174
rect 101008 114854 101328 114938
rect 101008 114618 101050 114854
rect 101286 114618 101328 114854
rect 101008 114586 101328 114618
rect 131728 115174 132048 115206
rect 131728 114938 131770 115174
rect 132006 114938 132048 115174
rect 131728 114854 132048 114938
rect 131728 114618 131770 114854
rect 132006 114618 132048 114854
rect 131728 114586 132048 114618
rect 162448 115174 162768 115206
rect 162448 114938 162490 115174
rect 162726 114938 162768 115174
rect 162448 114854 162768 114938
rect 162448 114618 162490 114854
rect 162726 114618 162768 114854
rect 162448 114586 162768 114618
rect 193168 115174 193488 115206
rect 193168 114938 193210 115174
rect 193446 114938 193488 115174
rect 193168 114854 193488 114938
rect 193168 114618 193210 114854
rect 193446 114618 193488 114854
rect 193168 114586 193488 114618
rect 223888 115174 224208 115206
rect 223888 114938 223930 115174
rect 224166 114938 224208 115174
rect 223888 114854 224208 114938
rect 223888 114618 223930 114854
rect 224166 114618 224208 114854
rect 223888 114586 224208 114618
rect 254608 115174 254928 115206
rect 254608 114938 254650 115174
rect 254886 114938 254928 115174
rect 254608 114854 254928 114938
rect 254608 114618 254650 114854
rect 254886 114618 254928 114854
rect 254608 114586 254928 114618
rect 285328 115174 285648 115206
rect 285328 114938 285370 115174
rect 285606 114938 285648 115174
rect 285328 114854 285648 114938
rect 285328 114618 285370 114854
rect 285606 114618 285648 114854
rect 285328 114586 285648 114618
rect 316048 115174 316368 115206
rect 316048 114938 316090 115174
rect 316326 114938 316368 115174
rect 316048 114854 316368 114938
rect 316048 114618 316090 114854
rect 316326 114618 316368 114854
rect 316048 114586 316368 114618
rect 54928 111454 55248 111486
rect 54928 111218 54970 111454
rect 55206 111218 55248 111454
rect 54928 111134 55248 111218
rect 54928 110898 54970 111134
rect 55206 110898 55248 111134
rect 54928 110866 55248 110898
rect 85648 111454 85968 111486
rect 85648 111218 85690 111454
rect 85926 111218 85968 111454
rect 85648 111134 85968 111218
rect 85648 110898 85690 111134
rect 85926 110898 85968 111134
rect 85648 110866 85968 110898
rect 116368 111454 116688 111486
rect 116368 111218 116410 111454
rect 116646 111218 116688 111454
rect 116368 111134 116688 111218
rect 116368 110898 116410 111134
rect 116646 110898 116688 111134
rect 116368 110866 116688 110898
rect 147088 111454 147408 111486
rect 147088 111218 147130 111454
rect 147366 111218 147408 111454
rect 147088 111134 147408 111218
rect 147088 110898 147130 111134
rect 147366 110898 147408 111134
rect 147088 110866 147408 110898
rect 177808 111454 178128 111486
rect 177808 111218 177850 111454
rect 178086 111218 178128 111454
rect 177808 111134 178128 111218
rect 177808 110898 177850 111134
rect 178086 110898 178128 111134
rect 177808 110866 178128 110898
rect 208528 111454 208848 111486
rect 208528 111218 208570 111454
rect 208806 111218 208848 111454
rect 208528 111134 208848 111218
rect 208528 110898 208570 111134
rect 208806 110898 208848 111134
rect 208528 110866 208848 110898
rect 239248 111454 239568 111486
rect 239248 111218 239290 111454
rect 239526 111218 239568 111454
rect 239248 111134 239568 111218
rect 239248 110898 239290 111134
rect 239526 110898 239568 111134
rect 239248 110866 239568 110898
rect 269968 111454 270288 111486
rect 269968 111218 270010 111454
rect 270246 111218 270288 111454
rect 269968 111134 270288 111218
rect 269968 110898 270010 111134
rect 270246 110898 270288 111134
rect 269968 110866 270288 110898
rect 300688 111454 301008 111486
rect 300688 111218 300730 111454
rect 300966 111218 301008 111454
rect 300688 111134 301008 111218
rect 300688 110898 300730 111134
rect 300966 110898 301008 111134
rect 300688 110866 301008 110898
rect 331408 111454 331728 111486
rect 331408 111218 331450 111454
rect 331686 111218 331728 111454
rect 331408 111134 331728 111218
rect 331408 110898 331450 111134
rect 331686 110898 331728 111134
rect 331408 110866 331728 110898
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 344394 94054 345014 129498
rect 348114 133774 348734 169218
rect 348114 133538 348146 133774
rect 348382 133538 348466 133774
rect 348702 133538 348734 133774
rect 348114 133454 348734 133538
rect 348114 133218 348146 133454
rect 348382 133218 348466 133454
rect 348702 133218 348734 133454
rect 346768 115174 347088 115206
rect 346768 114938 346810 115174
rect 347046 114938 347088 115174
rect 346768 114854 347088 114938
rect 346768 114618 346810 114854
rect 347046 114618 347088 114854
rect 346768 114586 347088 114618
rect 344394 93818 344426 94054
rect 344662 93818 344746 94054
rect 344982 93818 345014 94054
rect 344394 93734 345014 93818
rect 344394 93498 344426 93734
rect 344662 93498 344746 93734
rect 344982 93498 345014 93734
rect 70288 79174 70608 79206
rect 70288 78938 70330 79174
rect 70566 78938 70608 79174
rect 70288 78854 70608 78938
rect 70288 78618 70330 78854
rect 70566 78618 70608 78854
rect 70288 78586 70608 78618
rect 101008 79174 101328 79206
rect 101008 78938 101050 79174
rect 101286 78938 101328 79174
rect 101008 78854 101328 78938
rect 101008 78618 101050 78854
rect 101286 78618 101328 78854
rect 101008 78586 101328 78618
rect 131728 79174 132048 79206
rect 131728 78938 131770 79174
rect 132006 78938 132048 79174
rect 131728 78854 132048 78938
rect 131728 78618 131770 78854
rect 132006 78618 132048 78854
rect 131728 78586 132048 78618
rect 162448 79174 162768 79206
rect 162448 78938 162490 79174
rect 162726 78938 162768 79174
rect 162448 78854 162768 78938
rect 162448 78618 162490 78854
rect 162726 78618 162768 78854
rect 162448 78586 162768 78618
rect 193168 79174 193488 79206
rect 193168 78938 193210 79174
rect 193446 78938 193488 79174
rect 193168 78854 193488 78938
rect 193168 78618 193210 78854
rect 193446 78618 193488 78854
rect 193168 78586 193488 78618
rect 223888 79174 224208 79206
rect 223888 78938 223930 79174
rect 224166 78938 224208 79174
rect 223888 78854 224208 78938
rect 223888 78618 223930 78854
rect 224166 78618 224208 78854
rect 223888 78586 224208 78618
rect 254608 79174 254928 79206
rect 254608 78938 254650 79174
rect 254886 78938 254928 79174
rect 254608 78854 254928 78938
rect 254608 78618 254650 78854
rect 254886 78618 254928 78854
rect 254608 78586 254928 78618
rect 285328 79174 285648 79206
rect 285328 78938 285370 79174
rect 285606 78938 285648 79174
rect 285328 78854 285648 78938
rect 285328 78618 285370 78854
rect 285606 78618 285648 78854
rect 285328 78586 285648 78618
rect 316048 79174 316368 79206
rect 316048 78938 316090 79174
rect 316326 78938 316368 79174
rect 316048 78854 316368 78938
rect 316048 78618 316090 78854
rect 316326 78618 316368 78854
rect 316048 78586 316368 78618
rect 54928 75454 55248 75486
rect 54928 75218 54970 75454
rect 55206 75218 55248 75454
rect 54928 75134 55248 75218
rect 54928 74898 54970 75134
rect 55206 74898 55248 75134
rect 54928 74866 55248 74898
rect 85648 75454 85968 75486
rect 85648 75218 85690 75454
rect 85926 75218 85968 75454
rect 85648 75134 85968 75218
rect 85648 74898 85690 75134
rect 85926 74898 85968 75134
rect 85648 74866 85968 74898
rect 116368 75454 116688 75486
rect 116368 75218 116410 75454
rect 116646 75218 116688 75454
rect 116368 75134 116688 75218
rect 116368 74898 116410 75134
rect 116646 74898 116688 75134
rect 116368 74866 116688 74898
rect 147088 75454 147408 75486
rect 147088 75218 147130 75454
rect 147366 75218 147408 75454
rect 147088 75134 147408 75218
rect 147088 74898 147130 75134
rect 147366 74898 147408 75134
rect 147088 74866 147408 74898
rect 177808 75454 178128 75486
rect 177808 75218 177850 75454
rect 178086 75218 178128 75454
rect 177808 75134 178128 75218
rect 177808 74898 177850 75134
rect 178086 74898 178128 75134
rect 177808 74866 178128 74898
rect 208528 75454 208848 75486
rect 208528 75218 208570 75454
rect 208806 75218 208848 75454
rect 208528 75134 208848 75218
rect 208528 74898 208570 75134
rect 208806 74898 208848 75134
rect 208528 74866 208848 74898
rect 239248 75454 239568 75486
rect 239248 75218 239290 75454
rect 239526 75218 239568 75454
rect 239248 75134 239568 75218
rect 239248 74898 239290 75134
rect 239526 74898 239568 75134
rect 239248 74866 239568 74898
rect 269968 75454 270288 75486
rect 269968 75218 270010 75454
rect 270246 75218 270288 75454
rect 269968 75134 270288 75218
rect 269968 74898 270010 75134
rect 270246 74898 270288 75134
rect 269968 74866 270288 74898
rect 300688 75454 301008 75486
rect 300688 75218 300730 75454
rect 300966 75218 301008 75454
rect 300688 75134 301008 75218
rect 300688 74898 300730 75134
rect 300966 74898 301008 75134
rect 300688 74866 301008 74898
rect 331408 75454 331728 75486
rect 331408 75218 331450 75454
rect 331686 75218 331728 75454
rect 331408 75134 331728 75218
rect 331408 74898 331450 75134
rect 331686 74898 331728 75134
rect 331408 74866 331728 74898
rect 344394 58054 345014 93498
rect 348114 97774 348734 133218
rect 348114 97538 348146 97774
rect 348382 97538 348466 97774
rect 348702 97538 348734 97774
rect 348114 97454 348734 97538
rect 348114 97218 348146 97454
rect 348382 97218 348466 97454
rect 348702 97218 348734 97454
rect 346768 79174 347088 79206
rect 346768 78938 346810 79174
rect 347046 78938 347088 79174
rect 346768 78854 347088 78938
rect 346768 78618 346810 78854
rect 347046 78618 347088 78854
rect 346768 78586 347088 78618
rect 344394 57818 344426 58054
rect 344662 57818 344746 58054
rect 344982 57818 345014 58054
rect 344394 57734 345014 57818
rect 344394 57498 344426 57734
rect 344662 57498 344746 57734
rect 344982 57498 345014 57734
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 48954 -3226 49574 14058
rect 48954 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 49574 -3226
rect 48954 -3546 49574 -3462
rect 48954 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 49574 -3546
rect 48954 -7654 49574 -3782
rect 52674 54334 53294 56303
rect 52674 54098 52706 54334
rect 52942 54098 53026 54334
rect 53262 54098 53294 54334
rect 52674 54014 53294 54098
rect 52674 53778 52706 54014
rect 52942 53778 53026 54014
rect 53262 53778 53294 54014
rect 52674 18334 53294 53778
rect 52674 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 53294 18334
rect 52674 18014 53294 18098
rect 52674 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 53294 18014
rect 52674 -4186 53294 17778
rect 52674 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 53294 -4186
rect 52674 -4506 53294 -4422
rect 52674 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 53294 -4506
rect 52674 -7654 53294 -4742
rect 56394 22054 57014 56303
rect 56394 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 57014 22054
rect 56394 21734 57014 21818
rect 56394 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 57014 21734
rect 56394 -5146 57014 21498
rect 56394 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 57014 -5146
rect 56394 -5466 57014 -5382
rect 56394 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 57014 -5466
rect 56394 -7654 57014 -5702
rect 60114 25774 60734 56303
rect 60114 25538 60146 25774
rect 60382 25538 60466 25774
rect 60702 25538 60734 25774
rect 60114 25454 60734 25538
rect 60114 25218 60146 25454
rect 60382 25218 60466 25454
rect 60702 25218 60734 25454
rect 60114 -6106 60734 25218
rect 60114 -6342 60146 -6106
rect 60382 -6342 60466 -6106
rect 60702 -6342 60734 -6106
rect 60114 -6426 60734 -6342
rect 60114 -6662 60146 -6426
rect 60382 -6662 60466 -6426
rect 60702 -6662 60734 -6426
rect 60114 -7654 60734 -6662
rect 63834 29494 64454 56303
rect 63834 29258 63866 29494
rect 64102 29258 64186 29494
rect 64422 29258 64454 29494
rect 63834 29174 64454 29258
rect 63834 28938 63866 29174
rect 64102 28938 64186 29174
rect 64422 28938 64454 29174
rect 63834 -7066 64454 28938
rect 63834 -7302 63866 -7066
rect 64102 -7302 64186 -7066
rect 64422 -7302 64454 -7066
rect 63834 -7386 64454 -7302
rect 63834 -7622 63866 -7386
rect 64102 -7622 64186 -7386
rect 64422 -7622 64454 -7386
rect 63834 -7654 64454 -7622
rect 73794 39454 74414 56303
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 77514 43174 78134 56303
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -1306 78134 6618
rect 77514 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 78134 -1306
rect 77514 -1626 78134 -1542
rect 77514 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 78134 -1626
rect 77514 -7654 78134 -1862
rect 81234 46894 81854 56303
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -2266 81854 10338
rect 81234 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 81854 -2266
rect 81234 -2586 81854 -2502
rect 81234 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 81854 -2586
rect 81234 -7654 81854 -2822
rect 84954 50614 85574 56303
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 84954 -3226 85574 14058
rect 84954 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 85574 -3226
rect 84954 -3546 85574 -3462
rect 84954 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 85574 -3546
rect 84954 -7654 85574 -3782
rect 88674 54334 89294 56303
rect 88674 54098 88706 54334
rect 88942 54098 89026 54334
rect 89262 54098 89294 54334
rect 88674 54014 89294 54098
rect 88674 53778 88706 54014
rect 88942 53778 89026 54014
rect 89262 53778 89294 54014
rect 88674 18334 89294 53778
rect 88674 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 89294 18334
rect 88674 18014 89294 18098
rect 88674 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 89294 18014
rect 88674 -4186 89294 17778
rect 88674 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 89294 -4186
rect 88674 -4506 89294 -4422
rect 88674 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 89294 -4506
rect 88674 -7654 89294 -4742
rect 92394 22054 93014 56303
rect 92394 21818 92426 22054
rect 92662 21818 92746 22054
rect 92982 21818 93014 22054
rect 92394 21734 93014 21818
rect 92394 21498 92426 21734
rect 92662 21498 92746 21734
rect 92982 21498 93014 21734
rect 92394 -5146 93014 21498
rect 92394 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 93014 -5146
rect 92394 -5466 93014 -5382
rect 92394 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 93014 -5466
rect 92394 -7654 93014 -5702
rect 96114 25774 96734 56303
rect 96114 25538 96146 25774
rect 96382 25538 96466 25774
rect 96702 25538 96734 25774
rect 96114 25454 96734 25538
rect 96114 25218 96146 25454
rect 96382 25218 96466 25454
rect 96702 25218 96734 25454
rect 96114 -6106 96734 25218
rect 96114 -6342 96146 -6106
rect 96382 -6342 96466 -6106
rect 96702 -6342 96734 -6106
rect 96114 -6426 96734 -6342
rect 96114 -6662 96146 -6426
rect 96382 -6662 96466 -6426
rect 96702 -6662 96734 -6426
rect 96114 -7654 96734 -6662
rect 99834 29494 100454 56303
rect 99834 29258 99866 29494
rect 100102 29258 100186 29494
rect 100422 29258 100454 29494
rect 99834 29174 100454 29258
rect 99834 28938 99866 29174
rect 100102 28938 100186 29174
rect 100422 28938 100454 29174
rect 99834 -7066 100454 28938
rect 99834 -7302 99866 -7066
rect 100102 -7302 100186 -7066
rect 100422 -7302 100454 -7066
rect 99834 -7386 100454 -7302
rect 99834 -7622 99866 -7386
rect 100102 -7622 100186 -7386
rect 100422 -7622 100454 -7386
rect 99834 -7654 100454 -7622
rect 109794 39454 110414 56303
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 113514 43174 114134 56303
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -1306 114134 6618
rect 113514 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 114134 -1306
rect 113514 -1626 114134 -1542
rect 113514 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 114134 -1626
rect 113514 -7654 114134 -1862
rect 117234 46894 117854 56303
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -2266 117854 10338
rect 117234 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 117854 -2266
rect 117234 -2586 117854 -2502
rect 117234 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 117854 -2586
rect 117234 -7654 117854 -2822
rect 120954 50614 121574 56303
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 120954 -3226 121574 14058
rect 120954 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 121574 -3226
rect 120954 -3546 121574 -3462
rect 120954 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 121574 -3546
rect 120954 -7654 121574 -3782
rect 124674 54334 125294 56303
rect 124674 54098 124706 54334
rect 124942 54098 125026 54334
rect 125262 54098 125294 54334
rect 124674 54014 125294 54098
rect 124674 53778 124706 54014
rect 124942 53778 125026 54014
rect 125262 53778 125294 54014
rect 124674 18334 125294 53778
rect 124674 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 125294 18334
rect 124674 18014 125294 18098
rect 124674 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 125294 18014
rect 124674 -4186 125294 17778
rect 124674 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 125294 -4186
rect 124674 -4506 125294 -4422
rect 124674 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 125294 -4506
rect 124674 -7654 125294 -4742
rect 128394 22054 129014 56303
rect 128394 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 129014 22054
rect 128394 21734 129014 21818
rect 128394 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 129014 21734
rect 128394 -5146 129014 21498
rect 128394 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 129014 -5146
rect 128394 -5466 129014 -5382
rect 128394 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 129014 -5466
rect 128394 -7654 129014 -5702
rect 132114 25774 132734 56303
rect 132114 25538 132146 25774
rect 132382 25538 132466 25774
rect 132702 25538 132734 25774
rect 132114 25454 132734 25538
rect 132114 25218 132146 25454
rect 132382 25218 132466 25454
rect 132702 25218 132734 25454
rect 132114 -6106 132734 25218
rect 132114 -6342 132146 -6106
rect 132382 -6342 132466 -6106
rect 132702 -6342 132734 -6106
rect 132114 -6426 132734 -6342
rect 132114 -6662 132146 -6426
rect 132382 -6662 132466 -6426
rect 132702 -6662 132734 -6426
rect 132114 -7654 132734 -6662
rect 135834 29494 136454 56303
rect 135834 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 136454 29494
rect 135834 29174 136454 29258
rect 135834 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 136454 29174
rect 135834 -7066 136454 28938
rect 135834 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 136454 -7066
rect 135834 -7386 136454 -7302
rect 135834 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 136454 -7386
rect 135834 -7654 136454 -7622
rect 145794 39454 146414 56303
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 149514 43174 150134 56303
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -1306 150134 6618
rect 149514 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 150134 -1306
rect 149514 -1626 150134 -1542
rect 149514 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 150134 -1626
rect 149514 -7654 150134 -1862
rect 153234 46894 153854 56303
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -2266 153854 10338
rect 153234 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 153854 -2266
rect 153234 -2586 153854 -2502
rect 153234 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 153854 -2586
rect 153234 -7654 153854 -2822
rect 156954 50614 157574 56303
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 156954 -3226 157574 14058
rect 156954 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 157574 -3226
rect 156954 -3546 157574 -3462
rect 156954 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 157574 -3546
rect 156954 -7654 157574 -3782
rect 160674 54334 161294 56303
rect 160674 54098 160706 54334
rect 160942 54098 161026 54334
rect 161262 54098 161294 54334
rect 160674 54014 161294 54098
rect 160674 53778 160706 54014
rect 160942 53778 161026 54014
rect 161262 53778 161294 54014
rect 160674 18334 161294 53778
rect 160674 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 161294 18334
rect 160674 18014 161294 18098
rect 160674 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 161294 18014
rect 160674 -4186 161294 17778
rect 160674 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 161294 -4186
rect 160674 -4506 161294 -4422
rect 160674 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 161294 -4506
rect 160674 -7654 161294 -4742
rect 164394 22054 165014 56303
rect 164394 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 165014 22054
rect 164394 21734 165014 21818
rect 164394 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 165014 21734
rect 164394 -5146 165014 21498
rect 164394 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 165014 -5146
rect 164394 -5466 165014 -5382
rect 164394 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 165014 -5466
rect 164394 -7654 165014 -5702
rect 168114 25774 168734 56303
rect 168114 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 168734 25774
rect 168114 25454 168734 25538
rect 168114 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 168734 25454
rect 168114 -6106 168734 25218
rect 168114 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 168734 -6106
rect 168114 -6426 168734 -6342
rect 168114 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 168734 -6426
rect 168114 -7654 168734 -6662
rect 171834 29494 172454 56303
rect 171834 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 172454 29494
rect 171834 29174 172454 29258
rect 171834 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 172454 29174
rect 171834 -7066 172454 28938
rect 171834 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 172454 -7066
rect 171834 -7386 172454 -7302
rect 171834 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 172454 -7386
rect 171834 -7654 172454 -7622
rect 181794 39454 182414 56303
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 185514 43174 186134 56303
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -1306 186134 6618
rect 185514 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 186134 -1306
rect 185514 -1626 186134 -1542
rect 185514 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 186134 -1626
rect 185514 -7654 186134 -1862
rect 189234 46894 189854 56303
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 196674 54334 197294 56303
rect 196674 54098 196706 54334
rect 196942 54098 197026 54334
rect 197262 54098 197294 54334
rect 196674 54014 197294 54098
rect 196674 53778 196706 54014
rect 196942 53778 197026 54014
rect 197262 53778 197294 54014
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -2266 189854 10338
rect 189234 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 189854 -2266
rect 189234 -2586 189854 -2502
rect 189234 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 189854 -2586
rect 189234 -7654 189854 -2822
rect 192954 14614 193574 45068
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 192954 -3226 193574 14058
rect 192954 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 193574 -3226
rect 192954 -3546 193574 -3462
rect 192954 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 193574 -3546
rect 192954 -7654 193574 -3782
rect 196674 18334 197294 53778
rect 196674 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 197294 18334
rect 196674 18014 197294 18098
rect 196674 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 197294 18014
rect 196674 -4186 197294 17778
rect 196674 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 197294 -4186
rect 196674 -4506 197294 -4422
rect 196674 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 197294 -4506
rect 196674 -7654 197294 -4742
rect 200394 22054 201014 56303
rect 200394 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 201014 22054
rect 200394 21734 201014 21818
rect 200394 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 201014 21734
rect 200394 -5146 201014 21498
rect 200394 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 201014 -5146
rect 200394 -5466 201014 -5382
rect 200394 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 201014 -5466
rect 200394 -7654 201014 -5702
rect 204114 25774 204734 56303
rect 204114 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 204734 25774
rect 204114 25454 204734 25538
rect 204114 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 204734 25454
rect 204114 -6106 204734 25218
rect 204114 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 204734 -6106
rect 204114 -6426 204734 -6342
rect 204114 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 204734 -6426
rect 204114 -7654 204734 -6662
rect 207834 29494 208454 56303
rect 207834 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 208454 29494
rect 207834 29174 208454 29258
rect 207834 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 208454 29174
rect 207834 -7066 208454 28938
rect 207834 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 208454 -7066
rect 207834 -7386 208454 -7302
rect 207834 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 208454 -7386
rect 207834 -7654 208454 -7622
rect 217794 39454 218414 56303
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 221514 43174 222134 56303
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -1306 222134 6618
rect 221514 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 222134 -1306
rect 221514 -1626 222134 -1542
rect 221514 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 222134 -1626
rect 221514 -7654 222134 -1862
rect 225234 46894 225854 56303
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -2266 225854 10338
rect 225234 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 225854 -2266
rect 225234 -2586 225854 -2502
rect 225234 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 225854 -2586
rect 225234 -7654 225854 -2822
rect 228954 50614 229574 56303
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 228954 -3226 229574 14058
rect 228954 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 229574 -3226
rect 228954 -3546 229574 -3462
rect 228954 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 229574 -3546
rect 228954 -7654 229574 -3782
rect 232674 54334 233294 56303
rect 232674 54098 232706 54334
rect 232942 54098 233026 54334
rect 233262 54098 233294 54334
rect 232674 54014 233294 54098
rect 232674 53778 232706 54014
rect 232942 53778 233026 54014
rect 233262 53778 233294 54014
rect 232674 18334 233294 53778
rect 232674 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 233294 18334
rect 232674 18014 233294 18098
rect 232674 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 233294 18014
rect 232674 -4186 233294 17778
rect 232674 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 233294 -4186
rect 232674 -4506 233294 -4422
rect 232674 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 233294 -4506
rect 232674 -7654 233294 -4742
rect 236394 22054 237014 56303
rect 236394 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 237014 22054
rect 236394 21734 237014 21818
rect 236394 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 237014 21734
rect 236394 -5146 237014 21498
rect 236394 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 237014 -5146
rect 236394 -5466 237014 -5382
rect 236394 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 237014 -5466
rect 236394 -7654 237014 -5702
rect 240114 25774 240734 56303
rect 240114 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 240734 25774
rect 240114 25454 240734 25538
rect 240114 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 240734 25454
rect 240114 -6106 240734 25218
rect 240114 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 240734 -6106
rect 240114 -6426 240734 -6342
rect 240114 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 240734 -6426
rect 240114 -7654 240734 -6662
rect 243834 29494 244454 56303
rect 243834 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 244454 29494
rect 243834 29174 244454 29258
rect 243834 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 244454 29174
rect 243834 -7066 244454 28938
rect 243834 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 244454 -7066
rect 243834 -7386 244454 -7302
rect 243834 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 244454 -7386
rect 243834 -7654 244454 -7622
rect 253794 39454 254414 56303
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 257514 43174 258134 56303
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -1306 258134 6618
rect 257514 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 258134 -1306
rect 257514 -1626 258134 -1542
rect 257514 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 258134 -1626
rect 257514 -7654 258134 -1862
rect 261234 46894 261854 56303
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -2266 261854 10338
rect 261234 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 261854 -2266
rect 261234 -2586 261854 -2502
rect 261234 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 261854 -2586
rect 261234 -7654 261854 -2822
rect 264954 50614 265574 56303
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 264954 -3226 265574 14058
rect 264954 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 265574 -3226
rect 264954 -3546 265574 -3462
rect 264954 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 265574 -3546
rect 264954 -7654 265574 -3782
rect 268674 54334 269294 56303
rect 268674 54098 268706 54334
rect 268942 54098 269026 54334
rect 269262 54098 269294 54334
rect 268674 54014 269294 54098
rect 268674 53778 268706 54014
rect 268942 53778 269026 54014
rect 269262 53778 269294 54014
rect 268674 18334 269294 53778
rect 268674 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 269294 18334
rect 268674 18014 269294 18098
rect 268674 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 269294 18014
rect 268674 -4186 269294 17778
rect 268674 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 269294 -4186
rect 268674 -4506 269294 -4422
rect 268674 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 269294 -4506
rect 268674 -7654 269294 -4742
rect 272394 22054 273014 56303
rect 272394 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 273014 22054
rect 272394 21734 273014 21818
rect 272394 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 273014 21734
rect 272394 -5146 273014 21498
rect 272394 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 273014 -5146
rect 272394 -5466 273014 -5382
rect 272394 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 273014 -5466
rect 272394 -7654 273014 -5702
rect 276114 25774 276734 56303
rect 276114 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 276734 25774
rect 276114 25454 276734 25538
rect 276114 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 276734 25454
rect 276114 -6106 276734 25218
rect 276114 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 276734 -6106
rect 276114 -6426 276734 -6342
rect 276114 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 276734 -6426
rect 276114 -7654 276734 -6662
rect 279834 29494 280454 56303
rect 279834 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 280454 29494
rect 279834 29174 280454 29258
rect 279834 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 280454 29174
rect 279834 -7066 280454 28938
rect 279834 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 280454 -7066
rect 279834 -7386 280454 -7302
rect 279834 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 280454 -7386
rect 279834 -7654 280454 -7622
rect 289794 39454 290414 56303
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 293514 43174 294134 56303
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -1306 294134 6618
rect 293514 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 294134 -1306
rect 293514 -1626 294134 -1542
rect 293514 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 294134 -1626
rect 293514 -7654 294134 -1862
rect 297234 46894 297854 56303
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 304674 54334 305294 56303
rect 304674 54098 304706 54334
rect 304942 54098 305026 54334
rect 305262 54098 305294 54334
rect 304674 54014 305294 54098
rect 304674 53778 304706 54014
rect 304942 53778 305026 54014
rect 305262 53778 305294 54014
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -2266 297854 10338
rect 297234 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 297854 -2266
rect 297234 -2586 297854 -2502
rect 297234 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 297854 -2586
rect 297234 -7654 297854 -2822
rect 300954 14614 301574 45068
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 300954 -3226 301574 14058
rect 300954 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 301574 -3226
rect 300954 -3546 301574 -3462
rect 300954 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 301574 -3546
rect 300954 -7654 301574 -3782
rect 304674 18334 305294 53778
rect 304674 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 305294 18334
rect 304674 18014 305294 18098
rect 304674 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 305294 18014
rect 304674 -4186 305294 17778
rect 304674 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 305294 -4186
rect 304674 -4506 305294 -4422
rect 304674 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 305294 -4506
rect 304674 -7654 305294 -4742
rect 308394 22054 309014 56303
rect 308394 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 309014 22054
rect 308394 21734 309014 21818
rect 308394 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 309014 21734
rect 308394 -5146 309014 21498
rect 308394 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 309014 -5146
rect 308394 -5466 309014 -5382
rect 308394 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 309014 -5466
rect 308394 -7654 309014 -5702
rect 312114 25774 312734 56303
rect 312114 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 312734 25774
rect 312114 25454 312734 25538
rect 312114 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 312734 25454
rect 312114 -6106 312734 25218
rect 312114 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 312734 -6106
rect 312114 -6426 312734 -6342
rect 312114 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 312734 -6426
rect 312114 -7654 312734 -6662
rect 315834 29494 316454 45068
rect 315834 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 316454 29494
rect 315834 29174 316454 29258
rect 315834 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 316454 29174
rect 315834 -7066 316454 28938
rect 315834 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 316454 -7066
rect 315834 -7386 316454 -7302
rect 315834 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 316454 -7386
rect 315834 -7654 316454 -7622
rect 325794 39454 326414 56303
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 329514 43174 330134 56303
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -1306 330134 6618
rect 329514 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 330134 -1306
rect 329514 -1626 330134 -1542
rect 329514 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 330134 -1626
rect 329514 -7654 330134 -1862
rect 333234 46894 333854 56303
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -2266 333854 10338
rect 333234 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 333854 -2266
rect 333234 -2586 333854 -2502
rect 333234 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 333854 -2586
rect 333234 -7654 333854 -2822
rect 336954 50614 337574 56303
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 336954 -3226 337574 14058
rect 336954 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 337574 -3226
rect 336954 -3546 337574 -3462
rect 336954 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 337574 -3546
rect 336954 -7654 337574 -3782
rect 340674 54334 341294 56303
rect 340674 54098 340706 54334
rect 340942 54098 341026 54334
rect 341262 54098 341294 54334
rect 340674 54014 341294 54098
rect 340674 53778 340706 54014
rect 340942 53778 341026 54014
rect 341262 53778 341294 54014
rect 340674 18334 341294 53778
rect 340674 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 341294 18334
rect 340674 18014 341294 18098
rect 340674 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 341294 18014
rect 340674 -4186 341294 17778
rect 340674 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 341294 -4186
rect 340674 -4506 341294 -4422
rect 340674 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 341294 -4506
rect 340674 -7654 341294 -4742
rect 344394 22054 345014 57498
rect 344394 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 345014 22054
rect 344394 21734 345014 21818
rect 344394 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 345014 21734
rect 344394 -5146 345014 21498
rect 344394 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 345014 -5146
rect 344394 -5466 345014 -5382
rect 344394 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 345014 -5466
rect 344394 -7654 345014 -5702
rect 348114 61774 348734 97218
rect 348114 61538 348146 61774
rect 348382 61538 348466 61774
rect 348702 61538 348734 61774
rect 348114 61454 348734 61538
rect 348114 61218 348146 61454
rect 348382 61218 348466 61454
rect 348702 61218 348734 61454
rect 348114 25774 348734 61218
rect 348114 25538 348146 25774
rect 348382 25538 348466 25774
rect 348702 25538 348734 25774
rect 348114 25454 348734 25538
rect 348114 25218 348146 25454
rect 348382 25218 348466 25454
rect 348702 25218 348734 25454
rect 348114 -6106 348734 25218
rect 348114 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 348734 -6106
rect 348114 -6426 348734 -6342
rect 348114 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 348734 -6426
rect 348114 -7654 348734 -6662
rect 351834 711558 352454 711590
rect 351834 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 352454 711558
rect 351834 711238 352454 711322
rect 351834 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 352454 711238
rect 351834 677494 352454 711002
rect 351834 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 352454 677494
rect 351834 677174 352454 677258
rect 351834 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 352454 677174
rect 351834 641494 352454 676938
rect 351834 641258 351866 641494
rect 352102 641258 352186 641494
rect 352422 641258 352454 641494
rect 351834 641174 352454 641258
rect 351834 640938 351866 641174
rect 352102 640938 352186 641174
rect 352422 640938 352454 641174
rect 351834 605494 352454 640938
rect 351834 605258 351866 605494
rect 352102 605258 352186 605494
rect 352422 605258 352454 605494
rect 351834 605174 352454 605258
rect 351834 604938 351866 605174
rect 352102 604938 352186 605174
rect 352422 604938 352454 605174
rect 351834 569494 352454 604938
rect 351834 569258 351866 569494
rect 352102 569258 352186 569494
rect 352422 569258 352454 569494
rect 351834 569174 352454 569258
rect 351834 568938 351866 569174
rect 352102 568938 352186 569174
rect 352422 568938 352454 569174
rect 351834 533494 352454 568938
rect 351834 533258 351866 533494
rect 352102 533258 352186 533494
rect 352422 533258 352454 533494
rect 351834 533174 352454 533258
rect 351834 532938 351866 533174
rect 352102 532938 352186 533174
rect 352422 532938 352454 533174
rect 351834 497494 352454 532938
rect 351834 497258 351866 497494
rect 352102 497258 352186 497494
rect 352422 497258 352454 497494
rect 351834 497174 352454 497258
rect 351834 496938 351866 497174
rect 352102 496938 352186 497174
rect 352422 496938 352454 497174
rect 351834 461494 352454 496938
rect 351834 461258 351866 461494
rect 352102 461258 352186 461494
rect 352422 461258 352454 461494
rect 351834 461174 352454 461258
rect 351834 460938 351866 461174
rect 352102 460938 352186 461174
rect 352422 460938 352454 461174
rect 351834 425494 352454 460938
rect 351834 425258 351866 425494
rect 352102 425258 352186 425494
rect 352422 425258 352454 425494
rect 351834 425174 352454 425258
rect 351834 424938 351866 425174
rect 352102 424938 352186 425174
rect 352422 424938 352454 425174
rect 351834 389494 352454 424938
rect 351834 389258 351866 389494
rect 352102 389258 352186 389494
rect 352422 389258 352454 389494
rect 351834 389174 352454 389258
rect 351834 388938 351866 389174
rect 352102 388938 352186 389174
rect 352422 388938 352454 389174
rect 351834 353494 352454 388938
rect 351834 353258 351866 353494
rect 352102 353258 352186 353494
rect 352422 353258 352454 353494
rect 351834 353174 352454 353258
rect 351834 352938 351866 353174
rect 352102 352938 352186 353174
rect 352422 352938 352454 353174
rect 351834 317494 352454 352938
rect 351834 317258 351866 317494
rect 352102 317258 352186 317494
rect 352422 317258 352454 317494
rect 351834 317174 352454 317258
rect 351834 316938 351866 317174
rect 352102 316938 352186 317174
rect 352422 316938 352454 317174
rect 351834 281494 352454 316938
rect 351834 281258 351866 281494
rect 352102 281258 352186 281494
rect 352422 281258 352454 281494
rect 351834 281174 352454 281258
rect 351834 280938 351866 281174
rect 352102 280938 352186 281174
rect 352422 280938 352454 281174
rect 351834 245494 352454 280938
rect 351834 245258 351866 245494
rect 352102 245258 352186 245494
rect 352422 245258 352454 245494
rect 351834 245174 352454 245258
rect 351834 244938 351866 245174
rect 352102 244938 352186 245174
rect 352422 244938 352454 245174
rect 351834 209494 352454 244938
rect 351834 209258 351866 209494
rect 352102 209258 352186 209494
rect 352422 209258 352454 209494
rect 351834 209174 352454 209258
rect 351834 208938 351866 209174
rect 352102 208938 352186 209174
rect 352422 208938 352454 209174
rect 351834 173494 352454 208938
rect 351834 173258 351866 173494
rect 352102 173258 352186 173494
rect 352422 173258 352454 173494
rect 351834 173174 352454 173258
rect 351834 172938 351866 173174
rect 352102 172938 352186 173174
rect 352422 172938 352454 173174
rect 351834 137494 352454 172938
rect 351834 137258 351866 137494
rect 352102 137258 352186 137494
rect 352422 137258 352454 137494
rect 351834 137174 352454 137258
rect 351834 136938 351866 137174
rect 352102 136938 352186 137174
rect 352422 136938 352454 137174
rect 351834 101494 352454 136938
rect 351834 101258 351866 101494
rect 352102 101258 352186 101494
rect 352422 101258 352454 101494
rect 351834 101174 352454 101258
rect 351834 100938 351866 101174
rect 352102 100938 352186 101174
rect 352422 100938 352454 101174
rect 351834 65494 352454 100938
rect 351834 65258 351866 65494
rect 352102 65258 352186 65494
rect 352422 65258 352454 65494
rect 351834 65174 352454 65258
rect 351834 64938 351866 65174
rect 352102 64938 352186 65174
rect 352422 64938 352454 65174
rect 351834 29494 352454 64938
rect 351834 29258 351866 29494
rect 352102 29258 352186 29494
rect 352422 29258 352454 29494
rect 351834 29174 352454 29258
rect 351834 28938 351866 29174
rect 352102 28938 352186 29174
rect 352422 28938 352454 29174
rect 351834 -7066 352454 28938
rect 351834 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 352454 -7066
rect 351834 -7386 352454 -7302
rect 351834 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 352454 -7386
rect 351834 -7654 352454 -7622
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 365514 705798 366134 711590
rect 365514 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 366134 705798
rect 365514 705478 366134 705562
rect 365514 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 366134 705478
rect 365514 691174 366134 705242
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -1306 366134 6618
rect 365514 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 366134 -1306
rect 365514 -1626 366134 -1542
rect 365514 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 366134 -1626
rect 365514 -7654 366134 -1862
rect 369234 706758 369854 711590
rect 369234 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 369854 706758
rect 369234 706438 369854 706522
rect 369234 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 369854 706438
rect 369234 694894 369854 706202
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -2266 369854 10338
rect 369234 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 369854 -2266
rect 369234 -2586 369854 -2502
rect 369234 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 369854 -2586
rect 369234 -7654 369854 -2822
rect 372954 707718 373574 711590
rect 372954 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 373574 707718
rect 372954 707398 373574 707482
rect 372954 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 373574 707398
rect 372954 698614 373574 707162
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 372954 -3226 373574 14058
rect 372954 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 373574 -3226
rect 372954 -3546 373574 -3462
rect 372954 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 373574 -3546
rect 372954 -7654 373574 -3782
rect 376674 708678 377294 711590
rect 376674 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 377294 708678
rect 376674 708358 377294 708442
rect 376674 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 377294 708358
rect 376674 666334 377294 708122
rect 376674 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 377294 666334
rect 376674 666014 377294 666098
rect 376674 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 377294 666014
rect 376674 630334 377294 665778
rect 376674 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 377294 630334
rect 376674 630014 377294 630098
rect 376674 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 377294 630014
rect 376674 594334 377294 629778
rect 376674 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 377294 594334
rect 376674 594014 377294 594098
rect 376674 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 377294 594014
rect 376674 558334 377294 593778
rect 376674 558098 376706 558334
rect 376942 558098 377026 558334
rect 377262 558098 377294 558334
rect 376674 558014 377294 558098
rect 376674 557778 376706 558014
rect 376942 557778 377026 558014
rect 377262 557778 377294 558014
rect 376674 522334 377294 557778
rect 376674 522098 376706 522334
rect 376942 522098 377026 522334
rect 377262 522098 377294 522334
rect 376674 522014 377294 522098
rect 376674 521778 376706 522014
rect 376942 521778 377026 522014
rect 377262 521778 377294 522014
rect 376674 486334 377294 521778
rect 376674 486098 376706 486334
rect 376942 486098 377026 486334
rect 377262 486098 377294 486334
rect 376674 486014 377294 486098
rect 376674 485778 376706 486014
rect 376942 485778 377026 486014
rect 377262 485778 377294 486014
rect 376674 450334 377294 485778
rect 376674 450098 376706 450334
rect 376942 450098 377026 450334
rect 377262 450098 377294 450334
rect 376674 450014 377294 450098
rect 376674 449778 376706 450014
rect 376942 449778 377026 450014
rect 377262 449778 377294 450014
rect 376674 414334 377294 449778
rect 376674 414098 376706 414334
rect 376942 414098 377026 414334
rect 377262 414098 377294 414334
rect 376674 414014 377294 414098
rect 376674 413778 376706 414014
rect 376942 413778 377026 414014
rect 377262 413778 377294 414014
rect 376674 378334 377294 413778
rect 376674 378098 376706 378334
rect 376942 378098 377026 378334
rect 377262 378098 377294 378334
rect 376674 378014 377294 378098
rect 376674 377778 376706 378014
rect 376942 377778 377026 378014
rect 377262 377778 377294 378014
rect 376674 342334 377294 377778
rect 376674 342098 376706 342334
rect 376942 342098 377026 342334
rect 377262 342098 377294 342334
rect 376674 342014 377294 342098
rect 376674 341778 376706 342014
rect 376942 341778 377026 342014
rect 377262 341778 377294 342014
rect 376674 306334 377294 341778
rect 376674 306098 376706 306334
rect 376942 306098 377026 306334
rect 377262 306098 377294 306334
rect 376674 306014 377294 306098
rect 376674 305778 376706 306014
rect 376942 305778 377026 306014
rect 377262 305778 377294 306014
rect 376674 270334 377294 305778
rect 376674 270098 376706 270334
rect 376942 270098 377026 270334
rect 377262 270098 377294 270334
rect 376674 270014 377294 270098
rect 376674 269778 376706 270014
rect 376942 269778 377026 270014
rect 377262 269778 377294 270014
rect 376674 234334 377294 269778
rect 376674 234098 376706 234334
rect 376942 234098 377026 234334
rect 377262 234098 377294 234334
rect 376674 234014 377294 234098
rect 376674 233778 376706 234014
rect 376942 233778 377026 234014
rect 377262 233778 377294 234014
rect 376674 198334 377294 233778
rect 376674 198098 376706 198334
rect 376942 198098 377026 198334
rect 377262 198098 377294 198334
rect 376674 198014 377294 198098
rect 376674 197778 376706 198014
rect 376942 197778 377026 198014
rect 377262 197778 377294 198014
rect 376674 162334 377294 197778
rect 376674 162098 376706 162334
rect 376942 162098 377026 162334
rect 377262 162098 377294 162334
rect 376674 162014 377294 162098
rect 376674 161778 376706 162014
rect 376942 161778 377026 162014
rect 377262 161778 377294 162014
rect 376674 126334 377294 161778
rect 376674 126098 376706 126334
rect 376942 126098 377026 126334
rect 377262 126098 377294 126334
rect 376674 126014 377294 126098
rect 376674 125778 376706 126014
rect 376942 125778 377026 126014
rect 377262 125778 377294 126014
rect 376674 90334 377294 125778
rect 376674 90098 376706 90334
rect 376942 90098 377026 90334
rect 377262 90098 377294 90334
rect 376674 90014 377294 90098
rect 376674 89778 376706 90014
rect 376942 89778 377026 90014
rect 377262 89778 377294 90014
rect 376674 54334 377294 89778
rect 376674 54098 376706 54334
rect 376942 54098 377026 54334
rect 377262 54098 377294 54334
rect 376674 54014 377294 54098
rect 376674 53778 376706 54014
rect 376942 53778 377026 54014
rect 377262 53778 377294 54014
rect 376674 18334 377294 53778
rect 376674 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 377294 18334
rect 376674 18014 377294 18098
rect 376674 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 377294 18014
rect 376674 -4186 377294 17778
rect 376674 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 377294 -4186
rect 376674 -4506 377294 -4422
rect 376674 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 377294 -4506
rect 376674 -7654 377294 -4742
rect 380394 709638 381014 711590
rect 380394 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 381014 709638
rect 380394 709318 381014 709402
rect 380394 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 381014 709318
rect 380394 670054 381014 709082
rect 380394 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 381014 670054
rect 380394 669734 381014 669818
rect 380394 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 381014 669734
rect 380394 634054 381014 669498
rect 380394 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 381014 634054
rect 380394 633734 381014 633818
rect 380394 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 381014 633734
rect 380394 598054 381014 633498
rect 380394 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 381014 598054
rect 380394 597734 381014 597818
rect 380394 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 381014 597734
rect 380394 562054 381014 597498
rect 380394 561818 380426 562054
rect 380662 561818 380746 562054
rect 380982 561818 381014 562054
rect 380394 561734 381014 561818
rect 380394 561498 380426 561734
rect 380662 561498 380746 561734
rect 380982 561498 381014 561734
rect 380394 526054 381014 561498
rect 380394 525818 380426 526054
rect 380662 525818 380746 526054
rect 380982 525818 381014 526054
rect 380394 525734 381014 525818
rect 380394 525498 380426 525734
rect 380662 525498 380746 525734
rect 380982 525498 381014 525734
rect 380394 490054 381014 525498
rect 380394 489818 380426 490054
rect 380662 489818 380746 490054
rect 380982 489818 381014 490054
rect 380394 489734 381014 489818
rect 380394 489498 380426 489734
rect 380662 489498 380746 489734
rect 380982 489498 381014 489734
rect 380394 454054 381014 489498
rect 380394 453818 380426 454054
rect 380662 453818 380746 454054
rect 380982 453818 381014 454054
rect 380394 453734 381014 453818
rect 380394 453498 380426 453734
rect 380662 453498 380746 453734
rect 380982 453498 381014 453734
rect 380394 418054 381014 453498
rect 380394 417818 380426 418054
rect 380662 417818 380746 418054
rect 380982 417818 381014 418054
rect 380394 417734 381014 417818
rect 380394 417498 380426 417734
rect 380662 417498 380746 417734
rect 380982 417498 381014 417734
rect 380394 382054 381014 417498
rect 380394 381818 380426 382054
rect 380662 381818 380746 382054
rect 380982 381818 381014 382054
rect 380394 381734 381014 381818
rect 380394 381498 380426 381734
rect 380662 381498 380746 381734
rect 380982 381498 381014 381734
rect 380394 346054 381014 381498
rect 380394 345818 380426 346054
rect 380662 345818 380746 346054
rect 380982 345818 381014 346054
rect 380394 345734 381014 345818
rect 380394 345498 380426 345734
rect 380662 345498 380746 345734
rect 380982 345498 381014 345734
rect 380394 310054 381014 345498
rect 380394 309818 380426 310054
rect 380662 309818 380746 310054
rect 380982 309818 381014 310054
rect 380394 309734 381014 309818
rect 380394 309498 380426 309734
rect 380662 309498 380746 309734
rect 380982 309498 381014 309734
rect 380394 274054 381014 309498
rect 384114 710598 384734 711590
rect 384114 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 384734 710598
rect 384114 710278 384734 710362
rect 384114 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 384734 710278
rect 384114 673774 384734 710042
rect 384114 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 384734 673774
rect 384114 673454 384734 673538
rect 384114 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 384734 673454
rect 384114 637774 384734 673218
rect 384114 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 384734 637774
rect 384114 637454 384734 637538
rect 384114 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 384734 637454
rect 384114 601774 384734 637218
rect 384114 601538 384146 601774
rect 384382 601538 384466 601774
rect 384702 601538 384734 601774
rect 384114 601454 384734 601538
rect 384114 601218 384146 601454
rect 384382 601218 384466 601454
rect 384702 601218 384734 601454
rect 384114 565774 384734 601218
rect 384114 565538 384146 565774
rect 384382 565538 384466 565774
rect 384702 565538 384734 565774
rect 384114 565454 384734 565538
rect 384114 565218 384146 565454
rect 384382 565218 384466 565454
rect 384702 565218 384734 565454
rect 384114 529774 384734 565218
rect 384114 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 384734 529774
rect 384114 529454 384734 529538
rect 384114 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 384734 529454
rect 384114 493774 384734 529218
rect 384114 493538 384146 493774
rect 384382 493538 384466 493774
rect 384702 493538 384734 493774
rect 384114 493454 384734 493538
rect 384114 493218 384146 493454
rect 384382 493218 384466 493454
rect 384702 493218 384734 493454
rect 384114 457774 384734 493218
rect 384114 457538 384146 457774
rect 384382 457538 384466 457774
rect 384702 457538 384734 457774
rect 384114 457454 384734 457538
rect 384114 457218 384146 457454
rect 384382 457218 384466 457454
rect 384702 457218 384734 457454
rect 384114 421774 384734 457218
rect 384114 421538 384146 421774
rect 384382 421538 384466 421774
rect 384702 421538 384734 421774
rect 384114 421454 384734 421538
rect 384114 421218 384146 421454
rect 384382 421218 384466 421454
rect 384702 421218 384734 421454
rect 384114 385774 384734 421218
rect 384114 385538 384146 385774
rect 384382 385538 384466 385774
rect 384702 385538 384734 385774
rect 384114 385454 384734 385538
rect 384114 385218 384146 385454
rect 384382 385218 384466 385454
rect 384702 385218 384734 385454
rect 384114 349774 384734 385218
rect 384114 349538 384146 349774
rect 384382 349538 384466 349774
rect 384702 349538 384734 349774
rect 384114 349454 384734 349538
rect 384114 349218 384146 349454
rect 384382 349218 384466 349454
rect 384702 349218 384734 349454
rect 384114 313774 384734 349218
rect 384114 313538 384146 313774
rect 384382 313538 384466 313774
rect 384702 313538 384734 313774
rect 384114 313454 384734 313538
rect 384114 313218 384146 313454
rect 384382 313218 384466 313454
rect 384702 313218 384734 313454
rect 381491 305828 381557 305829
rect 381491 305764 381492 305828
rect 381556 305764 381557 305828
rect 381491 305763 381557 305764
rect 380394 273818 380426 274054
rect 380662 273818 380746 274054
rect 380982 273818 381014 274054
rect 380394 273734 381014 273818
rect 380394 273498 380426 273734
rect 380662 273498 380746 273734
rect 380982 273498 381014 273734
rect 380394 238054 381014 273498
rect 380394 237818 380426 238054
rect 380662 237818 380746 238054
rect 380982 237818 381014 238054
rect 380394 237734 381014 237818
rect 380394 237498 380426 237734
rect 380662 237498 380746 237734
rect 380982 237498 381014 237734
rect 380394 202054 381014 237498
rect 380394 201818 380426 202054
rect 380662 201818 380746 202054
rect 380982 201818 381014 202054
rect 380394 201734 381014 201818
rect 380394 201498 380426 201734
rect 380662 201498 380746 201734
rect 380982 201498 381014 201734
rect 380394 166054 381014 201498
rect 380394 165818 380426 166054
rect 380662 165818 380746 166054
rect 380982 165818 381014 166054
rect 380394 165734 381014 165818
rect 380394 165498 380426 165734
rect 380662 165498 380746 165734
rect 380982 165498 381014 165734
rect 380394 130054 381014 165498
rect 380394 129818 380426 130054
rect 380662 129818 380746 130054
rect 380982 129818 381014 130054
rect 380394 129734 381014 129818
rect 380394 129498 380426 129734
rect 380662 129498 380746 129734
rect 380982 129498 381014 129734
rect 380394 94054 381014 129498
rect 380394 93818 380426 94054
rect 380662 93818 380746 94054
rect 380982 93818 381014 94054
rect 380394 93734 381014 93818
rect 380394 93498 380426 93734
rect 380662 93498 380746 93734
rect 380982 93498 381014 93734
rect 380394 58054 381014 93498
rect 380394 57818 380426 58054
rect 380662 57818 380746 58054
rect 380982 57818 381014 58054
rect 380394 57734 381014 57818
rect 380394 57498 380426 57734
rect 380662 57498 380746 57734
rect 380982 57498 381014 57734
rect 380394 22054 381014 57498
rect 381494 44845 381554 305763
rect 384114 277774 384734 313218
rect 384114 277538 384146 277774
rect 384382 277538 384466 277774
rect 384702 277538 384734 277774
rect 384114 277454 384734 277538
rect 384114 277218 384146 277454
rect 384382 277218 384466 277454
rect 384702 277218 384734 277454
rect 384114 241774 384734 277218
rect 384114 241538 384146 241774
rect 384382 241538 384466 241774
rect 384702 241538 384734 241774
rect 384114 241454 384734 241538
rect 384114 241218 384146 241454
rect 384382 241218 384466 241454
rect 384702 241218 384734 241454
rect 384114 205774 384734 241218
rect 384114 205538 384146 205774
rect 384382 205538 384466 205774
rect 384702 205538 384734 205774
rect 384114 205454 384734 205538
rect 384114 205218 384146 205454
rect 384382 205218 384466 205454
rect 384702 205218 384734 205454
rect 384114 169774 384734 205218
rect 384114 169538 384146 169774
rect 384382 169538 384466 169774
rect 384702 169538 384734 169774
rect 384114 169454 384734 169538
rect 384114 169218 384146 169454
rect 384382 169218 384466 169454
rect 384702 169218 384734 169454
rect 384114 133774 384734 169218
rect 384114 133538 384146 133774
rect 384382 133538 384466 133774
rect 384702 133538 384734 133774
rect 384114 133454 384734 133538
rect 384114 133218 384146 133454
rect 384382 133218 384466 133454
rect 384702 133218 384734 133454
rect 384114 97774 384734 133218
rect 384114 97538 384146 97774
rect 384382 97538 384466 97774
rect 384702 97538 384734 97774
rect 384114 97454 384734 97538
rect 384114 97218 384146 97454
rect 384382 97218 384466 97454
rect 384702 97218 384734 97454
rect 384114 61774 384734 97218
rect 387834 711558 388454 711590
rect 387834 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 388454 711558
rect 387834 711238 388454 711322
rect 387834 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 388454 711238
rect 387834 677494 388454 711002
rect 387834 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 388454 677494
rect 387834 677174 388454 677258
rect 387834 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 388454 677174
rect 387834 641494 388454 676938
rect 387834 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 388454 641494
rect 387834 641174 388454 641258
rect 387834 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 388454 641174
rect 387834 605494 388454 640938
rect 387834 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 388454 605494
rect 387834 605174 388454 605258
rect 387834 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 388454 605174
rect 387834 569494 388454 604938
rect 387834 569258 387866 569494
rect 388102 569258 388186 569494
rect 388422 569258 388454 569494
rect 387834 569174 388454 569258
rect 387834 568938 387866 569174
rect 388102 568938 388186 569174
rect 388422 568938 388454 569174
rect 387834 533494 388454 568938
rect 387834 533258 387866 533494
rect 388102 533258 388186 533494
rect 388422 533258 388454 533494
rect 387834 533174 388454 533258
rect 387834 532938 387866 533174
rect 388102 532938 388186 533174
rect 388422 532938 388454 533174
rect 387834 497494 388454 532938
rect 387834 497258 387866 497494
rect 388102 497258 388186 497494
rect 388422 497258 388454 497494
rect 387834 497174 388454 497258
rect 387834 496938 387866 497174
rect 388102 496938 388186 497174
rect 388422 496938 388454 497174
rect 387834 461494 388454 496938
rect 387834 461258 387866 461494
rect 388102 461258 388186 461494
rect 388422 461258 388454 461494
rect 387834 461174 388454 461258
rect 387834 460938 387866 461174
rect 388102 460938 388186 461174
rect 388422 460938 388454 461174
rect 387834 425494 388454 460938
rect 387834 425258 387866 425494
rect 388102 425258 388186 425494
rect 388422 425258 388454 425494
rect 387834 425174 388454 425258
rect 387834 424938 387866 425174
rect 388102 424938 388186 425174
rect 388422 424938 388454 425174
rect 387834 389494 388454 424938
rect 387834 389258 387866 389494
rect 388102 389258 388186 389494
rect 388422 389258 388454 389494
rect 387834 389174 388454 389258
rect 387834 388938 387866 389174
rect 388102 388938 388186 389174
rect 388422 388938 388454 389174
rect 387834 353494 388454 388938
rect 387834 353258 387866 353494
rect 388102 353258 388186 353494
rect 388422 353258 388454 353494
rect 387834 353174 388454 353258
rect 387834 352938 387866 353174
rect 388102 352938 388186 353174
rect 388422 352938 388454 353174
rect 387834 317494 388454 352938
rect 387834 317258 387866 317494
rect 388102 317258 388186 317494
rect 388422 317258 388454 317494
rect 387834 317174 388454 317258
rect 387834 316938 387866 317174
rect 388102 316938 388186 317174
rect 388422 316938 388454 317174
rect 387834 281494 388454 316938
rect 387834 281258 387866 281494
rect 388102 281258 388186 281494
rect 388422 281258 388454 281494
rect 387834 281174 388454 281258
rect 387834 280938 387866 281174
rect 388102 280938 388186 281174
rect 388422 280938 388454 281174
rect 387834 245494 388454 280938
rect 387834 245258 387866 245494
rect 388102 245258 388186 245494
rect 388422 245258 388454 245494
rect 387834 245174 388454 245258
rect 387834 244938 387866 245174
rect 388102 244938 388186 245174
rect 388422 244938 388454 245174
rect 387834 209494 388454 244938
rect 387834 209258 387866 209494
rect 388102 209258 388186 209494
rect 388422 209258 388454 209494
rect 387834 209174 388454 209258
rect 387834 208938 387866 209174
rect 388102 208938 388186 209174
rect 388422 208938 388454 209174
rect 387834 173494 388454 208938
rect 387834 173258 387866 173494
rect 388102 173258 388186 173494
rect 388422 173258 388454 173494
rect 387834 173174 388454 173258
rect 387834 172938 387866 173174
rect 388102 172938 388186 173174
rect 388422 172938 388454 173174
rect 387834 137494 388454 172938
rect 387834 137258 387866 137494
rect 388102 137258 388186 137494
rect 388422 137258 388454 137494
rect 387834 137174 388454 137258
rect 387834 136938 387866 137174
rect 388102 136938 388186 137174
rect 388422 136938 388454 137174
rect 387834 101494 388454 136938
rect 387834 101258 387866 101494
rect 388102 101258 388186 101494
rect 388422 101258 388454 101494
rect 387834 101174 388454 101258
rect 387834 100938 387866 101174
rect 388102 100938 388186 101174
rect 388422 100938 388454 101174
rect 387834 92137 388454 100938
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 92137 398414 110898
rect 401514 705798 402134 711590
rect 401514 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 402134 705798
rect 401514 705478 402134 705562
rect 401514 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 402134 705478
rect 401514 691174 402134 705242
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 405234 706758 405854 711590
rect 405234 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 405854 706758
rect 405234 706438 405854 706522
rect 405234 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 405854 706438
rect 405234 694894 405854 706202
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 404417 327454 404737 327486
rect 404417 327218 404459 327454
rect 404695 327218 404737 327454
rect 404417 327134 404737 327218
rect 404417 326898 404459 327134
rect 404695 326898 404737 327134
rect 404417 326866 404737 326898
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 92137 402134 114618
rect 405234 298894 405854 334338
rect 408954 707718 409574 711590
rect 408954 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 409574 707718
rect 408954 707398 409574 707482
rect 408954 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 409574 707398
rect 408954 698614 409574 707162
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 407890 331174 408210 331206
rect 407890 330938 407932 331174
rect 408168 330938 408210 331174
rect 407890 330854 408210 330938
rect 407890 330618 407932 330854
rect 408168 330618 408210 330854
rect 407890 330586 408210 330618
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 104460 405854 118338
rect 408954 302614 409574 338058
rect 412674 708678 413294 711590
rect 412674 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 413294 708678
rect 412674 708358 413294 708442
rect 412674 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 413294 708358
rect 412674 666334 413294 708122
rect 412674 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 413294 666334
rect 412674 666014 413294 666098
rect 412674 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 413294 666014
rect 412674 630334 413294 665778
rect 412674 630098 412706 630334
rect 412942 630098 413026 630334
rect 413262 630098 413294 630334
rect 412674 630014 413294 630098
rect 412674 629778 412706 630014
rect 412942 629778 413026 630014
rect 413262 629778 413294 630014
rect 412674 594334 413294 629778
rect 412674 594098 412706 594334
rect 412942 594098 413026 594334
rect 413262 594098 413294 594334
rect 412674 594014 413294 594098
rect 412674 593778 412706 594014
rect 412942 593778 413026 594014
rect 413262 593778 413294 594014
rect 412674 558334 413294 593778
rect 412674 558098 412706 558334
rect 412942 558098 413026 558334
rect 413262 558098 413294 558334
rect 412674 558014 413294 558098
rect 412674 557778 412706 558014
rect 412942 557778 413026 558014
rect 413262 557778 413294 558014
rect 412674 522334 413294 557778
rect 412674 522098 412706 522334
rect 412942 522098 413026 522334
rect 413262 522098 413294 522334
rect 412674 522014 413294 522098
rect 412674 521778 412706 522014
rect 412942 521778 413026 522014
rect 413262 521778 413294 522014
rect 412674 486334 413294 521778
rect 412674 486098 412706 486334
rect 412942 486098 413026 486334
rect 413262 486098 413294 486334
rect 412674 486014 413294 486098
rect 412674 485778 412706 486014
rect 412942 485778 413026 486014
rect 413262 485778 413294 486014
rect 412674 450334 413294 485778
rect 412674 450098 412706 450334
rect 412942 450098 413026 450334
rect 413262 450098 413294 450334
rect 412674 450014 413294 450098
rect 412674 449778 412706 450014
rect 412942 449778 413026 450014
rect 413262 449778 413294 450014
rect 412674 414334 413294 449778
rect 412674 414098 412706 414334
rect 412942 414098 413026 414334
rect 413262 414098 413294 414334
rect 412674 414014 413294 414098
rect 412674 413778 412706 414014
rect 412942 413778 413026 414014
rect 413262 413778 413294 414014
rect 412674 378334 413294 413778
rect 412674 378098 412706 378334
rect 412942 378098 413026 378334
rect 413262 378098 413294 378334
rect 412674 378014 413294 378098
rect 412674 377778 412706 378014
rect 412942 377778 413026 378014
rect 413262 377778 413294 378014
rect 412674 342334 413294 377778
rect 412674 342098 412706 342334
rect 412942 342098 413026 342334
rect 413262 342098 413294 342334
rect 412674 342014 413294 342098
rect 412674 341778 412706 342014
rect 412942 341778 413026 342014
rect 413262 341778 413294 342014
rect 411363 327454 411683 327486
rect 411363 327218 411405 327454
rect 411641 327218 411683 327454
rect 411363 327134 411683 327218
rect 411363 326898 411405 327134
rect 411641 326898 411683 327134
rect 411363 326866 411683 326898
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 412674 306334 413294 341778
rect 416394 709638 417014 711590
rect 416394 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 417014 709638
rect 416394 709318 417014 709402
rect 416394 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 417014 709318
rect 416394 670054 417014 709082
rect 416394 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 417014 670054
rect 416394 669734 417014 669818
rect 416394 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 417014 669734
rect 416394 634054 417014 669498
rect 416394 633818 416426 634054
rect 416662 633818 416746 634054
rect 416982 633818 417014 634054
rect 416394 633734 417014 633818
rect 416394 633498 416426 633734
rect 416662 633498 416746 633734
rect 416982 633498 417014 633734
rect 416394 598054 417014 633498
rect 416394 597818 416426 598054
rect 416662 597818 416746 598054
rect 416982 597818 417014 598054
rect 416394 597734 417014 597818
rect 416394 597498 416426 597734
rect 416662 597498 416746 597734
rect 416982 597498 417014 597734
rect 416394 562054 417014 597498
rect 416394 561818 416426 562054
rect 416662 561818 416746 562054
rect 416982 561818 417014 562054
rect 416394 561734 417014 561818
rect 416394 561498 416426 561734
rect 416662 561498 416746 561734
rect 416982 561498 417014 561734
rect 416394 526054 417014 561498
rect 416394 525818 416426 526054
rect 416662 525818 416746 526054
rect 416982 525818 417014 526054
rect 416394 525734 417014 525818
rect 416394 525498 416426 525734
rect 416662 525498 416746 525734
rect 416982 525498 417014 525734
rect 416394 490054 417014 525498
rect 416394 489818 416426 490054
rect 416662 489818 416746 490054
rect 416982 489818 417014 490054
rect 416394 489734 417014 489818
rect 416394 489498 416426 489734
rect 416662 489498 416746 489734
rect 416982 489498 417014 489734
rect 416394 454054 417014 489498
rect 416394 453818 416426 454054
rect 416662 453818 416746 454054
rect 416982 453818 417014 454054
rect 416394 453734 417014 453818
rect 416394 453498 416426 453734
rect 416662 453498 416746 453734
rect 416982 453498 417014 453734
rect 416394 418054 417014 453498
rect 416394 417818 416426 418054
rect 416662 417818 416746 418054
rect 416982 417818 417014 418054
rect 416394 417734 417014 417818
rect 416394 417498 416426 417734
rect 416662 417498 416746 417734
rect 416982 417498 417014 417734
rect 416394 382054 417014 417498
rect 416394 381818 416426 382054
rect 416662 381818 416746 382054
rect 416982 381818 417014 382054
rect 416394 381734 417014 381818
rect 416394 381498 416426 381734
rect 416662 381498 416746 381734
rect 416982 381498 417014 381734
rect 416394 346054 417014 381498
rect 416394 345818 416426 346054
rect 416662 345818 416746 346054
rect 416982 345818 417014 346054
rect 416394 345734 417014 345818
rect 416394 345498 416426 345734
rect 416662 345498 416746 345734
rect 416982 345498 417014 345734
rect 414836 331174 415156 331206
rect 414836 330938 414878 331174
rect 415114 330938 415156 331174
rect 414836 330854 415156 330938
rect 414836 330618 414878 330854
rect 415114 330618 415156 330854
rect 414836 330586 415156 330618
rect 412674 306098 412706 306334
rect 412942 306098 413026 306334
rect 413262 306098 413294 306334
rect 412674 306014 413294 306098
rect 412674 305778 412706 306014
rect 412942 305778 413026 306014
rect 413262 305778 413294 306014
rect 412674 270334 413294 305778
rect 412674 270098 412706 270334
rect 412942 270098 413026 270334
rect 413262 270098 413294 270334
rect 412674 270014 413294 270098
rect 412674 269778 412706 270014
rect 412942 269778 413026 270014
rect 413262 269778 413294 270014
rect 412674 234334 413294 269778
rect 412674 234098 412706 234334
rect 412942 234098 413026 234334
rect 413262 234098 413294 234334
rect 412674 234014 413294 234098
rect 412674 233778 412706 234014
rect 412942 233778 413026 234014
rect 413262 233778 413294 234014
rect 412674 198334 413294 233778
rect 412674 198098 412706 198334
rect 412942 198098 413026 198334
rect 413262 198098 413294 198334
rect 412674 198014 413294 198098
rect 412674 197778 412706 198014
rect 412942 197778 413026 198014
rect 413262 197778 413294 198014
rect 412674 162334 413294 197778
rect 412674 162098 412706 162334
rect 412942 162098 413026 162334
rect 413262 162098 413294 162334
rect 412674 162014 413294 162098
rect 412674 161778 412706 162014
rect 412942 161778 413026 162014
rect 413262 161778 413294 162014
rect 412674 161465 413294 161778
rect 416394 310054 417014 345498
rect 420114 710598 420734 711590
rect 420114 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 420734 710598
rect 420114 710278 420734 710362
rect 420114 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 420734 710278
rect 420114 673774 420734 710042
rect 420114 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 420734 673774
rect 420114 673454 420734 673538
rect 420114 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 420734 673454
rect 420114 637774 420734 673218
rect 420114 637538 420146 637774
rect 420382 637538 420466 637774
rect 420702 637538 420734 637774
rect 420114 637454 420734 637538
rect 420114 637218 420146 637454
rect 420382 637218 420466 637454
rect 420702 637218 420734 637454
rect 420114 601774 420734 637218
rect 420114 601538 420146 601774
rect 420382 601538 420466 601774
rect 420702 601538 420734 601774
rect 420114 601454 420734 601538
rect 420114 601218 420146 601454
rect 420382 601218 420466 601454
rect 420702 601218 420734 601454
rect 420114 565774 420734 601218
rect 420114 565538 420146 565774
rect 420382 565538 420466 565774
rect 420702 565538 420734 565774
rect 420114 565454 420734 565538
rect 420114 565218 420146 565454
rect 420382 565218 420466 565454
rect 420702 565218 420734 565454
rect 420114 529774 420734 565218
rect 420114 529538 420146 529774
rect 420382 529538 420466 529774
rect 420702 529538 420734 529774
rect 420114 529454 420734 529538
rect 420114 529218 420146 529454
rect 420382 529218 420466 529454
rect 420702 529218 420734 529454
rect 420114 493774 420734 529218
rect 420114 493538 420146 493774
rect 420382 493538 420466 493774
rect 420702 493538 420734 493774
rect 420114 493454 420734 493538
rect 420114 493218 420146 493454
rect 420382 493218 420466 493454
rect 420702 493218 420734 493454
rect 420114 457774 420734 493218
rect 420114 457538 420146 457774
rect 420382 457538 420466 457774
rect 420702 457538 420734 457774
rect 420114 457454 420734 457538
rect 420114 457218 420146 457454
rect 420382 457218 420466 457454
rect 420702 457218 420734 457454
rect 420114 421774 420734 457218
rect 423834 711558 424454 711590
rect 423834 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 424454 711558
rect 423834 711238 424454 711322
rect 423834 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 424454 711238
rect 423834 677494 424454 711002
rect 423834 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 424454 677494
rect 423834 677174 424454 677258
rect 423834 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 424454 677174
rect 423834 641494 424454 676938
rect 423834 641258 423866 641494
rect 424102 641258 424186 641494
rect 424422 641258 424454 641494
rect 423834 641174 424454 641258
rect 423834 640938 423866 641174
rect 424102 640938 424186 641174
rect 424422 640938 424454 641174
rect 423834 605494 424454 640938
rect 423834 605258 423866 605494
rect 424102 605258 424186 605494
rect 424422 605258 424454 605494
rect 423834 605174 424454 605258
rect 423834 604938 423866 605174
rect 424102 604938 424186 605174
rect 424422 604938 424454 605174
rect 423834 569494 424454 604938
rect 423834 569258 423866 569494
rect 424102 569258 424186 569494
rect 424422 569258 424454 569494
rect 423834 569174 424454 569258
rect 423834 568938 423866 569174
rect 424102 568938 424186 569174
rect 424422 568938 424454 569174
rect 423834 533494 424454 568938
rect 423834 533258 423866 533494
rect 424102 533258 424186 533494
rect 424422 533258 424454 533494
rect 423834 533174 424454 533258
rect 423834 532938 423866 533174
rect 424102 532938 424186 533174
rect 424422 532938 424454 533174
rect 423834 497494 424454 532938
rect 423834 497258 423866 497494
rect 424102 497258 424186 497494
rect 424422 497258 424454 497494
rect 423834 497174 424454 497258
rect 423834 496938 423866 497174
rect 424102 496938 424186 497174
rect 424422 496938 424454 497174
rect 423834 461494 424454 496938
rect 423834 461258 423866 461494
rect 424102 461258 424186 461494
rect 424422 461258 424454 461494
rect 423834 461174 424454 461258
rect 423834 460938 423866 461174
rect 424102 460938 424186 461174
rect 424422 460938 424454 461174
rect 423834 444412 424454 460938
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 443377 434414 470898
rect 437514 705798 438134 711590
rect 437514 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 438134 705798
rect 437514 705478 438134 705562
rect 437514 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 438134 705478
rect 437514 691174 438134 705242
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 444412 438134 474618
rect 441234 706758 441854 711590
rect 441234 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 441854 706758
rect 441234 706438 441854 706522
rect 441234 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 441854 706438
rect 441234 694894 441854 706202
rect 444954 707718 445574 711590
rect 444954 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 445574 707718
rect 444954 707398 445574 707482
rect 444954 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 445574 707398
rect 444235 700500 444301 700501
rect 444235 700436 444236 700500
rect 444300 700436 444301 700500
rect 444235 700435 444301 700436
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 443377 441854 478338
rect 426624 439174 426944 439206
rect 426624 438938 426666 439174
rect 426902 438938 426944 439174
rect 426624 438854 426944 438938
rect 426624 438618 426666 438854
rect 426902 438618 426944 438854
rect 426624 438586 426944 438618
rect 432305 439174 432625 439206
rect 432305 438938 432347 439174
rect 432583 438938 432625 439174
rect 432305 438854 432625 438938
rect 432305 438618 432347 438854
rect 432583 438618 432625 438854
rect 432305 438586 432625 438618
rect 437986 439174 438306 439206
rect 437986 438938 438028 439174
rect 438264 438938 438306 439174
rect 437986 438854 438306 438938
rect 437986 438618 438028 438854
rect 438264 438618 438306 438854
rect 437986 438586 438306 438618
rect 443667 439174 443987 439206
rect 443667 438938 443709 439174
rect 443945 438938 443987 439174
rect 443667 438854 443987 438938
rect 443667 438618 443709 438854
rect 443945 438618 443987 438854
rect 443667 438586 443987 438618
rect 423784 435454 424104 435486
rect 423784 435218 423826 435454
rect 424062 435218 424104 435454
rect 423784 435134 424104 435218
rect 423784 434898 423826 435134
rect 424062 434898 424104 435134
rect 423784 434866 424104 434898
rect 429465 435454 429785 435486
rect 429465 435218 429507 435454
rect 429743 435218 429785 435454
rect 429465 435134 429785 435218
rect 429465 434898 429507 435134
rect 429743 434898 429785 435134
rect 429465 434866 429785 434898
rect 435146 435454 435466 435486
rect 435146 435218 435188 435454
rect 435424 435218 435466 435454
rect 435146 435134 435466 435218
rect 435146 434898 435188 435134
rect 435424 434898 435466 435134
rect 435146 434866 435466 434898
rect 440827 435454 441147 435486
rect 440827 435218 440869 435454
rect 441105 435218 441147 435454
rect 440827 435134 441147 435218
rect 440827 434898 440869 435134
rect 441105 434898 441147 435134
rect 440827 434866 441147 434898
rect 420114 421538 420146 421774
rect 420382 421538 420466 421774
rect 420702 421538 420734 421774
rect 420114 421454 420734 421538
rect 420114 421218 420146 421454
rect 420382 421218 420466 421454
rect 420702 421218 420734 421454
rect 420114 385774 420734 421218
rect 420114 385538 420146 385774
rect 420382 385538 420466 385774
rect 420702 385538 420734 385774
rect 420114 385454 420734 385538
rect 420114 385218 420146 385454
rect 420382 385218 420466 385454
rect 420702 385218 420734 385454
rect 420114 349774 420734 385218
rect 420114 349538 420146 349774
rect 420382 349538 420466 349774
rect 420702 349538 420734 349774
rect 420114 349454 420734 349538
rect 420114 349218 420146 349454
rect 420382 349218 420466 349454
rect 420702 349218 420734 349454
rect 418309 327454 418629 327486
rect 418309 327218 418351 327454
rect 418587 327218 418629 327454
rect 418309 327134 418629 327218
rect 418309 326898 418351 327134
rect 418587 326898 418629 327134
rect 418309 326866 418629 326898
rect 416394 309818 416426 310054
rect 416662 309818 416746 310054
rect 416982 309818 417014 310054
rect 416394 309734 417014 309818
rect 416394 309498 416426 309734
rect 416662 309498 416746 309734
rect 416982 309498 417014 309734
rect 416394 274054 417014 309498
rect 416394 273818 416426 274054
rect 416662 273818 416746 274054
rect 416982 273818 417014 274054
rect 416394 273734 417014 273818
rect 416394 273498 416426 273734
rect 416662 273498 416746 273734
rect 416982 273498 417014 273734
rect 416394 238054 417014 273498
rect 416394 237818 416426 238054
rect 416662 237818 416746 238054
rect 416982 237818 417014 238054
rect 416394 237734 417014 237818
rect 416394 237498 416426 237734
rect 416662 237498 416746 237734
rect 416982 237498 417014 237734
rect 416394 202054 417014 237498
rect 416394 201818 416426 202054
rect 416662 201818 416746 202054
rect 416982 201818 417014 202054
rect 416394 201734 417014 201818
rect 416394 201498 416426 201734
rect 416662 201498 416746 201734
rect 416982 201498 417014 201734
rect 416394 166054 417014 201498
rect 416394 165818 416426 166054
rect 416662 165818 416746 166054
rect 416982 165818 417014 166054
rect 416394 165734 417014 165818
rect 416394 165498 416426 165734
rect 416662 165498 416746 165734
rect 416982 165498 417014 165734
rect 416394 161465 417014 165498
rect 420114 313774 420734 349218
rect 423834 389494 424454 420068
rect 423834 389258 423866 389494
rect 424102 389258 424186 389494
rect 424422 389258 424454 389494
rect 423834 389174 424454 389258
rect 423834 388938 423866 389174
rect 424102 388938 424186 389174
rect 424422 388938 424454 389174
rect 423834 353494 424454 388938
rect 423834 353258 423866 353494
rect 424102 353258 424186 353494
rect 424422 353258 424454 353494
rect 423834 353174 424454 353258
rect 423834 352938 423866 353174
rect 424102 352938 424186 353174
rect 424422 352938 424454 353174
rect 421051 334524 421117 334525
rect 421051 334460 421052 334524
rect 421116 334460 421117 334524
rect 421051 334459 421117 334460
rect 420114 313538 420146 313774
rect 420382 313538 420466 313774
rect 420702 313538 420734 313774
rect 420114 313454 420734 313538
rect 420114 313218 420146 313454
rect 420382 313218 420466 313454
rect 420702 313218 420734 313454
rect 420114 277774 420734 313218
rect 420114 277538 420146 277774
rect 420382 277538 420466 277774
rect 420702 277538 420734 277774
rect 420114 277454 420734 277538
rect 420114 277218 420146 277454
rect 420382 277218 420466 277454
rect 420702 277218 420734 277454
rect 420114 241774 420734 277218
rect 420114 241538 420146 241774
rect 420382 241538 420466 241774
rect 420702 241538 420734 241774
rect 420114 241454 420734 241538
rect 420114 241218 420146 241454
rect 420382 241218 420466 241454
rect 420702 241218 420734 241454
rect 420114 205774 420734 241218
rect 420114 205538 420146 205774
rect 420382 205538 420466 205774
rect 420702 205538 420734 205774
rect 420114 205454 420734 205538
rect 420114 205218 420146 205454
rect 420382 205218 420466 205454
rect 420702 205218 420734 205454
rect 420114 169774 420734 205218
rect 420114 169538 420146 169774
rect 420382 169538 420466 169774
rect 420702 169538 420734 169774
rect 420114 169454 420734 169538
rect 420114 169218 420146 169454
rect 420382 169218 420466 169454
rect 420702 169218 420734 169454
rect 420114 161465 420734 169218
rect 421054 162757 421114 334459
rect 421782 331174 422102 331206
rect 421782 330938 421824 331174
rect 422060 330938 422102 331174
rect 421782 330854 422102 330938
rect 421782 330618 421824 330854
rect 422060 330618 422102 330854
rect 421782 330586 422102 330618
rect 423834 317494 424454 352938
rect 433794 399454 434414 420423
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 428411 334524 428477 334525
rect 428411 334460 428412 334524
rect 428476 334460 428477 334524
rect 428411 334459 428477 334460
rect 425255 327454 425575 327486
rect 425255 327218 425297 327454
rect 425533 327218 425575 327454
rect 425255 327134 425575 327218
rect 425255 326898 425297 327134
rect 425533 326898 425575 327134
rect 425255 326866 425575 326898
rect 423834 317258 423866 317494
rect 424102 317258 424186 317494
rect 424422 317258 424454 317494
rect 423834 317174 424454 317258
rect 423834 316938 423866 317174
rect 424102 316938 424186 317174
rect 424422 316938 424454 317174
rect 423834 281494 424454 316938
rect 423834 281258 423866 281494
rect 424102 281258 424186 281494
rect 424422 281258 424454 281494
rect 423834 281174 424454 281258
rect 423834 280938 423866 281174
rect 424102 280938 424186 281174
rect 424422 280938 424454 281174
rect 423834 245494 424454 280938
rect 423834 245258 423866 245494
rect 424102 245258 424186 245494
rect 424422 245258 424454 245494
rect 423834 245174 424454 245258
rect 423834 244938 423866 245174
rect 424102 244938 424186 245174
rect 424422 244938 424454 245174
rect 423834 209494 424454 244938
rect 423834 209258 423866 209494
rect 424102 209258 424186 209494
rect 424422 209258 424454 209494
rect 423834 209174 424454 209258
rect 423834 208938 423866 209174
rect 424102 208938 424186 209174
rect 424422 208938 424454 209174
rect 423834 173494 424454 208938
rect 423834 173258 423866 173494
rect 424102 173258 424186 173494
rect 424422 173258 424454 173494
rect 423834 173174 424454 173258
rect 423834 172938 423866 173174
rect 424102 172938 424186 173174
rect 424422 172938 424454 173174
rect 421051 162756 421117 162757
rect 421051 162692 421052 162756
rect 421116 162692 421117 162756
rect 421051 162691 421117 162692
rect 423834 161465 424454 172938
rect 428414 162757 428474 334459
rect 428728 331174 429048 331206
rect 428728 330938 428770 331174
rect 429006 330938 429048 331174
rect 428728 330854 429048 330938
rect 428728 330618 428770 330854
rect 429006 330618 429048 330854
rect 428728 330586 429048 330618
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 428411 162756 428477 162757
rect 428411 162692 428412 162756
rect 428476 162692 428477 162756
rect 428411 162691 428477 162692
rect 433794 161465 434414 182898
rect 437514 403174 438134 420068
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 161465 438134 186618
rect 441234 406894 441854 420423
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 444238 321061 444298 700435
rect 444954 698614 445574 707162
rect 448674 708678 449294 711590
rect 448674 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 449294 708678
rect 448674 708358 449294 708442
rect 448674 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 449294 708358
rect 447731 700364 447797 700365
rect 447731 700300 447732 700364
rect 447796 700300 447797 700364
rect 447731 700299 447797 700300
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 446259 683908 446325 683909
rect 446259 683844 446260 683908
rect 446324 683844 446325 683908
rect 446259 683843 446325 683844
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444235 321060 444301 321061
rect 444235 320996 444236 321060
rect 444300 320996 444301 321060
rect 444235 320995 444301 320996
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 161465 441854 190338
rect 444954 302614 445574 338058
rect 446262 319837 446322 683843
rect 446443 683772 446509 683773
rect 446443 683708 446444 683772
rect 446508 683708 446509 683772
rect 446443 683707 446509 683708
rect 446259 319836 446325 319837
rect 446259 319772 446260 319836
rect 446324 319772 446325 319836
rect 446259 319771 446325 319772
rect 446446 319565 446506 683707
rect 447734 321333 447794 700299
rect 447915 682820 447981 682821
rect 447915 682756 447916 682820
rect 447980 682756 447981 682820
rect 447915 682755 447981 682756
rect 447731 321332 447797 321333
rect 447731 321268 447732 321332
rect 447796 321268 447797 321332
rect 447731 321267 447797 321268
rect 447918 320109 447978 682755
rect 448674 666334 449294 708122
rect 452394 709638 453014 711590
rect 452394 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 453014 709638
rect 452394 709318 453014 709402
rect 452394 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 453014 709318
rect 450491 700636 450557 700637
rect 450491 700572 450492 700636
rect 450556 700572 450557 700636
rect 450491 700571 450557 700572
rect 448674 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 449294 666334
rect 448674 666014 449294 666098
rect 448674 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 449294 666014
rect 448674 630334 449294 665778
rect 448674 630098 448706 630334
rect 448942 630098 449026 630334
rect 449262 630098 449294 630334
rect 448674 630014 449294 630098
rect 448674 629778 448706 630014
rect 448942 629778 449026 630014
rect 449262 629778 449294 630014
rect 448674 594334 449294 629778
rect 448674 594098 448706 594334
rect 448942 594098 449026 594334
rect 449262 594098 449294 594334
rect 448674 594014 449294 594098
rect 448674 593778 448706 594014
rect 448942 593778 449026 594014
rect 449262 593778 449294 594014
rect 448674 558334 449294 593778
rect 448674 558098 448706 558334
rect 448942 558098 449026 558334
rect 449262 558098 449294 558334
rect 448674 558014 449294 558098
rect 448674 557778 448706 558014
rect 448942 557778 449026 558014
rect 449262 557778 449294 558014
rect 448674 522334 449294 557778
rect 448674 522098 448706 522334
rect 448942 522098 449026 522334
rect 449262 522098 449294 522334
rect 448674 522014 449294 522098
rect 448674 521778 448706 522014
rect 448942 521778 449026 522014
rect 449262 521778 449294 522014
rect 448674 486334 449294 521778
rect 448674 486098 448706 486334
rect 448942 486098 449026 486334
rect 449262 486098 449294 486334
rect 448674 486014 449294 486098
rect 448674 485778 448706 486014
rect 448942 485778 449026 486014
rect 449262 485778 449294 486014
rect 448674 450334 449294 485778
rect 448674 450098 448706 450334
rect 448942 450098 449026 450334
rect 449262 450098 449294 450334
rect 448674 450014 449294 450098
rect 448674 449778 448706 450014
rect 448942 449778 449026 450014
rect 449262 449778 449294 450014
rect 448674 414334 449294 449778
rect 448674 414098 448706 414334
rect 448942 414098 449026 414334
rect 449262 414098 449294 414334
rect 448674 414014 449294 414098
rect 448674 413778 448706 414014
rect 448942 413778 449026 414014
rect 449262 413778 449294 414014
rect 448674 378334 449294 413778
rect 448674 378098 448706 378334
rect 448942 378098 449026 378334
rect 449262 378098 449294 378334
rect 448674 378014 449294 378098
rect 448674 377778 448706 378014
rect 448942 377778 449026 378014
rect 449262 377778 449294 378014
rect 448674 342334 449294 377778
rect 448674 342098 448706 342334
rect 448942 342098 449026 342334
rect 449262 342098 449294 342334
rect 448674 342014 449294 342098
rect 448674 341778 448706 342014
rect 448942 341778 449026 342014
rect 449262 341778 449294 342014
rect 447915 320108 447981 320109
rect 447915 320044 447916 320108
rect 447980 320044 447981 320108
rect 447915 320043 447981 320044
rect 446443 319564 446509 319565
rect 446443 319500 446444 319564
rect 446508 319500 446509 319564
rect 446443 319499 446509 319500
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 161465 445574 194058
rect 448674 306334 449294 341778
rect 450494 320925 450554 700571
rect 450675 684044 450741 684045
rect 450675 683980 450676 684044
rect 450740 683980 450741 684044
rect 450675 683979 450741 683980
rect 450491 320924 450557 320925
rect 450491 320860 450492 320924
rect 450556 320860 450557 320924
rect 450491 320859 450557 320860
rect 450678 319973 450738 683979
rect 452394 670054 453014 709082
rect 452394 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 453014 670054
rect 452394 669734 453014 669818
rect 452394 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 453014 669734
rect 452394 634054 453014 669498
rect 452394 633818 452426 634054
rect 452662 633818 452746 634054
rect 452982 633818 453014 634054
rect 452394 633734 453014 633818
rect 452394 633498 452426 633734
rect 452662 633498 452746 633734
rect 452982 633498 453014 633734
rect 452394 598054 453014 633498
rect 452394 597818 452426 598054
rect 452662 597818 452746 598054
rect 452982 597818 453014 598054
rect 452394 597734 453014 597818
rect 452394 597498 452426 597734
rect 452662 597498 452746 597734
rect 452982 597498 453014 597734
rect 452394 562054 453014 597498
rect 452394 561818 452426 562054
rect 452662 561818 452746 562054
rect 452982 561818 453014 562054
rect 452394 561734 453014 561818
rect 452394 561498 452426 561734
rect 452662 561498 452746 561734
rect 452982 561498 453014 561734
rect 452394 526054 453014 561498
rect 452394 525818 452426 526054
rect 452662 525818 452746 526054
rect 452982 525818 453014 526054
rect 452394 525734 453014 525818
rect 452394 525498 452426 525734
rect 452662 525498 452746 525734
rect 452982 525498 453014 525734
rect 452394 517884 453014 525498
rect 456114 710598 456734 711590
rect 456114 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 456734 710598
rect 456114 710278 456734 710362
rect 456114 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 456734 710278
rect 456114 673774 456734 710042
rect 456114 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 456734 673774
rect 456114 673454 456734 673538
rect 456114 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 456734 673454
rect 456114 637774 456734 673218
rect 459834 711558 460454 711590
rect 459834 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 460454 711558
rect 459834 711238 460454 711322
rect 459834 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 460454 711238
rect 459834 677494 460454 711002
rect 459834 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 460454 677494
rect 459834 677174 460454 677258
rect 459834 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 460454 677174
rect 459834 668801 460454 676938
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 668801 470414 686898
rect 473514 705798 474134 711590
rect 473514 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 474134 705798
rect 473514 705478 474134 705562
rect 473514 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 474134 705478
rect 473514 691174 474134 705242
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 668801 474134 690618
rect 477234 706758 477854 711590
rect 477234 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 477854 706758
rect 477234 706438 477854 706522
rect 477234 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 477854 706438
rect 477234 694894 477854 706202
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 668801 477854 694338
rect 480954 707718 481574 711590
rect 480954 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 481574 707718
rect 480954 707398 481574 707482
rect 480954 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 481574 707398
rect 480954 698614 481574 707162
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 668801 481574 698058
rect 488394 709638 489014 711590
rect 488394 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 489014 709638
rect 488394 709318 489014 709402
rect 488394 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 489014 709318
rect 488394 670054 489014 709082
rect 488394 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 489014 670054
rect 488394 669734 489014 669818
rect 488394 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 489014 669734
rect 488394 668801 489014 669498
rect 492114 710598 492734 711590
rect 492114 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 492734 710598
rect 492114 710278 492734 710362
rect 492114 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 492734 710278
rect 492114 673774 492734 710042
rect 492114 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 492734 673774
rect 492114 673454 492734 673538
rect 492114 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 492734 673454
rect 492114 668801 492734 673218
rect 495834 711558 496454 711590
rect 495834 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 496454 711558
rect 495834 711238 496454 711322
rect 495834 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 496454 711238
rect 495834 677494 496454 711002
rect 495834 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 496454 677494
rect 495834 677174 496454 677258
rect 495834 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 496454 677174
rect 495834 668801 496454 676938
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 668801 506414 686898
rect 509514 705798 510134 711590
rect 509514 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 510134 705798
rect 509514 705478 510134 705562
rect 509514 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 510134 705478
rect 509514 691174 510134 705242
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 668801 510134 690618
rect 513234 706758 513854 711590
rect 513234 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 513854 706758
rect 513234 706438 513854 706522
rect 513234 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 513854 706438
rect 513234 694894 513854 706202
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 668801 513854 694338
rect 516954 707718 517574 711590
rect 516954 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 517574 707718
rect 516954 707398 517574 707482
rect 516954 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 517574 707398
rect 516954 698614 517574 707162
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 668801 517574 698058
rect 520674 708678 521294 711590
rect 520674 708442 520706 708678
rect 520942 708442 521026 708678
rect 521262 708442 521294 708678
rect 520674 708358 521294 708442
rect 520674 708122 520706 708358
rect 520942 708122 521026 708358
rect 521262 708122 521294 708358
rect 520674 666334 521294 708122
rect 520674 666098 520706 666334
rect 520942 666098 521026 666334
rect 521262 666098 521294 666334
rect 520674 666014 521294 666098
rect 520674 665778 520706 666014
rect 520942 665778 521026 666014
rect 521262 665778 521294 666014
rect 458035 665276 458101 665277
rect 458035 665212 458036 665276
rect 458100 665212 458101 665276
rect 458035 665211 458101 665212
rect 457851 662556 457917 662557
rect 457851 662492 457852 662556
rect 457916 662492 457917 662556
rect 457851 662491 457917 662492
rect 456114 637538 456146 637774
rect 456382 637538 456466 637774
rect 456702 637538 456734 637774
rect 456114 637454 456734 637538
rect 456114 637218 456146 637454
rect 456382 637218 456466 637454
rect 456702 637218 456734 637454
rect 456114 601774 456734 637218
rect 456114 601538 456146 601774
rect 456382 601538 456466 601774
rect 456702 601538 456734 601774
rect 456114 601454 456734 601538
rect 456114 601218 456146 601454
rect 456382 601218 456466 601454
rect 456702 601218 456734 601454
rect 456114 565774 456734 601218
rect 456114 565538 456146 565774
rect 456382 565538 456466 565774
rect 456702 565538 456734 565774
rect 456114 565454 456734 565538
rect 456114 565218 456146 565454
rect 456382 565218 456466 565454
rect 456702 565218 456734 565454
rect 456114 529774 456734 565218
rect 456114 529538 456146 529774
rect 456382 529538 456466 529774
rect 456702 529538 456734 529774
rect 456114 529454 456734 529538
rect 456114 529218 456146 529454
rect 456382 529218 456466 529454
rect 456702 529218 456734 529454
rect 456114 517884 456734 529218
rect 457854 521117 457914 662491
rect 458038 522341 458098 665211
rect 479568 655174 479888 655206
rect 479568 654938 479610 655174
rect 479846 654938 479888 655174
rect 479568 654854 479888 654938
rect 479568 654618 479610 654854
rect 479846 654618 479888 654854
rect 479568 654586 479888 654618
rect 510288 655174 510608 655206
rect 510288 654938 510330 655174
rect 510566 654938 510608 655174
rect 510288 654854 510608 654938
rect 510288 654618 510330 654854
rect 510566 654618 510608 654854
rect 510288 654586 510608 654618
rect 464208 651454 464528 651486
rect 464208 651218 464250 651454
rect 464486 651218 464528 651454
rect 464208 651134 464528 651218
rect 464208 650898 464250 651134
rect 464486 650898 464528 651134
rect 464208 650866 464528 650898
rect 494928 651454 495248 651486
rect 494928 651218 494970 651454
rect 495206 651218 495248 651454
rect 494928 651134 495248 651218
rect 494928 650898 494970 651134
rect 495206 650898 495248 651134
rect 494928 650866 495248 650898
rect 459139 630732 459205 630733
rect 459139 630668 459140 630732
rect 459204 630668 459205 630732
rect 459139 630667 459205 630668
rect 458035 522340 458101 522341
rect 458035 522276 458036 522340
rect 458100 522276 458101 522340
rect 458035 522275 458101 522276
rect 457851 521116 457917 521117
rect 457851 521052 457852 521116
rect 457916 521052 457917 521116
rect 457851 521051 457917 521052
rect 453382 511174 453702 511206
rect 453382 510938 453424 511174
rect 453660 510938 453702 511174
rect 453382 510854 453702 510938
rect 453382 510618 453424 510854
rect 453660 510618 453702 510854
rect 453382 510586 453702 510618
rect 455820 511174 456140 511206
rect 455820 510938 455862 511174
rect 456098 510938 456140 511174
rect 455820 510854 456140 510938
rect 455820 510618 455862 510854
rect 456098 510618 456140 510854
rect 455820 510586 456140 510618
rect 458258 511174 458578 511206
rect 458258 510938 458300 511174
rect 458536 510938 458578 511174
rect 458258 510854 458578 510938
rect 458258 510618 458300 510854
rect 458536 510618 458578 510854
rect 458258 510586 458578 510618
rect 452163 507454 452483 507486
rect 452163 507218 452205 507454
rect 452441 507218 452483 507454
rect 452163 507134 452483 507218
rect 452163 506898 452205 507134
rect 452441 506898 452483 507134
rect 452163 506866 452483 506898
rect 454601 507454 454921 507486
rect 454601 507218 454643 507454
rect 454879 507218 454921 507454
rect 454601 507134 454921 507218
rect 454601 506898 454643 507134
rect 454879 506898 454921 507134
rect 454601 506866 454921 506898
rect 457039 507454 457359 507486
rect 457039 507218 457081 507454
rect 457317 507218 457359 507454
rect 457039 507134 457359 507218
rect 457039 506898 457081 507134
rect 457317 506898 457359 507134
rect 457039 506866 457359 506898
rect 452394 490054 453014 500068
rect 452394 489818 452426 490054
rect 452662 489818 452746 490054
rect 452982 489818 453014 490054
rect 452394 489734 453014 489818
rect 452394 489498 452426 489734
rect 452662 489498 452746 489734
rect 452982 489498 453014 489734
rect 452394 454054 453014 489498
rect 452394 453818 452426 454054
rect 452662 453818 452746 454054
rect 452982 453818 453014 454054
rect 452394 453734 453014 453818
rect 452394 453498 452426 453734
rect 452662 453498 452746 453734
rect 452982 453498 453014 453734
rect 452394 418054 453014 453498
rect 452394 417818 452426 418054
rect 452662 417818 452746 418054
rect 452982 417818 453014 418054
rect 452394 417734 453014 417818
rect 452394 417498 452426 417734
rect 452662 417498 452746 417734
rect 452982 417498 453014 417734
rect 452394 382054 453014 417498
rect 452394 381818 452426 382054
rect 452662 381818 452746 382054
rect 452982 381818 453014 382054
rect 452394 381734 453014 381818
rect 452394 381498 452426 381734
rect 452662 381498 452746 381734
rect 452982 381498 453014 381734
rect 452394 346054 453014 381498
rect 456114 493774 456734 500068
rect 456114 493538 456146 493774
rect 456382 493538 456466 493774
rect 456702 493538 456734 493774
rect 456114 493454 456734 493538
rect 456114 493218 456146 493454
rect 456382 493218 456466 493454
rect 456702 493218 456734 493454
rect 456114 457774 456734 493218
rect 456114 457538 456146 457774
rect 456382 457538 456466 457774
rect 456702 457538 456734 457774
rect 456114 457454 456734 457538
rect 456114 457218 456146 457454
rect 456382 457218 456466 457454
rect 456702 457218 456734 457454
rect 456114 421774 456734 457218
rect 456114 421538 456146 421774
rect 456382 421538 456466 421774
rect 456702 421538 456734 421774
rect 456114 421454 456734 421538
rect 456114 421218 456146 421454
rect 456382 421218 456466 421454
rect 456702 421218 456734 421454
rect 456114 385774 456734 421218
rect 459142 391237 459202 630667
rect 520674 630334 521294 665778
rect 520674 630098 520706 630334
rect 520942 630098 521026 630334
rect 521262 630098 521294 630334
rect 520674 630014 521294 630098
rect 520674 629778 520706 630014
rect 520942 629778 521026 630014
rect 521262 629778 521294 630014
rect 479568 619174 479888 619206
rect 479568 618938 479610 619174
rect 479846 618938 479888 619174
rect 479568 618854 479888 618938
rect 479568 618618 479610 618854
rect 479846 618618 479888 618854
rect 479568 618586 479888 618618
rect 510288 619174 510608 619206
rect 510288 618938 510330 619174
rect 510566 618938 510608 619174
rect 510288 618854 510608 618938
rect 510288 618618 510330 618854
rect 510566 618618 510608 618854
rect 510288 618586 510608 618618
rect 464208 615454 464528 615486
rect 464208 615218 464250 615454
rect 464486 615218 464528 615454
rect 464208 615134 464528 615218
rect 464208 614898 464250 615134
rect 464486 614898 464528 615134
rect 464208 614866 464528 614898
rect 494928 615454 495248 615486
rect 494928 615218 494970 615454
rect 495206 615218 495248 615454
rect 494928 615134 495248 615218
rect 494928 614898 494970 615134
rect 495206 614898 495248 615134
rect 494928 614866 495248 614898
rect 459834 569494 460454 600287
rect 459834 569258 459866 569494
rect 460102 569258 460186 569494
rect 460422 569258 460454 569494
rect 459834 569174 460454 569258
rect 459834 568938 459866 569174
rect 460102 568938 460186 569174
rect 460422 568938 460454 569174
rect 459834 533494 460454 568938
rect 459834 533258 459866 533494
rect 460102 533258 460186 533494
rect 460422 533258 460454 533494
rect 459834 533174 460454 533258
rect 459834 532938 459866 533174
rect 460102 532938 460186 533174
rect 460422 532938 460454 533174
rect 459834 517884 460454 532938
rect 469794 579454 470414 600287
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 460696 511174 461016 511206
rect 460696 510938 460738 511174
rect 460974 510938 461016 511174
rect 460696 510854 461016 510938
rect 460696 510618 460738 510854
rect 460974 510618 461016 510854
rect 460696 510586 461016 510618
rect 459477 507454 459797 507486
rect 459477 507218 459519 507454
rect 459755 507218 459797 507454
rect 459477 507134 459797 507218
rect 459477 506898 459519 507134
rect 459755 506898 459797 507134
rect 459477 506866 459797 506898
rect 469794 507454 470414 542898
rect 473514 583174 474134 600287
rect 474779 599588 474845 599589
rect 474779 599524 474780 599588
rect 474844 599524 474845 599588
rect 474779 599523 474845 599524
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 472019 519620 472085 519621
rect 472019 519556 472020 519620
rect 472084 519556 472085 519620
rect 472019 519555 472085 519556
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 459834 497494 460454 500068
rect 459834 497258 459866 497494
rect 460102 497258 460186 497494
rect 460422 497258 460454 497494
rect 459834 497174 460454 497258
rect 459834 496938 459866 497174
rect 460102 496938 460186 497174
rect 460422 496938 460454 497174
rect 459834 461494 460454 496938
rect 459834 461258 459866 461494
rect 460102 461258 460186 461494
rect 460422 461258 460454 461494
rect 459834 461174 460454 461258
rect 459834 460938 459866 461174
rect 460102 460938 460186 461174
rect 460422 460938 460454 461174
rect 459834 425494 460454 460938
rect 459834 425258 459866 425494
rect 460102 425258 460186 425494
rect 460422 425258 460454 425494
rect 459834 425174 460454 425258
rect 459834 424938 459866 425174
rect 460102 424938 460186 425174
rect 460422 424938 460454 425174
rect 459139 391236 459205 391237
rect 459139 391172 459140 391236
rect 459204 391172 459205 391236
rect 459139 391171 459205 391172
rect 456114 385538 456146 385774
rect 456382 385538 456466 385774
rect 456702 385538 456734 385774
rect 456114 385454 456734 385538
rect 456114 385218 456146 385454
rect 456382 385218 456466 385454
rect 456702 385218 456734 385454
rect 454208 363454 454528 363486
rect 454208 363218 454250 363454
rect 454486 363218 454528 363454
rect 454208 363134 454528 363218
rect 454208 362898 454250 363134
rect 454486 362898 454528 363134
rect 454208 362866 454528 362898
rect 452394 345818 452426 346054
rect 452662 345818 452746 346054
rect 452982 345818 453014 346054
rect 452394 345734 453014 345818
rect 452394 345498 452426 345734
rect 452662 345498 452746 345734
rect 452982 345498 453014 345734
rect 450675 319972 450741 319973
rect 450675 319908 450676 319972
rect 450740 319908 450741 319972
rect 450675 319907 450741 319908
rect 448674 306098 448706 306334
rect 448942 306098 449026 306334
rect 449262 306098 449294 306334
rect 448674 306014 449294 306098
rect 448674 305778 448706 306014
rect 448942 305778 449026 306014
rect 449262 305778 449294 306014
rect 448674 270334 449294 305778
rect 448674 270098 448706 270334
rect 448942 270098 449026 270334
rect 449262 270098 449294 270334
rect 448674 270014 449294 270098
rect 448674 269778 448706 270014
rect 448942 269778 449026 270014
rect 449262 269778 449294 270014
rect 448674 234334 449294 269778
rect 448674 234098 448706 234334
rect 448942 234098 449026 234334
rect 449262 234098 449294 234334
rect 448674 234014 449294 234098
rect 448674 233778 448706 234014
rect 448942 233778 449026 234014
rect 449262 233778 449294 234014
rect 448674 198334 449294 233778
rect 448674 198098 448706 198334
rect 448942 198098 449026 198334
rect 449262 198098 449294 198334
rect 448674 198014 449294 198098
rect 448674 197778 448706 198014
rect 448942 197778 449026 198014
rect 449262 197778 449294 198014
rect 448674 162334 449294 197778
rect 448674 162098 448706 162334
rect 448942 162098 449026 162334
rect 449262 162098 449294 162334
rect 448674 162014 449294 162098
rect 448674 161778 448706 162014
rect 448942 161778 449026 162014
rect 449262 161778 449294 162014
rect 448674 161465 449294 161778
rect 452394 310054 453014 345498
rect 456114 349774 456734 385218
rect 456114 349538 456146 349774
rect 456382 349538 456466 349774
rect 456702 349538 456734 349774
rect 456114 349454 456734 349538
rect 456114 349218 456146 349454
rect 456382 349218 456466 349454
rect 456702 349218 456734 349454
rect 454208 327454 454528 327486
rect 454208 327218 454250 327454
rect 454486 327218 454528 327454
rect 454208 327134 454528 327218
rect 454208 326898 454250 327134
rect 454486 326898 454528 327134
rect 454208 326866 454528 326898
rect 452394 309818 452426 310054
rect 452662 309818 452746 310054
rect 452982 309818 453014 310054
rect 452394 309734 453014 309818
rect 452394 309498 452426 309734
rect 452662 309498 452746 309734
rect 452982 309498 453014 309734
rect 452394 274054 453014 309498
rect 452394 273818 452426 274054
rect 452662 273818 452746 274054
rect 452982 273818 453014 274054
rect 452394 273734 453014 273818
rect 452394 273498 452426 273734
rect 452662 273498 452746 273734
rect 452982 273498 453014 273734
rect 452394 238054 453014 273498
rect 452394 237818 452426 238054
rect 452662 237818 452746 238054
rect 452982 237818 453014 238054
rect 452394 237734 453014 237818
rect 452394 237498 452426 237734
rect 452662 237498 452746 237734
rect 452982 237498 453014 237734
rect 452394 202054 453014 237498
rect 452394 201818 452426 202054
rect 452662 201818 452746 202054
rect 452982 201818 453014 202054
rect 452394 201734 453014 201818
rect 452394 201498 452426 201734
rect 452662 201498 452746 201734
rect 452982 201498 453014 201734
rect 452394 166054 453014 201498
rect 452394 165818 452426 166054
rect 452662 165818 452746 166054
rect 452982 165818 453014 166054
rect 452394 165734 453014 165818
rect 452394 165498 452426 165734
rect 452662 165498 452746 165734
rect 452982 165498 453014 165734
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 429568 151174 429888 151206
rect 429568 150938 429610 151174
rect 429846 150938 429888 151174
rect 429568 150854 429888 150938
rect 429568 150618 429610 150854
rect 429846 150618 429888 150854
rect 429568 150586 429888 150618
rect 414208 147454 414528 147486
rect 414208 147218 414250 147454
rect 414486 147218 414528 147454
rect 414208 147134 414528 147218
rect 414208 146898 414250 147134
rect 414486 146898 414528 147134
rect 414208 146866 414528 146898
rect 444928 147454 445248 147486
rect 444928 147218 444970 147454
rect 445206 147218 445248 147454
rect 444928 147134 445248 147218
rect 444928 146898 444970 147134
rect 445206 146898 445248 147134
rect 444928 146866 445248 146898
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 92137 409574 122058
rect 452394 130054 453014 165498
rect 452394 129818 452426 130054
rect 452662 129818 452746 130054
rect 452982 129818 453014 130054
rect 452394 129734 453014 129818
rect 452394 129498 452426 129734
rect 452662 129498 452746 129734
rect 452982 129498 453014 129734
rect 416394 94054 417014 120423
rect 416394 93818 416426 94054
rect 416662 93818 416746 94054
rect 416982 93818 417014 94054
rect 416394 93734 417014 93818
rect 416394 93498 416426 93734
rect 416662 93498 416746 93734
rect 416982 93498 417014 93734
rect 416394 92137 417014 93498
rect 420114 97774 420734 120423
rect 420114 97538 420146 97774
rect 420382 97538 420466 97774
rect 420702 97538 420734 97774
rect 420114 97454 420734 97538
rect 420114 97218 420146 97454
rect 420382 97218 420466 97454
rect 420702 97218 420734 97454
rect 420114 92137 420734 97218
rect 423834 101494 424454 120423
rect 423834 101258 423866 101494
rect 424102 101258 424186 101494
rect 424422 101258 424454 101494
rect 423834 101174 424454 101258
rect 423834 100938 423866 101174
rect 424102 100938 424186 101174
rect 424422 100938 424454 101174
rect 423834 92137 424454 100938
rect 452394 94054 453014 129498
rect 452394 93818 452426 94054
rect 452662 93818 452746 94054
rect 452982 93818 453014 94054
rect 452394 93734 453014 93818
rect 452394 93498 452426 93734
rect 452662 93498 452746 93734
rect 452982 93498 453014 93734
rect 452394 92137 453014 93498
rect 456114 313774 456734 349218
rect 456114 313538 456146 313774
rect 456382 313538 456466 313774
rect 456702 313538 456734 313774
rect 456114 313454 456734 313538
rect 456114 313218 456146 313454
rect 456382 313218 456466 313454
rect 456702 313218 456734 313454
rect 456114 277774 456734 313218
rect 456114 277538 456146 277774
rect 456382 277538 456466 277774
rect 456702 277538 456734 277774
rect 456114 277454 456734 277538
rect 456114 277218 456146 277454
rect 456382 277218 456466 277454
rect 456702 277218 456734 277454
rect 456114 241774 456734 277218
rect 456114 241538 456146 241774
rect 456382 241538 456466 241774
rect 456702 241538 456734 241774
rect 456114 241454 456734 241538
rect 456114 241218 456146 241454
rect 456382 241218 456466 241454
rect 456702 241218 456734 241454
rect 456114 205774 456734 241218
rect 456114 205538 456146 205774
rect 456382 205538 456466 205774
rect 456702 205538 456734 205774
rect 456114 205454 456734 205538
rect 456114 205218 456146 205454
rect 456382 205218 456466 205454
rect 456702 205218 456734 205454
rect 456114 169774 456734 205218
rect 456114 169538 456146 169774
rect 456382 169538 456466 169774
rect 456702 169538 456734 169774
rect 456114 169454 456734 169538
rect 456114 169218 456146 169454
rect 456382 169218 456466 169454
rect 456702 169218 456734 169454
rect 456114 133774 456734 169218
rect 456114 133538 456146 133774
rect 456382 133538 456466 133774
rect 456702 133538 456734 133774
rect 456114 133454 456734 133538
rect 456114 133218 456146 133454
rect 456382 133218 456466 133454
rect 456702 133218 456734 133454
rect 456114 97774 456734 133218
rect 456114 97538 456146 97774
rect 456382 97538 456466 97774
rect 456702 97538 456734 97774
rect 456114 97454 456734 97538
rect 456114 97218 456146 97454
rect 456382 97218 456466 97454
rect 456702 97218 456734 97454
rect 456114 92137 456734 97218
rect 459834 389494 460454 424938
rect 459834 389258 459866 389494
rect 460102 389258 460186 389494
rect 460422 389258 460454 389494
rect 459834 389174 460454 389258
rect 459834 388938 459866 389174
rect 460102 388938 460186 389174
rect 460422 388938 460454 389174
rect 459834 353494 460454 388938
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 385580 470414 398898
rect 472022 389061 472082 519555
rect 473514 511174 474134 546618
rect 474411 520980 474477 520981
rect 474411 520916 474412 520980
rect 474476 520916 474477 520980
rect 474411 520915 474477 520916
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 453692 474134 474618
rect 473416 435454 473736 435486
rect 473416 435218 473458 435454
rect 473694 435218 473736 435454
rect 473416 435134 473736 435218
rect 473416 434898 473458 435134
rect 473694 434898 473736 435134
rect 473416 434866 473736 434898
rect 474414 389061 474474 520915
rect 474595 519484 474661 519485
rect 474595 519420 474596 519484
rect 474660 519420 474661 519484
rect 474595 519419 474661 519420
rect 472019 389060 472085 389061
rect 472019 388996 472020 389060
rect 472084 388996 472085 389060
rect 472019 388995 472085 388996
rect 474411 389060 474477 389061
rect 474411 388996 474412 389060
rect 474476 388996 474477 389060
rect 474411 388995 474477 388996
rect 474598 388925 474658 519419
rect 474782 389061 474842 599523
rect 476435 598228 476501 598229
rect 476435 598164 476436 598228
rect 476500 598164 476501 598228
rect 476435 598163 476501 598164
rect 475888 439174 476208 439206
rect 475888 438938 475930 439174
rect 476166 438938 476208 439174
rect 475888 438854 476208 438938
rect 475888 438618 475930 438854
rect 476166 438618 476208 438854
rect 475888 438586 476208 438618
rect 476438 389061 476498 598163
rect 477234 586894 477854 600287
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 480954 590614 481574 600287
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 478827 543012 478893 543013
rect 478827 542948 478828 543012
rect 478892 542948 478893 543012
rect 478827 542947 478893 542948
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 478361 435454 478681 435486
rect 478361 435218 478403 435454
rect 478639 435218 478681 435454
rect 478361 435134 478681 435218
rect 478361 434898 478403 435134
rect 478639 434898 478681 435134
rect 478361 434866 478681 434898
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 474779 389060 474845 389061
rect 474779 388996 474780 389060
rect 474844 388996 474845 389060
rect 474779 388995 474845 388996
rect 476435 389060 476501 389061
rect 476435 388996 476436 389060
rect 476500 388996 476501 389060
rect 476435 388995 476501 388996
rect 474595 388924 474661 388925
rect 474595 388860 474596 388924
rect 474660 388860 474661 388924
rect 474595 388859 474661 388860
rect 477234 385225 477854 406338
rect 478830 389061 478890 542947
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 484674 594334 485294 600287
rect 484674 594098 484706 594334
rect 484942 594098 485026 594334
rect 485262 594098 485294 594334
rect 484674 594014 485294 594098
rect 484674 593778 484706 594014
rect 484942 593778 485026 594014
rect 485262 593778 485294 594014
rect 484674 558334 485294 593778
rect 484674 558098 484706 558334
rect 484942 558098 485026 558334
rect 485262 558098 485294 558334
rect 484674 558014 485294 558098
rect 484674 557778 484706 558014
rect 484942 557778 485026 558014
rect 485262 557778 485294 558014
rect 484674 522334 485294 557778
rect 484674 522098 484706 522334
rect 484942 522098 485026 522334
rect 485262 522098 485294 522334
rect 484674 522014 485294 522098
rect 484674 521778 484706 522014
rect 484942 521778 485026 522014
rect 485262 521778 485294 522014
rect 484674 517884 485294 521778
rect 488394 598054 489014 600287
rect 488394 597818 488426 598054
rect 488662 597818 488746 598054
rect 488982 597818 489014 598054
rect 488394 597734 489014 597818
rect 488394 597498 488426 597734
rect 488662 597498 488746 597734
rect 488982 597498 489014 597734
rect 488394 562054 489014 597498
rect 488394 561818 488426 562054
rect 488662 561818 488746 562054
rect 488982 561818 489014 562054
rect 488394 561734 489014 561818
rect 488394 561498 488426 561734
rect 488662 561498 488746 561734
rect 488982 561498 489014 561734
rect 488394 526054 489014 561498
rect 488394 525818 488426 526054
rect 488662 525818 488746 526054
rect 488982 525818 489014 526054
rect 488394 525734 489014 525818
rect 488394 525498 488426 525734
rect 488662 525498 488746 525734
rect 488982 525498 489014 525734
rect 488394 517884 489014 525498
rect 492114 565774 492734 600287
rect 492114 565538 492146 565774
rect 492382 565538 492466 565774
rect 492702 565538 492734 565774
rect 492114 565454 492734 565538
rect 492114 565218 492146 565454
rect 492382 565218 492466 565454
rect 492702 565218 492734 565454
rect 492114 529774 492734 565218
rect 492114 529538 492146 529774
rect 492382 529538 492466 529774
rect 492702 529538 492734 529774
rect 492114 529454 492734 529538
rect 492114 529218 492146 529454
rect 492382 529218 492466 529454
rect 492702 529218 492734 529454
rect 483382 511174 483702 511206
rect 483382 510938 483424 511174
rect 483660 510938 483702 511174
rect 483382 510854 483702 510938
rect 483382 510618 483424 510854
rect 483660 510618 483702 510854
rect 483382 510586 483702 510618
rect 485820 511174 486140 511206
rect 485820 510938 485862 511174
rect 486098 510938 486140 511174
rect 485820 510854 486140 510938
rect 485820 510618 485862 510854
rect 486098 510618 486140 510854
rect 485820 510586 486140 510618
rect 488258 511174 488578 511206
rect 488258 510938 488300 511174
rect 488536 510938 488578 511174
rect 488258 510854 488578 510938
rect 488258 510618 488300 510854
rect 488536 510618 488578 510854
rect 488258 510586 488578 510618
rect 490696 511174 491016 511206
rect 490696 510938 490738 511174
rect 490974 510938 491016 511174
rect 490696 510854 491016 510938
rect 490696 510618 490738 510854
rect 490974 510618 491016 510854
rect 490696 510586 491016 510618
rect 482163 507454 482483 507486
rect 482163 507218 482205 507454
rect 482441 507218 482483 507454
rect 482163 507134 482483 507218
rect 482163 506898 482205 507134
rect 482441 506898 482483 507134
rect 482163 506866 482483 506898
rect 484601 507454 484921 507486
rect 484601 507218 484643 507454
rect 484879 507218 484921 507454
rect 484601 507134 484921 507218
rect 484601 506898 484643 507134
rect 484879 506898 484921 507134
rect 484601 506866 484921 506898
rect 487039 507454 487359 507486
rect 487039 507218 487081 507454
rect 487317 507218 487359 507454
rect 487039 507134 487359 507218
rect 487039 506898 487081 507134
rect 487317 506898 487359 507134
rect 487039 506866 487359 506898
rect 489477 507454 489797 507486
rect 489477 507218 489519 507454
rect 489755 507218 489797 507454
rect 489477 507134 489797 507218
rect 489477 506898 489519 507134
rect 489755 506898 489797 507134
rect 489477 506866 489797 506898
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 453692 481574 482058
rect 484674 486334 485294 500068
rect 484674 486098 484706 486334
rect 484942 486098 485026 486334
rect 485262 486098 485294 486334
rect 484674 486014 485294 486098
rect 484674 485778 484706 486014
rect 484942 485778 485026 486014
rect 485262 485778 485294 486014
rect 484674 450334 485294 485778
rect 488394 490054 489014 500068
rect 488394 489818 488426 490054
rect 488662 489818 488746 490054
rect 488982 489818 489014 490054
rect 488394 489734 489014 489818
rect 488394 489498 488426 489734
rect 488662 489498 488746 489734
rect 488982 489498 489014 489734
rect 488394 454007 489014 489498
rect 487107 453932 487173 453933
rect 487107 453868 487108 453932
rect 487172 453868 487173 453932
rect 487107 453867 487173 453868
rect 484674 450098 484706 450334
rect 484942 450098 485026 450334
rect 485262 450098 485294 450334
rect 484674 450014 485294 450098
rect 484674 449778 484706 450014
rect 484942 449778 485026 450014
rect 485262 449778 485294 450014
rect 480833 439174 481153 439206
rect 480833 438938 480875 439174
rect 481111 438938 481153 439174
rect 480833 438854 481153 438938
rect 480833 438618 480875 438854
rect 481111 438618 481153 438854
rect 480833 438586 481153 438618
rect 483306 435454 483626 435486
rect 483306 435218 483348 435454
rect 483584 435218 483626 435454
rect 483306 435134 483626 435218
rect 483306 434898 483348 435134
rect 483584 434898 483626 435134
rect 483306 434866 483626 434898
rect 484674 414334 485294 449778
rect 485778 439174 486098 439206
rect 485778 438938 485820 439174
rect 486056 438938 486098 439174
rect 485778 438854 486098 438938
rect 485778 438618 485820 438854
rect 486056 438618 486098 438854
rect 485778 438586 486098 438618
rect 484674 414098 484706 414334
rect 484942 414098 485026 414334
rect 485262 414098 485294 414334
rect 484674 414014 485294 414098
rect 484674 413778 484706 414014
rect 484942 413778 485026 414014
rect 485262 413778 485294 414014
rect 478827 389060 478893 389061
rect 478827 388996 478828 389060
rect 478892 388996 478893 389060
rect 478827 388995 478893 388996
rect 484674 385580 485294 413778
rect 487110 385661 487170 453867
rect 488394 453771 488426 454007
rect 488662 453771 488746 454007
rect 488982 453771 489014 454007
rect 488394 453692 489014 453771
rect 492114 493774 492734 529218
rect 492114 493538 492146 493774
rect 492382 493538 492466 493774
rect 492702 493538 492734 493774
rect 492114 493454 492734 493538
rect 492114 493218 492146 493454
rect 492382 493218 492466 493454
rect 492702 493218 492734 493454
rect 492114 457774 492734 493218
rect 492114 457538 492146 457774
rect 492382 457538 492466 457774
rect 492702 457538 492734 457774
rect 492114 457454 492734 457538
rect 492114 457218 492146 457454
rect 492382 457218 492466 457454
rect 492702 457218 492734 457454
rect 490723 439174 491043 439206
rect 490723 438938 490765 439174
rect 491001 438938 491043 439174
rect 490723 438854 491043 438938
rect 490723 438618 490765 438854
rect 491001 438618 491043 438854
rect 490723 438586 491043 438618
rect 488251 435454 488571 435486
rect 488251 435218 488293 435454
rect 488529 435218 488571 435454
rect 488251 435134 488571 435218
rect 488251 434898 488293 435134
rect 488529 434898 488571 435134
rect 488251 434866 488571 434898
rect 492114 421774 492734 457218
rect 492114 421538 492146 421774
rect 492382 421538 492466 421774
rect 492702 421538 492734 421774
rect 492114 421454 492734 421538
rect 492114 421218 492146 421454
rect 492382 421218 492466 421454
rect 492702 421218 492734 421454
rect 487107 385660 487173 385661
rect 487107 385596 487108 385660
rect 487172 385596 487173 385660
rect 487107 385595 487173 385596
rect 492114 385225 492734 421218
rect 495834 569494 496454 600287
rect 495834 569258 495866 569494
rect 496102 569258 496186 569494
rect 496422 569258 496454 569494
rect 495834 569174 496454 569258
rect 495834 568938 495866 569174
rect 496102 568938 496186 569174
rect 496422 568938 496454 569174
rect 495834 533494 496454 568938
rect 495834 533258 495866 533494
rect 496102 533258 496186 533494
rect 496422 533258 496454 533494
rect 495834 533174 496454 533258
rect 495834 532938 495866 533174
rect 496102 532938 496186 533174
rect 496422 532938 496454 533174
rect 495834 497494 496454 532938
rect 495834 497258 495866 497494
rect 496102 497258 496186 497494
rect 496422 497258 496454 497494
rect 495834 497174 496454 497258
rect 495834 496938 495866 497174
rect 496102 496938 496186 497174
rect 496422 496938 496454 497174
rect 495834 461494 496454 496938
rect 495834 461258 495866 461494
rect 496102 461258 496186 461494
rect 496422 461258 496454 461494
rect 495834 461174 496454 461258
rect 495834 460938 495866 461174
rect 496102 460938 496186 461174
rect 496422 460938 496454 461174
rect 495834 425494 496454 460938
rect 495834 425258 495866 425494
rect 496102 425258 496186 425494
rect 496422 425258 496454 425494
rect 495834 425174 496454 425258
rect 495834 424938 495866 425174
rect 496102 424938 496186 425174
rect 496422 424938 496454 425174
rect 495834 389494 496454 424938
rect 495834 389258 495866 389494
rect 496102 389258 496186 389494
rect 496422 389258 496454 389494
rect 495834 389174 496454 389258
rect 495834 388938 495866 389174
rect 496102 388938 496186 389174
rect 496422 388938 496454 389174
rect 495834 385225 496454 388938
rect 505794 579454 506414 600287
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 469568 367174 469888 367206
rect 469568 366938 469610 367174
rect 469846 366938 469888 367174
rect 469568 366854 469888 366938
rect 469568 366618 469610 366854
rect 469846 366618 469888 366854
rect 469568 366586 469888 366618
rect 500288 367174 500608 367206
rect 500288 366938 500330 367174
rect 500566 366938 500608 367174
rect 500288 366854 500608 366938
rect 500288 366618 500330 366854
rect 500566 366618 500608 366854
rect 500288 366586 500608 366618
rect 484928 363454 485248 363486
rect 484928 363218 484970 363454
rect 485206 363218 485248 363454
rect 484928 363134 485248 363218
rect 484928 362898 484970 363134
rect 485206 362898 485248 363134
rect 484928 362866 485248 362898
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 459834 353258 459866 353494
rect 460102 353258 460186 353494
rect 460422 353258 460454 353494
rect 459834 353174 460454 353258
rect 459834 352938 459866 353174
rect 460102 352938 460186 353174
rect 460422 352938 460454 353174
rect 459834 317494 460454 352938
rect 469568 331174 469888 331206
rect 469568 330938 469610 331174
rect 469846 330938 469888 331174
rect 469568 330854 469888 330938
rect 469568 330618 469610 330854
rect 469846 330618 469888 330854
rect 469568 330586 469888 330618
rect 500288 331174 500608 331206
rect 500288 330938 500330 331174
rect 500566 330938 500608 331174
rect 500288 330854 500608 330938
rect 500288 330618 500330 330854
rect 500566 330618 500608 330854
rect 500288 330586 500608 330618
rect 484928 327454 485248 327486
rect 484928 327218 484970 327454
rect 485206 327218 485248 327454
rect 484928 327134 485248 327218
rect 484928 326898 484970 327134
rect 485206 326898 485248 327134
rect 484928 326866 485248 326898
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 459834 317258 459866 317494
rect 460102 317258 460186 317494
rect 460422 317258 460454 317494
rect 459834 317174 460454 317258
rect 459834 316938 459866 317174
rect 460102 316938 460186 317174
rect 460422 316938 460454 317174
rect 459834 281494 460454 316938
rect 459834 281258 459866 281494
rect 460102 281258 460186 281494
rect 460422 281258 460454 281494
rect 459834 281174 460454 281258
rect 459834 280938 459866 281174
rect 460102 280938 460186 281174
rect 460422 280938 460454 281174
rect 459834 245494 460454 280938
rect 477234 298894 477854 320655
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 259417 477854 262338
rect 480954 302614 481574 320655
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 259417 481574 266058
rect 484674 306334 485294 320655
rect 484674 306098 484706 306334
rect 484942 306098 485026 306334
rect 485262 306098 485294 306334
rect 484674 306014 485294 306098
rect 484674 305778 484706 306014
rect 484942 305778 485026 306014
rect 485262 305778 485294 306014
rect 484674 270334 485294 305778
rect 484674 270098 484706 270334
rect 484942 270098 485026 270334
rect 485262 270098 485294 270334
rect 484674 270014 485294 270098
rect 484674 269778 484706 270014
rect 484942 269778 485026 270014
rect 485262 269778 485294 270014
rect 484674 259417 485294 269778
rect 488394 310054 489014 320655
rect 488394 309818 488426 310054
rect 488662 309818 488746 310054
rect 488982 309818 489014 310054
rect 488394 309734 489014 309818
rect 488394 309498 488426 309734
rect 488662 309498 488746 309734
rect 488982 309498 489014 309734
rect 488394 274054 489014 309498
rect 488394 273818 488426 274054
rect 488662 273818 488746 274054
rect 488982 273818 489014 274054
rect 488394 273734 489014 273818
rect 488394 273498 488426 273734
rect 488662 273498 488746 273734
rect 488982 273498 489014 273734
rect 488394 259417 489014 273498
rect 492114 313774 492734 320655
rect 492114 313538 492146 313774
rect 492382 313538 492466 313774
rect 492702 313538 492734 313774
rect 492114 313454 492734 313538
rect 492114 313218 492146 313454
rect 492382 313218 492466 313454
rect 492702 313218 492734 313454
rect 492114 277774 492734 313218
rect 492114 277538 492146 277774
rect 492382 277538 492466 277774
rect 492702 277538 492734 277774
rect 492114 277454 492734 277538
rect 492114 277218 492146 277454
rect 492382 277218 492466 277454
rect 492702 277218 492734 277454
rect 492114 259417 492734 277218
rect 495834 317494 496454 320655
rect 495834 317258 495866 317494
rect 496102 317258 496186 317494
rect 496422 317258 496454 317494
rect 495834 317174 496454 317258
rect 495834 316938 495866 317174
rect 496102 316938 496186 317174
rect 496422 316938 496454 317174
rect 495834 281494 496454 316938
rect 495834 281258 495866 281494
rect 496102 281258 496186 281494
rect 496422 281258 496454 281494
rect 495834 281174 496454 281258
rect 495834 280938 495866 281174
rect 496102 280938 496186 281174
rect 496422 280938 496454 281174
rect 495834 259417 496454 280938
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 259417 506414 290898
rect 509514 583174 510134 600287
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 513234 586894 513854 600287
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 510659 342820 510725 342821
rect 510659 342756 510660 342820
rect 510724 342756 510725 342820
rect 510659 342755 510725 342756
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 510291 324868 510357 324869
rect 510291 324804 510292 324868
rect 510356 324804 510357 324868
rect 510291 324803 510357 324804
rect 510294 321877 510354 324803
rect 510475 323780 510541 323781
rect 510475 323716 510476 323780
rect 510540 323716 510541 323780
rect 510475 323715 510541 323716
rect 510291 321876 510357 321877
rect 510291 321812 510292 321876
rect 510356 321812 510357 321876
rect 510291 321811 510357 321812
rect 510478 306237 510538 323715
rect 510475 306236 510541 306237
rect 510475 306172 510476 306236
rect 510540 306172 510541 306236
rect 510475 306171 510541 306172
rect 510662 305829 510722 342755
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 510843 327588 510909 327589
rect 510843 327524 510844 327588
rect 510908 327524 510909 327588
rect 510843 327523 510909 327524
rect 510846 321333 510906 327523
rect 511211 326500 511277 326501
rect 511211 326436 511212 326500
rect 511276 326436 511277 326500
rect 511211 326435 511277 326436
rect 511027 325956 511093 325957
rect 511027 325892 511028 325956
rect 511092 325892 511093 325956
rect 511027 325891 511093 325892
rect 511030 321741 511090 325891
rect 511027 321740 511093 321741
rect 511027 321676 511028 321740
rect 511092 321676 511093 321740
rect 511027 321675 511093 321676
rect 510843 321332 510909 321333
rect 510843 321268 510844 321332
rect 510908 321268 510909 321332
rect 510843 321267 510909 321268
rect 511214 316050 511274 326435
rect 510846 315990 511274 316050
rect 510846 305965 510906 315990
rect 510843 305964 510909 305965
rect 510843 305900 510844 305964
rect 510908 305900 510909 305964
rect 510843 305899 510909 305900
rect 510659 305828 510725 305829
rect 510659 305764 510660 305828
rect 510724 305764 510725 305828
rect 510659 305763 510725 305764
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259417 510134 294618
rect 513234 298894 513854 334338
rect 516954 590614 517574 600287
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 514891 333028 514957 333029
rect 514891 332964 514892 333028
rect 514956 332964 514957 333028
rect 514891 332963 514957 332964
rect 514339 330852 514405 330853
rect 514339 330788 514340 330852
rect 514404 330788 514405 330852
rect 514339 330787 514405 330788
rect 514155 328132 514221 328133
rect 514155 328068 514156 328132
rect 514220 328068 514221 328132
rect 514155 328067 514221 328068
rect 514158 302973 514218 328067
rect 514342 320925 514402 330787
rect 514707 330308 514773 330309
rect 514707 330244 514708 330308
rect 514772 330244 514773 330308
rect 514707 330243 514773 330244
rect 514339 320924 514405 320925
rect 514339 320860 514340 320924
rect 514404 320860 514405 320924
rect 514339 320859 514405 320860
rect 514155 302972 514221 302973
rect 514155 302908 514156 302972
rect 514220 302908 514221 302972
rect 514155 302907 514221 302908
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 514710 291821 514770 330243
rect 514894 300117 514954 332963
rect 516954 302614 517574 338058
rect 520674 594334 521294 629778
rect 520674 594098 520706 594334
rect 520942 594098 521026 594334
rect 521262 594098 521294 594334
rect 520674 594014 521294 594098
rect 520674 593778 520706 594014
rect 520942 593778 521026 594014
rect 521262 593778 521294 594014
rect 520674 558334 521294 593778
rect 520674 558098 520706 558334
rect 520942 558098 521026 558334
rect 521262 558098 521294 558334
rect 520674 558014 521294 558098
rect 520674 557778 520706 558014
rect 520942 557778 521026 558014
rect 521262 557778 521294 558014
rect 520674 522334 521294 557778
rect 520674 522098 520706 522334
rect 520942 522098 521026 522334
rect 521262 522098 521294 522334
rect 520674 522014 521294 522098
rect 520674 521778 520706 522014
rect 520942 521778 521026 522014
rect 521262 521778 521294 522014
rect 520674 486334 521294 521778
rect 520674 486098 520706 486334
rect 520942 486098 521026 486334
rect 521262 486098 521294 486334
rect 520674 486014 521294 486098
rect 520674 485778 520706 486014
rect 520942 485778 521026 486014
rect 521262 485778 521294 486014
rect 520674 450334 521294 485778
rect 520674 450098 520706 450334
rect 520942 450098 521026 450334
rect 521262 450098 521294 450334
rect 520674 450014 521294 450098
rect 520674 449778 520706 450014
rect 520942 449778 521026 450014
rect 521262 449778 521294 450014
rect 520674 414334 521294 449778
rect 520674 414098 520706 414334
rect 520942 414098 521026 414334
rect 521262 414098 521294 414334
rect 520674 414014 521294 414098
rect 520674 413778 520706 414014
rect 520942 413778 521026 414014
rect 521262 413778 521294 414014
rect 520674 378334 521294 413778
rect 520674 378098 520706 378334
rect 520942 378098 521026 378334
rect 521262 378098 521294 378334
rect 520674 378014 521294 378098
rect 520674 377778 520706 378014
rect 520942 377778 521026 378014
rect 521262 377778 521294 378014
rect 520674 342334 521294 377778
rect 520674 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 521294 342334
rect 520674 342014 521294 342098
rect 520674 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 521294 342014
rect 517835 329220 517901 329221
rect 517835 329156 517836 329220
rect 517900 329156 517901 329220
rect 517835 329155 517901 329156
rect 517838 320789 517898 329155
rect 517835 320788 517901 320789
rect 517835 320724 517836 320788
rect 517900 320724 517901 320788
rect 517835 320723 517901 320724
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 514891 300116 514957 300117
rect 514891 300052 514892 300116
rect 514956 300052 514957 300116
rect 514891 300051 514957 300052
rect 514707 291820 514773 291821
rect 514707 291756 514708 291820
rect 514772 291756 514773 291820
rect 514707 291755 514773 291756
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 259417 513854 262338
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 259417 517574 266058
rect 520674 306334 521294 341778
rect 520674 306098 520706 306334
rect 520942 306098 521026 306334
rect 521262 306098 521294 306334
rect 520674 306014 521294 306098
rect 520674 305778 520706 306014
rect 520942 305778 521026 306014
rect 521262 305778 521294 306014
rect 520674 270334 521294 305778
rect 520674 270098 520706 270334
rect 520942 270098 521026 270334
rect 521262 270098 521294 270334
rect 520674 270014 521294 270098
rect 520674 269778 520706 270014
rect 520942 269778 521026 270014
rect 521262 269778 521294 270014
rect 520674 259417 521294 269778
rect 524394 709638 525014 711590
rect 524394 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 525014 709638
rect 524394 709318 525014 709402
rect 524394 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 525014 709318
rect 524394 670054 525014 709082
rect 528114 710598 528734 711590
rect 528114 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 528734 710598
rect 528114 710278 528734 710362
rect 528114 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 528734 710278
rect 526299 699820 526365 699821
rect 526299 699756 526300 699820
rect 526364 699756 526365 699820
rect 526299 699755 526365 699756
rect 524394 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 525014 670054
rect 524394 669734 525014 669818
rect 524394 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 525014 669734
rect 524394 634054 525014 669498
rect 525648 651454 525968 651486
rect 525648 651218 525690 651454
rect 525926 651218 525968 651454
rect 525648 651134 525968 651218
rect 525648 650898 525690 651134
rect 525926 650898 525968 651134
rect 525648 650866 525968 650898
rect 524394 633818 524426 634054
rect 524662 633818 524746 634054
rect 524982 633818 525014 634054
rect 524394 633734 525014 633818
rect 524394 633498 524426 633734
rect 524662 633498 524746 633734
rect 524982 633498 525014 633734
rect 524394 598054 525014 633498
rect 525648 615454 525968 615486
rect 525648 615218 525690 615454
rect 525926 615218 525968 615454
rect 525648 615134 525968 615218
rect 525648 614898 525690 615134
rect 525926 614898 525968 615134
rect 525648 614866 525968 614898
rect 524394 597818 524426 598054
rect 524662 597818 524746 598054
rect 524982 597818 525014 598054
rect 524394 597734 525014 597818
rect 524394 597498 524426 597734
rect 524662 597498 524746 597734
rect 524982 597498 525014 597734
rect 524394 562054 525014 597498
rect 524394 561818 524426 562054
rect 524662 561818 524746 562054
rect 524982 561818 525014 562054
rect 524394 561734 525014 561818
rect 524394 561498 524426 561734
rect 524662 561498 524746 561734
rect 524982 561498 525014 561734
rect 524394 526054 525014 561498
rect 524394 525818 524426 526054
rect 524662 525818 524746 526054
rect 524982 525818 525014 526054
rect 524394 525734 525014 525818
rect 524394 525498 524426 525734
rect 524662 525498 524746 525734
rect 524982 525498 525014 525734
rect 524394 490054 525014 525498
rect 524394 489818 524426 490054
rect 524662 489818 524746 490054
rect 524982 489818 525014 490054
rect 524394 489734 525014 489818
rect 524394 489498 524426 489734
rect 524662 489498 524746 489734
rect 524982 489498 525014 489734
rect 524394 454054 525014 489498
rect 524394 453818 524426 454054
rect 524662 453818 524746 454054
rect 524982 453818 525014 454054
rect 524394 453734 525014 453818
rect 524394 453498 524426 453734
rect 524662 453498 524746 453734
rect 524982 453498 525014 453734
rect 524394 418054 525014 453498
rect 525164 435454 525484 435486
rect 525164 435218 525206 435454
rect 525442 435218 525484 435454
rect 525164 435134 525484 435218
rect 525164 434898 525206 435134
rect 525442 434898 525484 435134
rect 525164 434866 525484 434898
rect 524394 417818 524426 418054
rect 524662 417818 524746 418054
rect 524982 417818 525014 418054
rect 524394 417734 525014 417818
rect 524394 417498 524426 417734
rect 524662 417498 524746 417734
rect 524982 417498 525014 417734
rect 524394 382054 525014 417498
rect 524394 381818 524426 382054
rect 524662 381818 524746 382054
rect 524982 381818 525014 382054
rect 524394 381734 525014 381818
rect 524394 381498 524426 381734
rect 524662 381498 524746 381734
rect 524982 381498 525014 381734
rect 524394 346054 525014 381498
rect 524394 345818 524426 346054
rect 524662 345818 524746 346054
rect 524982 345818 525014 346054
rect 524394 345734 525014 345818
rect 524394 345498 524426 345734
rect 524662 345498 524746 345734
rect 524982 345498 525014 345734
rect 524394 310054 525014 345498
rect 526302 320109 526362 699755
rect 528114 673774 528734 710042
rect 528114 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 528734 673774
rect 528114 673454 528734 673538
rect 528114 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 528734 673454
rect 528114 637774 528734 673218
rect 528114 637538 528146 637774
rect 528382 637538 528466 637774
rect 528702 637538 528734 637774
rect 528114 637454 528734 637538
rect 528114 637218 528146 637454
rect 528382 637218 528466 637454
rect 528702 637218 528734 637454
rect 528114 601774 528734 637218
rect 528114 601538 528146 601774
rect 528382 601538 528466 601774
rect 528702 601538 528734 601774
rect 528114 601454 528734 601538
rect 528114 601218 528146 601454
rect 528382 601218 528466 601454
rect 528702 601218 528734 601454
rect 528114 565774 528734 601218
rect 528114 565538 528146 565774
rect 528382 565538 528466 565774
rect 528702 565538 528734 565774
rect 528114 565454 528734 565538
rect 528114 565218 528146 565454
rect 528382 565218 528466 565454
rect 528702 565218 528734 565454
rect 528114 529774 528734 565218
rect 528114 529538 528146 529774
rect 528382 529538 528466 529774
rect 528702 529538 528734 529774
rect 528114 529454 528734 529538
rect 528114 529218 528146 529454
rect 528382 529218 528466 529454
rect 528702 529218 528734 529454
rect 528114 493774 528734 529218
rect 528114 493538 528146 493774
rect 528382 493538 528466 493774
rect 528702 493538 528734 493774
rect 528114 493454 528734 493538
rect 528114 493218 528146 493454
rect 528382 493218 528466 493454
rect 528702 493218 528734 493454
rect 528114 457774 528734 493218
rect 528114 457538 528146 457774
rect 528382 457538 528466 457774
rect 528702 457538 528734 457774
rect 528114 457454 528734 457538
rect 528114 457218 528146 457454
rect 528382 457218 528466 457454
rect 528702 457218 528734 457454
rect 528114 421774 528734 457218
rect 531834 711558 532454 711590
rect 531834 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 532454 711558
rect 531834 711238 532454 711322
rect 531834 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 532454 711238
rect 531834 677494 532454 711002
rect 531834 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 532454 677494
rect 531834 677174 532454 677258
rect 531834 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 532454 677174
rect 531834 641494 532454 676938
rect 531834 641258 531866 641494
rect 532102 641258 532186 641494
rect 532422 641258 532454 641494
rect 531834 641174 532454 641258
rect 531834 640938 531866 641174
rect 532102 640938 532186 641174
rect 532422 640938 532454 641174
rect 531834 605494 532454 640938
rect 531834 605258 531866 605494
rect 532102 605258 532186 605494
rect 532422 605258 532454 605494
rect 531834 605174 532454 605258
rect 531834 604938 531866 605174
rect 532102 604938 532186 605174
rect 532422 604938 532454 605174
rect 531834 569494 532454 604938
rect 531834 569258 531866 569494
rect 532102 569258 532186 569494
rect 532422 569258 532454 569494
rect 531834 569174 532454 569258
rect 531834 568938 531866 569174
rect 532102 568938 532186 569174
rect 532422 568938 532454 569174
rect 531834 533494 532454 568938
rect 531834 533258 531866 533494
rect 532102 533258 532186 533494
rect 532422 533258 532454 533494
rect 531834 533174 532454 533258
rect 531834 532938 531866 533174
rect 532102 532938 532186 533174
rect 532422 532938 532454 533174
rect 531834 497494 532454 532938
rect 531834 497258 531866 497494
rect 532102 497258 532186 497494
rect 532422 497258 532454 497494
rect 531834 497174 532454 497258
rect 531834 496938 531866 497174
rect 532102 496938 532186 497174
rect 532422 496938 532454 497174
rect 531834 461494 532454 496938
rect 531834 461258 531866 461494
rect 532102 461258 532186 461494
rect 532422 461258 532454 461494
rect 531834 461174 532454 461258
rect 531834 460938 531866 461174
rect 532102 460938 532186 461174
rect 532422 460938 532454 461174
rect 529384 439174 529704 439206
rect 529384 438938 529426 439174
rect 529662 438938 529704 439174
rect 529384 438854 529704 438938
rect 529384 438618 529426 438854
rect 529662 438618 529704 438854
rect 529384 438586 529704 438618
rect 528114 421538 528146 421774
rect 528382 421538 528466 421774
rect 528702 421538 528734 421774
rect 528114 421454 528734 421538
rect 528114 421218 528146 421454
rect 528382 421218 528466 421454
rect 528702 421218 528734 421454
rect 528114 385774 528734 421218
rect 528114 385538 528146 385774
rect 528382 385538 528466 385774
rect 528702 385538 528734 385774
rect 528114 385454 528734 385538
rect 528114 385218 528146 385454
rect 528382 385218 528466 385454
rect 528702 385218 528734 385454
rect 528114 349774 528734 385218
rect 528114 349538 528146 349774
rect 528382 349538 528466 349774
rect 528702 349538 528734 349774
rect 528114 349454 528734 349538
rect 528114 349218 528146 349454
rect 528382 349218 528466 349454
rect 528702 349218 528734 349454
rect 526299 320108 526365 320109
rect 526299 320044 526300 320108
rect 526364 320044 526365 320108
rect 526299 320043 526365 320044
rect 524394 309818 524426 310054
rect 524662 309818 524746 310054
rect 524982 309818 525014 310054
rect 524394 309734 525014 309818
rect 524394 309498 524426 309734
rect 524662 309498 524746 309734
rect 524982 309498 525014 309734
rect 524394 274054 525014 309498
rect 524394 273818 524426 274054
rect 524662 273818 524746 274054
rect 524982 273818 525014 274054
rect 524394 273734 525014 273818
rect 524394 273498 524426 273734
rect 524662 273498 524746 273734
rect 524982 273498 525014 273734
rect 524394 259417 525014 273498
rect 528114 313774 528734 349218
rect 528114 313538 528146 313774
rect 528382 313538 528466 313774
rect 528702 313538 528734 313774
rect 528114 313454 528734 313538
rect 528114 313218 528146 313454
rect 528382 313218 528466 313454
rect 528702 313218 528734 313454
rect 528114 277774 528734 313218
rect 528114 277538 528146 277774
rect 528382 277538 528466 277774
rect 528702 277538 528734 277774
rect 528114 277454 528734 277538
rect 528114 277218 528146 277454
rect 528382 277218 528466 277454
rect 528702 277218 528734 277454
rect 528114 259417 528734 277218
rect 531834 425494 532454 460938
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 460836 542414 470898
rect 545514 705798 546134 711590
rect 545514 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 546134 705798
rect 545514 705478 546134 705562
rect 545514 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 546134 705478
rect 545514 691174 546134 705242
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 537825 439174 538145 439206
rect 537825 438938 537867 439174
rect 538103 438938 538145 439174
rect 537825 438854 538145 438938
rect 537825 438618 537867 438854
rect 538103 438618 538145 438854
rect 537825 438586 538145 438618
rect 545514 439174 546134 474618
rect 549234 706758 549854 711590
rect 549234 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 549854 706758
rect 549234 706438 549854 706522
rect 549234 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 549854 706438
rect 549234 694894 549854 706202
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 533605 435454 533925 435486
rect 533605 435218 533647 435454
rect 533883 435218 533925 435454
rect 533605 435134 533925 435218
rect 533605 434898 533647 435134
rect 533883 434898 533925 435134
rect 533605 434866 533925 434898
rect 542046 435454 542366 435486
rect 542046 435218 542088 435454
rect 542324 435218 542366 435454
rect 542046 435134 542366 435218
rect 542046 434898 542088 435134
rect 542324 434898 542366 435134
rect 542046 434866 542366 434898
rect 531834 425258 531866 425494
rect 532102 425258 532186 425494
rect 532422 425258 532454 425494
rect 531834 425174 532454 425258
rect 531834 424938 531866 425174
rect 532102 424938 532186 425174
rect 532422 424938 532454 425174
rect 531834 389494 532454 424938
rect 531834 389258 531866 389494
rect 532102 389258 532186 389494
rect 532422 389258 532454 389494
rect 531834 389174 532454 389258
rect 531834 388938 531866 389174
rect 532102 388938 532186 389174
rect 532422 388938 532454 389174
rect 531834 353494 532454 388938
rect 531834 353258 531866 353494
rect 532102 353258 532186 353494
rect 532422 353258 532454 353494
rect 531834 353174 532454 353258
rect 531834 352938 531866 353174
rect 532102 352938 532186 353174
rect 532422 352938 532454 353174
rect 531834 317494 532454 352938
rect 531834 317258 531866 317494
rect 532102 317258 532186 317494
rect 532422 317258 532454 317494
rect 531834 317174 532454 317258
rect 531834 316938 531866 317174
rect 532102 316938 532186 317174
rect 532422 316938 532454 317174
rect 531834 281494 532454 316938
rect 541794 399454 542414 425068
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 538259 313988 538325 313989
rect 538259 313924 538260 313988
rect 538324 313924 538325 313988
rect 538259 313923 538325 313924
rect 531834 281258 531866 281494
rect 532102 281258 532186 281494
rect 532422 281258 532454 281494
rect 531834 281174 532454 281258
rect 531834 280938 531866 281174
rect 532102 280938 532186 281174
rect 532422 280938 532454 281174
rect 479568 259174 479888 259206
rect 479568 258938 479610 259174
rect 479846 258938 479888 259174
rect 479568 258854 479888 258938
rect 479568 258618 479610 258854
rect 479846 258618 479888 258854
rect 479568 258586 479888 258618
rect 510288 259174 510608 259206
rect 510288 258938 510330 259174
rect 510566 258938 510608 259174
rect 510288 258854 510608 258938
rect 510288 258618 510330 258854
rect 510566 258618 510608 258854
rect 510288 258586 510608 258618
rect 464208 255454 464528 255486
rect 464208 255218 464250 255454
rect 464486 255218 464528 255454
rect 464208 255134 464528 255218
rect 464208 254898 464250 255134
rect 464486 254898 464528 255134
rect 464208 254866 464528 254898
rect 494928 255454 495248 255486
rect 494928 255218 494970 255454
rect 495206 255218 495248 255454
rect 494928 255134 495248 255218
rect 494928 254898 494970 255134
rect 495206 254898 495248 255134
rect 494928 254866 495248 254898
rect 525648 255454 525968 255486
rect 525648 255218 525690 255454
rect 525926 255218 525968 255454
rect 525648 255134 525968 255218
rect 525648 254898 525690 255134
rect 525926 254898 525968 255134
rect 525648 254866 525968 254898
rect 459834 245258 459866 245494
rect 460102 245258 460186 245494
rect 460422 245258 460454 245494
rect 459834 245174 460454 245258
rect 459834 244938 459866 245174
rect 460102 244938 460186 245174
rect 460422 244938 460454 245174
rect 459834 209494 460454 244938
rect 531834 245494 532454 280938
rect 531834 245258 531866 245494
rect 532102 245258 532186 245494
rect 532422 245258 532454 245494
rect 531834 245174 532454 245258
rect 531834 244938 531866 245174
rect 532102 244938 532186 245174
rect 532422 244938 532454 245174
rect 479568 223174 479888 223206
rect 479568 222938 479610 223174
rect 479846 222938 479888 223174
rect 479568 222854 479888 222938
rect 479568 222618 479610 222854
rect 479846 222618 479888 222854
rect 479568 222586 479888 222618
rect 510288 223174 510608 223206
rect 510288 222938 510330 223174
rect 510566 222938 510608 223174
rect 510288 222854 510608 222938
rect 510288 222618 510330 222854
rect 510566 222618 510608 222854
rect 510288 222586 510608 222618
rect 464208 219454 464528 219486
rect 464208 219218 464250 219454
rect 464486 219218 464528 219454
rect 464208 219134 464528 219218
rect 464208 218898 464250 219134
rect 464486 218898 464528 219134
rect 464208 218866 464528 218898
rect 494928 219454 495248 219486
rect 494928 219218 494970 219454
rect 495206 219218 495248 219454
rect 494928 219134 495248 219218
rect 494928 218898 494970 219134
rect 495206 218898 495248 219134
rect 494928 218866 495248 218898
rect 525648 219454 525968 219486
rect 525648 219218 525690 219454
rect 525926 219218 525968 219454
rect 525648 219134 525968 219218
rect 525648 218898 525690 219134
rect 525926 218898 525968 219134
rect 525648 218866 525968 218898
rect 459834 209258 459866 209494
rect 460102 209258 460186 209494
rect 460422 209258 460454 209494
rect 459834 209174 460454 209258
rect 459834 208938 459866 209174
rect 460102 208938 460186 209174
rect 460422 208938 460454 209174
rect 459834 173494 460454 208938
rect 531834 209494 532454 244938
rect 531834 209258 531866 209494
rect 532102 209258 532186 209494
rect 532422 209258 532454 209494
rect 531834 209174 532454 209258
rect 531834 208938 531866 209174
rect 532102 208938 532186 209174
rect 532422 208938 532454 209174
rect 459834 173258 459866 173494
rect 460102 173258 460186 173494
rect 460422 173258 460454 173494
rect 459834 173174 460454 173258
rect 459834 172938 459866 173174
rect 460102 172938 460186 173174
rect 460422 172938 460454 173174
rect 459834 137494 460454 172938
rect 459834 137258 459866 137494
rect 460102 137258 460186 137494
rect 460422 137258 460454 137494
rect 459834 137174 460454 137258
rect 459834 136938 459866 137174
rect 460102 136938 460186 137174
rect 460422 136938 460454 137174
rect 459834 101494 460454 136938
rect 459834 101258 459866 101494
rect 460102 101258 460186 101494
rect 460422 101258 460454 101494
rect 459834 101174 460454 101258
rect 459834 100938 459866 101174
rect 460102 100938 460186 101174
rect 460422 100938 460454 101174
rect 405568 79174 405888 79206
rect 405568 78938 405610 79174
rect 405846 78938 405888 79174
rect 405568 78854 405888 78938
rect 405568 78618 405610 78854
rect 405846 78618 405888 78854
rect 405568 78586 405888 78618
rect 436288 79174 436608 79206
rect 436288 78938 436330 79174
rect 436566 78938 436608 79174
rect 436288 78854 436608 78938
rect 436288 78618 436330 78854
rect 436566 78618 436608 78854
rect 436288 78586 436608 78618
rect 390208 75454 390528 75486
rect 390208 75218 390250 75454
rect 390486 75218 390528 75454
rect 390208 75134 390528 75218
rect 390208 74898 390250 75134
rect 390486 74898 390528 75134
rect 390208 74866 390528 74898
rect 420928 75454 421248 75486
rect 420928 75218 420970 75454
rect 421206 75218 421248 75454
rect 420928 75134 421248 75218
rect 420928 74898 420970 75134
rect 421206 74898 421248 75134
rect 420928 74866 421248 74898
rect 451648 75454 451968 75486
rect 451648 75218 451690 75454
rect 451926 75218 451968 75454
rect 451648 75134 451968 75218
rect 451648 74898 451690 75134
rect 451926 74898 451968 75134
rect 451648 74866 451968 74898
rect 384114 61538 384146 61774
rect 384382 61538 384466 61774
rect 384702 61538 384734 61774
rect 384114 61454 384734 61538
rect 384114 61218 384146 61454
rect 384382 61218 384466 61454
rect 384702 61218 384734 61454
rect 381491 44844 381557 44845
rect 381491 44780 381492 44844
rect 381556 44780 381557 44844
rect 381491 44779 381557 44780
rect 380394 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 381014 22054
rect 380394 21734 381014 21818
rect 380394 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 381014 21734
rect 380394 -5146 381014 21498
rect 380394 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 381014 -5146
rect 380394 -5466 381014 -5382
rect 380394 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 381014 -5466
rect 380394 -7654 381014 -5702
rect 384114 25774 384734 61218
rect 459834 65494 460454 100938
rect 459834 65258 459866 65494
rect 460102 65258 460186 65494
rect 460422 65258 460454 65494
rect 459834 65174 460454 65258
rect 459834 64938 459866 65174
rect 460102 64938 460186 65174
rect 460422 64938 460454 65174
rect 405568 43174 405888 43206
rect 405568 42938 405610 43174
rect 405846 42938 405888 43174
rect 405568 42854 405888 42938
rect 405568 42618 405610 42854
rect 405846 42618 405888 42854
rect 405568 42586 405888 42618
rect 436288 43174 436608 43206
rect 436288 42938 436330 43174
rect 436566 42938 436608 43174
rect 436288 42854 436608 42938
rect 436288 42618 436330 42854
rect 436566 42618 436608 42854
rect 436288 42586 436608 42618
rect 390208 39454 390528 39486
rect 390208 39218 390250 39454
rect 390486 39218 390528 39454
rect 390208 39134 390528 39218
rect 390208 38898 390250 39134
rect 390486 38898 390528 39134
rect 390208 38866 390528 38898
rect 420928 39454 421248 39486
rect 420928 39218 420970 39454
rect 421206 39218 421248 39454
rect 420928 39134 421248 39218
rect 420928 38898 420970 39134
rect 421206 38898 421248 39134
rect 420928 38866 421248 38898
rect 451648 39454 451968 39486
rect 451648 39218 451690 39454
rect 451926 39218 451968 39454
rect 451648 39134 451968 39218
rect 451648 38898 451690 39134
rect 451926 38898 451968 39134
rect 451648 38866 451968 38898
rect 384114 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 384734 25774
rect 384114 25454 384734 25538
rect 384114 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 384734 25454
rect 384114 -6106 384734 25218
rect 384114 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 384734 -6106
rect 384114 -6426 384734 -6342
rect 384114 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 384734 -6426
rect 384114 -7654 384734 -6662
rect 387834 29494 388454 31919
rect 387834 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 388454 29494
rect 387834 29174 388454 29258
rect 387834 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 388454 29174
rect 387834 -7066 388454 28938
rect 387834 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 388454 -7066
rect 387834 -7386 388454 -7302
rect 387834 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 388454 -7386
rect 387834 -7654 388454 -7622
rect 397794 3454 398414 31919
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 401514 7174 402134 31919
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -1306 402134 6618
rect 401514 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 402134 -1306
rect 401514 -1626 402134 -1542
rect 401514 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 402134 -1626
rect 401514 -7654 402134 -1862
rect 405234 10894 405854 30068
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -2266 405854 10338
rect 405234 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 405854 -2266
rect 405234 -2586 405854 -2502
rect 405234 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 405854 -2586
rect 405234 -7654 405854 -2822
rect 408954 14614 409574 31919
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 408954 -3226 409574 14058
rect 408954 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 409574 -3226
rect 408954 -3546 409574 -3462
rect 408954 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 409574 -3546
rect 408954 -7654 409574 -3782
rect 412674 18334 413294 31919
rect 412674 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 413294 18334
rect 412674 18014 413294 18098
rect 412674 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 413294 18014
rect 412674 -4186 413294 17778
rect 412674 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 413294 -4186
rect 412674 -4506 413294 -4422
rect 412674 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 413294 -4506
rect 412674 -7654 413294 -4742
rect 416394 22054 417014 31919
rect 416394 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 417014 22054
rect 416394 21734 417014 21818
rect 416394 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 417014 21734
rect 416394 -5146 417014 21498
rect 416394 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 417014 -5146
rect 416394 -5466 417014 -5382
rect 416394 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 417014 -5466
rect 416394 -7654 417014 -5702
rect 420114 25774 420734 31919
rect 420114 25538 420146 25774
rect 420382 25538 420466 25774
rect 420702 25538 420734 25774
rect 420114 25454 420734 25538
rect 420114 25218 420146 25454
rect 420382 25218 420466 25454
rect 420702 25218 420734 25454
rect 420114 -6106 420734 25218
rect 420114 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 420734 -6106
rect 420114 -6426 420734 -6342
rect 420114 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 420734 -6426
rect 420114 -7654 420734 -6662
rect 423834 29494 424454 31919
rect 423834 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 424454 29494
rect 423834 29174 424454 29258
rect 423834 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 424454 29174
rect 423834 -7066 424454 28938
rect 423834 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 424454 -7066
rect 423834 -7386 424454 -7302
rect 423834 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 424454 -7386
rect 423834 -7654 424454 -7622
rect 433794 3454 434414 31919
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 437514 7174 438134 31919
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -1306 438134 6618
rect 437514 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 438134 -1306
rect 437514 -1626 438134 -1542
rect 437514 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 438134 -1626
rect 437514 -7654 438134 -1862
rect 441234 10894 441854 31919
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -2266 441854 10338
rect 441234 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 441854 -2266
rect 441234 -2586 441854 -2502
rect 441234 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 441854 -2586
rect 441234 -7654 441854 -2822
rect 444954 14614 445574 31919
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 444954 -3226 445574 14058
rect 444954 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 445574 -3226
rect 444954 -3546 445574 -3462
rect 444954 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 445574 -3546
rect 444954 -7654 445574 -3782
rect 448674 18334 449294 31919
rect 448674 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 449294 18334
rect 448674 18014 449294 18098
rect 448674 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 449294 18014
rect 448674 -4186 449294 17778
rect 448674 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 449294 -4186
rect 448674 -4506 449294 -4422
rect 448674 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 449294 -4506
rect 448674 -7654 449294 -4742
rect 452394 22054 453014 31919
rect 452394 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 453014 22054
rect 452394 21734 453014 21818
rect 452394 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 453014 21734
rect 452394 -5146 453014 21498
rect 452394 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 453014 -5146
rect 452394 -5466 453014 -5382
rect 452394 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 453014 -5466
rect 452394 -7654 453014 -5702
rect 456114 25774 456734 31919
rect 456114 25538 456146 25774
rect 456382 25538 456466 25774
rect 456702 25538 456734 25774
rect 456114 25454 456734 25538
rect 456114 25218 456146 25454
rect 456382 25218 456466 25454
rect 456702 25218 456734 25454
rect 456114 -6106 456734 25218
rect 456114 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 456734 -6106
rect 456114 -6426 456734 -6342
rect 456114 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 456734 -6426
rect 456114 -7654 456734 -6662
rect 459834 29494 460454 64938
rect 459834 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 460454 29494
rect 459834 29174 460454 29258
rect 459834 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 460454 29174
rect 459834 -7066 460454 28938
rect 459834 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 460454 -7066
rect 459834 -7386 460454 -7302
rect 459834 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 460454 -7386
rect 459834 -7654 460454 -7622
rect 469794 183454 470414 201919
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 473514 187174 474134 201919
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -1306 474134 6618
rect 473514 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 474134 -1306
rect 473514 -1626 474134 -1542
rect 473514 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 474134 -1626
rect 473514 -7654 474134 -1862
rect 477234 190894 477854 201919
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -2266 477854 10338
rect 477234 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 477854 -2266
rect 477234 -2586 477854 -2502
rect 477234 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 477854 -2586
rect 477234 -7654 477854 -2822
rect 480954 194614 481574 201919
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 484674 198334 485294 201919
rect 484674 198098 484706 198334
rect 484942 198098 485026 198334
rect 485262 198098 485294 198334
rect 484674 198014 485294 198098
rect 484674 197778 484706 198014
rect 484942 197778 485026 198014
rect 485262 197778 485294 198014
rect 484674 162334 485294 197778
rect 484674 162098 484706 162334
rect 484942 162098 485026 162334
rect 485262 162098 485294 162334
rect 484674 162014 485294 162098
rect 484674 161778 484706 162014
rect 484942 161778 485026 162014
rect 485262 161778 485294 162014
rect 484674 126334 485294 161778
rect 484674 126098 484706 126334
rect 484942 126098 485026 126334
rect 485262 126098 485294 126334
rect 484674 126014 485294 126098
rect 484674 125778 484706 126014
rect 484942 125778 485026 126014
rect 485262 125778 485294 126014
rect 484208 111454 484528 111486
rect 484208 111218 484250 111454
rect 484486 111218 484528 111454
rect 484208 111134 484528 111218
rect 484208 110898 484250 111134
rect 484486 110898 484528 111134
rect 484208 110866 484528 110898
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 480954 -3226 481574 14058
rect 480954 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 481574 -3226
rect 480954 -3546 481574 -3462
rect 480954 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 481574 -3546
rect 480954 -7654 481574 -3782
rect 484674 90334 485294 125778
rect 484674 90098 484706 90334
rect 484942 90098 485026 90334
rect 485262 90098 485294 90334
rect 484674 90014 485294 90098
rect 484674 89778 484706 90014
rect 484942 89778 485026 90014
rect 485262 89778 485294 90014
rect 484674 54334 485294 89778
rect 484674 54098 484706 54334
rect 484942 54098 485026 54334
rect 485262 54098 485294 54334
rect 484674 54014 485294 54098
rect 484674 53778 484706 54014
rect 484942 53778 485026 54014
rect 485262 53778 485294 54014
rect 484674 18334 485294 53778
rect 484674 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 485294 18334
rect 484674 18014 485294 18098
rect 484674 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 485294 18014
rect 484674 -4186 485294 17778
rect 484674 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 485294 -4186
rect 484674 -4506 485294 -4422
rect 484674 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 485294 -4506
rect 484674 -7654 485294 -4742
rect 488394 166054 489014 201919
rect 488394 165818 488426 166054
rect 488662 165818 488746 166054
rect 488982 165818 489014 166054
rect 488394 165734 489014 165818
rect 488394 165498 488426 165734
rect 488662 165498 488746 165734
rect 488982 165498 489014 165734
rect 488394 130054 489014 165498
rect 505794 183454 506414 201919
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 139417 506414 146898
rect 509514 187174 510134 201919
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 139417 510134 150618
rect 513234 190894 513854 201919
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 139417 513854 154338
rect 516954 194614 517574 201919
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 139417 517574 158058
rect 520674 198334 521294 201919
rect 520674 198098 520706 198334
rect 520942 198098 521026 198334
rect 521262 198098 521294 198334
rect 520674 198014 521294 198098
rect 520674 197778 520706 198014
rect 520942 197778 521026 198014
rect 521262 197778 521294 198014
rect 520674 162334 521294 197778
rect 520674 162098 520706 162334
rect 520942 162098 521026 162334
rect 521262 162098 521294 162334
rect 520674 162014 521294 162098
rect 520674 161778 520706 162014
rect 520942 161778 521026 162014
rect 521262 161778 521294 162014
rect 520674 139417 521294 161778
rect 524394 166054 525014 201919
rect 524394 165818 524426 166054
rect 524662 165818 524746 166054
rect 524982 165818 525014 166054
rect 524394 165734 525014 165818
rect 524394 165498 524426 165734
rect 524662 165498 524746 165734
rect 524982 165498 525014 165734
rect 524394 139417 525014 165498
rect 531834 173494 532454 208938
rect 531834 173258 531866 173494
rect 532102 173258 532186 173494
rect 532422 173258 532454 173494
rect 531834 173174 532454 173258
rect 531834 172938 531866 173174
rect 532102 172938 532186 173174
rect 532422 172938 532454 173174
rect 531834 139417 532454 172938
rect 538262 151830 538322 313923
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 538262 151770 539426 151830
rect 488394 129818 488426 130054
rect 488662 129818 488746 130054
rect 488982 129818 489014 130054
rect 488394 129734 489014 129818
rect 488394 129498 488426 129734
rect 488662 129498 488746 129734
rect 488982 129498 489014 129734
rect 488394 94054 489014 129498
rect 539366 129301 539426 151770
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 539363 129300 539429 129301
rect 539363 129236 539364 129300
rect 539428 129236 539429 129300
rect 539363 129235 539429 129236
rect 499568 115174 499888 115206
rect 499568 114938 499610 115174
rect 499846 114938 499888 115174
rect 499568 114854 499888 114938
rect 499568 114618 499610 114854
rect 499846 114618 499888 114854
rect 499568 114586 499888 114618
rect 530288 115174 530608 115206
rect 530288 114938 530330 115174
rect 530566 114938 530608 115174
rect 530288 114854 530608 114938
rect 530288 114618 530330 114854
rect 530566 114618 530608 114854
rect 530288 114586 530608 114618
rect 514928 111454 515248 111486
rect 514928 111218 514970 111454
rect 515206 111218 515248 111454
rect 514928 111134 515248 111218
rect 514928 110898 514970 111134
rect 515206 110898 515248 111134
rect 514928 110866 515248 110898
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 488394 93818 488426 94054
rect 488662 93818 488746 94054
rect 488982 93818 489014 94054
rect 488394 93734 489014 93818
rect 488394 93498 488426 93734
rect 488662 93498 488746 93734
rect 488982 93498 489014 93734
rect 488394 58054 489014 93498
rect 488394 57818 488426 58054
rect 488662 57818 488746 58054
rect 488982 57818 489014 58054
rect 488394 57734 489014 57818
rect 488394 57498 488426 57734
rect 488662 57498 488746 57734
rect 488982 57498 489014 57734
rect 488394 22054 489014 57498
rect 488394 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 489014 22054
rect 488394 21734 489014 21818
rect 488394 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 489014 21734
rect 488394 -5146 489014 21498
rect 488394 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 489014 -5146
rect 488394 -5466 489014 -5382
rect 488394 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 489014 -5466
rect 488394 -7654 489014 -5702
rect 492114 61774 492734 83687
rect 492114 61538 492146 61774
rect 492382 61538 492466 61774
rect 492702 61538 492734 61774
rect 492114 61454 492734 61538
rect 492114 61218 492146 61454
rect 492382 61218 492466 61454
rect 492702 61218 492734 61454
rect 492114 25774 492734 61218
rect 492114 25538 492146 25774
rect 492382 25538 492466 25774
rect 492702 25538 492734 25774
rect 492114 25454 492734 25538
rect 492114 25218 492146 25454
rect 492382 25218 492466 25454
rect 492702 25218 492734 25454
rect 492114 -6106 492734 25218
rect 492114 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 492734 -6106
rect 492114 -6426 492734 -6342
rect 492114 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 492734 -6426
rect 492114 -7654 492734 -6662
rect 495834 65494 496454 83687
rect 495834 65258 495866 65494
rect 496102 65258 496186 65494
rect 496422 65258 496454 65494
rect 495834 65174 496454 65258
rect 495834 64938 495866 65174
rect 496102 64938 496186 65174
rect 496422 64938 496454 65174
rect 495834 29494 496454 64938
rect 495834 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 496454 29494
rect 495834 29174 496454 29258
rect 495834 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 496454 29174
rect 495834 -7066 496454 28938
rect 495834 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 496454 -7066
rect 495834 -7386 496454 -7302
rect 495834 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 496454 -7386
rect 495834 -7654 496454 -7622
rect 505794 75454 506414 83687
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 509514 79174 510134 83687
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -1306 510134 6618
rect 509514 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 510134 -1306
rect 509514 -1626 510134 -1542
rect 509514 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 510134 -1626
rect 509514 -7654 510134 -1862
rect 513234 82894 513854 83687
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -2266 513854 10338
rect 513234 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 513854 -2266
rect 513234 -2586 513854 -2502
rect 513234 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 513854 -2586
rect 513234 -7654 513854 -2822
rect 516954 50614 517574 83687
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 516954 -3226 517574 14058
rect 516954 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 517574 -3226
rect 516954 -3546 517574 -3462
rect 516954 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 517574 -3546
rect 516954 -7654 517574 -3782
rect 520674 54334 521294 83687
rect 520674 54098 520706 54334
rect 520942 54098 521026 54334
rect 521262 54098 521294 54334
rect 520674 54014 521294 54098
rect 520674 53778 520706 54014
rect 520942 53778 521026 54014
rect 521262 53778 521294 54014
rect 520674 18334 521294 53778
rect 520674 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 521294 18334
rect 520674 18014 521294 18098
rect 520674 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 521294 18014
rect 520674 -4186 521294 17778
rect 520674 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 521294 -4186
rect 520674 -4506 521294 -4422
rect 520674 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 521294 -4506
rect 520674 -7654 521294 -4742
rect 524394 58054 525014 83687
rect 524394 57818 524426 58054
rect 524662 57818 524746 58054
rect 524982 57818 525014 58054
rect 524394 57734 525014 57818
rect 524394 57498 524426 57734
rect 524662 57498 524746 57734
rect 524982 57498 525014 57734
rect 524394 22054 525014 57498
rect 524394 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 525014 22054
rect 524394 21734 525014 21818
rect 524394 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 525014 21734
rect 524394 -5146 525014 21498
rect 524394 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 525014 -5146
rect 524394 -5466 525014 -5382
rect 524394 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 525014 -5466
rect 524394 -7654 525014 -5702
rect 528114 61774 528734 83687
rect 528114 61538 528146 61774
rect 528382 61538 528466 61774
rect 528702 61538 528734 61774
rect 528114 61454 528734 61538
rect 528114 61218 528146 61454
rect 528382 61218 528466 61454
rect 528702 61218 528734 61454
rect 528114 25774 528734 61218
rect 528114 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 528734 25774
rect 528114 25454 528734 25538
rect 528114 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 528734 25454
rect 528114 -6106 528734 25218
rect 528114 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 528734 -6106
rect 528114 -6426 528734 -6342
rect 528114 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 528734 -6426
rect 528114 -7654 528734 -6662
rect 531834 65494 532454 83687
rect 531834 65258 531866 65494
rect 532102 65258 532186 65494
rect 532422 65258 532454 65494
rect 531834 65174 532454 65258
rect 531834 64938 531866 65174
rect 532102 64938 532186 65174
rect 532422 64938 532454 65174
rect 531834 29494 532454 64938
rect 531834 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 532454 29494
rect 531834 29174 532454 29258
rect 531834 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 532454 29174
rect 531834 -7066 532454 28938
rect 531834 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 532454 -7066
rect 531834 -7386 532454 -7302
rect 531834 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 532454 -7386
rect 531834 -7654 532454 -7622
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 545514 403174 546134 438618
rect 546266 439174 546586 439206
rect 546266 438938 546308 439174
rect 546544 438938 546586 439174
rect 546266 438854 546586 438938
rect 546266 438618 546308 438854
rect 546544 438618 546586 438854
rect 546266 438586 546586 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 51692 546134 78618
rect 549234 406894 549854 442338
rect 552954 707718 553574 711590
rect 552954 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 553574 707718
rect 552954 707398 553574 707482
rect 552954 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 553574 707398
rect 552954 698614 553574 707162
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 550487 435454 550807 435486
rect 550487 435218 550529 435454
rect 550765 435218 550807 435454
rect 550487 435134 550807 435218
rect 550487 434898 550529 435134
rect 550765 434898 550807 435134
rect 550487 434866 550807 434898
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 552954 410614 553574 446058
rect 556674 708678 557294 711590
rect 556674 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 557294 708678
rect 556674 708358 557294 708442
rect 556674 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 557294 708358
rect 556674 666334 557294 708122
rect 560394 709638 561014 711590
rect 560394 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 561014 709638
rect 560394 709318 561014 709402
rect 560394 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 561014 709318
rect 559419 699820 559485 699821
rect 559419 699756 559420 699820
rect 559484 699756 559485 699820
rect 559419 699755 559485 699756
rect 556674 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 557294 666334
rect 556674 666014 557294 666098
rect 556674 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 557294 666014
rect 556674 630334 557294 665778
rect 556674 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 557294 630334
rect 556674 630014 557294 630098
rect 556674 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 557294 630014
rect 556674 594334 557294 629778
rect 556674 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 557294 594334
rect 556674 594014 557294 594098
rect 556674 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 557294 594014
rect 556674 558334 557294 593778
rect 556674 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 557294 558334
rect 556674 558014 557294 558098
rect 556674 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 557294 558014
rect 556674 522334 557294 557778
rect 556674 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 557294 522334
rect 556674 522014 557294 522098
rect 556674 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 557294 522014
rect 556674 486334 557294 521778
rect 556674 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 557294 486334
rect 556674 486014 557294 486098
rect 556674 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 557294 486014
rect 556674 450334 557294 485778
rect 556674 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 557294 450334
rect 556674 450014 557294 450098
rect 556674 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 557294 450014
rect 554707 439174 555027 439206
rect 554707 438938 554749 439174
rect 554985 438938 555027 439174
rect 554707 438854 555027 438938
rect 554707 438618 554749 438854
rect 554985 438618 555027 438854
rect 554707 438586 555027 438618
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 377884 553574 410058
rect 556674 414334 557294 449778
rect 556674 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 557294 414334
rect 556674 414014 557294 414098
rect 556674 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 557294 414014
rect 556674 378243 557294 413778
rect 556674 378007 556706 378243
rect 556942 378007 557026 378243
rect 557262 378007 557294 378243
rect 556674 377884 557294 378007
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 554876 367174 555196 367206
rect 554876 366938 554918 367174
rect 555154 366938 555196 367174
rect 554876 366854 555196 366938
rect 554876 366618 554918 366854
rect 555154 366618 555196 366854
rect 554876 366586 555196 366618
rect 558809 367174 559129 367206
rect 558809 366938 558851 367174
rect 559087 366938 559129 367174
rect 558809 366854 559129 366938
rect 558809 366618 558851 366854
rect 559087 366618 559129 366854
rect 558809 366586 559129 366618
rect 552910 363454 553230 363486
rect 552910 363218 552952 363454
rect 553188 363218 553230 363454
rect 552910 363134 553230 363218
rect 552910 362898 552952 363134
rect 553188 362898 553230 363134
rect 552910 362866 553230 362898
rect 556843 363454 557163 363486
rect 556843 363218 556885 363454
rect 557121 363218 557163 363454
rect 556843 363134 557163 363218
rect 556843 362898 556885 363134
rect 557121 362898 557163 363134
rect 556843 362866 557163 362898
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 552954 338614 553574 360068
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 51692 553574 86058
rect 556674 342334 557294 360068
rect 556674 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 557294 342334
rect 556674 342014 557294 342098
rect 556674 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 557294 342014
rect 556674 306334 557294 341778
rect 559422 321469 559482 699755
rect 560394 670054 561014 709082
rect 560394 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 561014 670054
rect 560394 669734 561014 669818
rect 560394 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 561014 669734
rect 560394 634054 561014 669498
rect 560394 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 561014 634054
rect 560394 633734 561014 633818
rect 560394 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 561014 633734
rect 560394 598054 561014 633498
rect 560394 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 561014 598054
rect 560394 597734 561014 597818
rect 560394 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 561014 597734
rect 560394 562054 561014 597498
rect 560394 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 561014 562054
rect 560394 561734 561014 561818
rect 560394 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 561014 561734
rect 560394 526054 561014 561498
rect 560394 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 561014 526054
rect 560394 525734 561014 525818
rect 560394 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 561014 525734
rect 560394 490054 561014 525498
rect 560394 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 561014 490054
rect 560394 489734 561014 489818
rect 560394 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 561014 489734
rect 560394 454054 561014 489498
rect 560394 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 561014 454054
rect 560394 453734 561014 453818
rect 560394 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 561014 453734
rect 560394 418054 561014 453498
rect 560394 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 561014 418054
rect 560394 417734 561014 417818
rect 560394 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 561014 417734
rect 560394 382054 561014 417498
rect 560394 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 561014 382054
rect 560394 381734 561014 381818
rect 560394 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 561014 381734
rect 560394 377884 561014 381498
rect 564114 710598 564734 711590
rect 564114 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 564734 710598
rect 564114 710278 564734 710362
rect 564114 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 564734 710278
rect 564114 673774 564734 710042
rect 564114 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 564734 673774
rect 564114 673454 564734 673538
rect 564114 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 564734 673454
rect 564114 637774 564734 673218
rect 564114 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 564734 637774
rect 564114 637454 564734 637538
rect 564114 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 564734 637454
rect 564114 601774 564734 637218
rect 564114 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 564734 601774
rect 564114 601454 564734 601538
rect 564114 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 564734 601454
rect 564114 565774 564734 601218
rect 564114 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 564734 565774
rect 564114 565454 564734 565538
rect 564114 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 564734 565454
rect 564114 529774 564734 565218
rect 564114 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 564734 529774
rect 564114 529454 564734 529538
rect 564114 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 564734 529454
rect 564114 493774 564734 529218
rect 564114 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 564734 493774
rect 564114 493454 564734 493538
rect 564114 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 564734 493454
rect 564114 457774 564734 493218
rect 564114 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 564734 457774
rect 564114 457454 564734 457538
rect 564114 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 564734 457454
rect 564114 421774 564734 457218
rect 564114 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 564734 421774
rect 564114 421454 564734 421538
rect 564114 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 564734 421454
rect 564114 385774 564734 421218
rect 564114 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 564734 385774
rect 564114 385454 564734 385538
rect 564114 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 564734 385454
rect 564114 377884 564734 385218
rect 567834 711558 568454 711590
rect 567834 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 568454 711558
rect 567834 711238 568454 711322
rect 567834 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 568454 711238
rect 567834 677494 568454 711002
rect 567834 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 568454 677494
rect 567834 677174 568454 677258
rect 567834 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 568454 677174
rect 567834 641494 568454 676938
rect 567834 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 568454 641494
rect 567834 641174 568454 641258
rect 567834 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 568454 641174
rect 567834 605494 568454 640938
rect 567834 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 568454 605494
rect 567834 605174 568454 605258
rect 567834 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 568454 605174
rect 567834 569494 568454 604938
rect 567834 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 568454 569494
rect 567834 569174 568454 569258
rect 567834 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 568454 569174
rect 567834 533494 568454 568938
rect 567834 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 568454 533494
rect 567834 533174 568454 533258
rect 567834 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 568454 533174
rect 567834 497494 568454 532938
rect 567834 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 568454 497494
rect 567834 497174 568454 497258
rect 567834 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 568454 497174
rect 567834 461494 568454 496938
rect 567834 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 568454 461494
rect 567834 461174 568454 461258
rect 567834 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 568454 461174
rect 567834 425494 568454 460938
rect 567834 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 568454 425494
rect 567834 425174 568454 425258
rect 567834 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 568454 425174
rect 567834 389494 568454 424938
rect 567834 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 568454 389494
rect 567834 389174 568454 389258
rect 567834 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 568454 389174
rect 562742 367174 563062 367206
rect 562742 366938 562784 367174
rect 563020 366938 563062 367174
rect 562742 366854 563062 366938
rect 562742 366618 562784 366854
rect 563020 366618 563062 366854
rect 562742 366586 563062 366618
rect 566675 367174 566995 367206
rect 566675 366938 566717 367174
rect 566953 366938 566995 367174
rect 566675 366854 566995 366938
rect 566675 366618 566717 366854
rect 566953 366618 566995 366854
rect 566675 366586 566995 366618
rect 560776 363454 561096 363486
rect 560776 363218 560818 363454
rect 561054 363218 561096 363454
rect 560776 363134 561096 363218
rect 560776 362898 560818 363134
rect 561054 362898 561096 363134
rect 560776 362866 561096 362898
rect 564709 363454 565029 363486
rect 564709 363218 564751 363454
rect 564987 363218 565029 363454
rect 564709 363134 565029 363218
rect 564709 362898 564751 363134
rect 564987 362898 565029 363134
rect 564709 362866 565029 362898
rect 560394 346054 561014 360068
rect 560394 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 561014 346054
rect 560394 345734 561014 345818
rect 560394 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 561014 345734
rect 559419 321468 559485 321469
rect 559419 321404 559420 321468
rect 559484 321404 559485 321468
rect 559419 321403 559485 321404
rect 556674 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 557294 306334
rect 556674 306014 557294 306098
rect 556674 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 557294 306014
rect 556674 270334 557294 305778
rect 556674 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 557294 270334
rect 556674 270014 557294 270098
rect 556674 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 557294 270014
rect 556674 234334 557294 269778
rect 556674 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 557294 234334
rect 556674 234014 557294 234098
rect 556674 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 557294 234014
rect 556674 198334 557294 233778
rect 556674 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 557294 198334
rect 556674 198014 557294 198098
rect 556674 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 557294 198014
rect 556674 162334 557294 197778
rect 556674 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 557294 162334
rect 556674 162014 557294 162098
rect 556674 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 557294 162014
rect 556674 126334 557294 161778
rect 556674 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 557294 126334
rect 556674 126014 557294 126098
rect 556674 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 557294 126014
rect 556674 90334 557294 125778
rect 556674 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 557294 90334
rect 556674 90014 557294 90098
rect 556674 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 557294 90014
rect 556674 54334 557294 89778
rect 556674 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 557294 54334
rect 556674 54014 557294 54098
rect 556674 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 557294 54014
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 545888 43174 546208 43206
rect 545888 42938 545930 43174
rect 546166 42938 546208 43174
rect 545888 42854 546208 42938
rect 545888 42618 545930 42854
rect 546166 42618 546208 42854
rect 545888 42586 546208 42618
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 543416 39454 543736 39486
rect 543416 39218 543458 39454
rect 543694 39218 543736 39454
rect 543416 39134 543736 39218
rect 543416 38898 543458 39134
rect 543694 38898 543736 39134
rect 543416 38866 543736 38898
rect 548361 39454 548681 39486
rect 548361 39218 548403 39454
rect 548639 39218 548681 39454
rect 548361 39134 548681 39218
rect 548361 38898 548403 39134
rect 548639 38898 548681 39134
rect 548361 38866 548681 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 545514 7174 546134 30068
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -1306 546134 6618
rect 545514 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 546134 -1306
rect 545514 -1626 546134 -1542
rect 545514 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 546134 -1626
rect 545514 -7654 546134 -1862
rect 549234 10894 549854 46338
rect 550833 43174 551153 43206
rect 550833 42938 550875 43174
rect 551111 42938 551153 43174
rect 550833 42854 551153 42938
rect 550833 42618 550875 42854
rect 551111 42618 551153 42854
rect 550833 42586 551153 42618
rect 555778 43174 556098 43206
rect 555778 42938 555820 43174
rect 556056 42938 556098 43174
rect 555778 42854 556098 42938
rect 555778 42618 555820 42854
rect 556056 42618 556098 42854
rect 555778 42586 556098 42618
rect 553306 39454 553626 39486
rect 553306 39218 553348 39454
rect 553584 39218 553626 39454
rect 553306 39134 553626 39218
rect 553306 38898 553348 39134
rect 553584 38898 553626 39134
rect 553306 38866 553626 38898
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -2266 549854 10338
rect 549234 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 549854 -2266
rect 549234 -2586 549854 -2502
rect 549234 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 549854 -2586
rect 549234 -7654 549854 -2822
rect 552954 14614 553574 30068
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 552954 -3226 553574 14058
rect 552954 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 553574 -3226
rect 552954 -3546 553574 -3462
rect 552954 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 553574 -3546
rect 552954 -7654 553574 -3782
rect 556674 18334 557294 53778
rect 560394 310054 561014 345498
rect 560394 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 561014 310054
rect 560394 309734 561014 309818
rect 560394 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 561014 309734
rect 560394 274054 561014 309498
rect 560394 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 561014 274054
rect 560394 273734 561014 273818
rect 560394 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 561014 273734
rect 560394 238054 561014 273498
rect 560394 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 561014 238054
rect 560394 237734 561014 237818
rect 560394 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 561014 237734
rect 560394 202054 561014 237498
rect 560394 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 561014 202054
rect 560394 201734 561014 201818
rect 560394 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 561014 201734
rect 560394 166054 561014 201498
rect 560394 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 561014 166054
rect 560394 165734 561014 165818
rect 560394 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 561014 165734
rect 560394 130054 561014 165498
rect 560394 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 561014 130054
rect 560394 129734 561014 129818
rect 560394 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 561014 129734
rect 560394 94054 561014 129498
rect 560394 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 561014 94054
rect 560394 93734 561014 93818
rect 560394 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 561014 93734
rect 560394 58054 561014 93498
rect 560394 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 561014 58054
rect 560394 57734 561014 57818
rect 560394 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 561014 57734
rect 560394 51692 561014 57498
rect 564114 349774 564734 360068
rect 564114 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 564734 349774
rect 564114 349454 564734 349538
rect 564114 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 564734 349454
rect 564114 313774 564734 349218
rect 564114 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 564734 313774
rect 564114 313454 564734 313538
rect 564114 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 564734 313454
rect 564114 277774 564734 313218
rect 564114 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 564734 277774
rect 564114 277454 564734 277538
rect 564114 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 564734 277454
rect 564114 241774 564734 277218
rect 564114 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 564734 241774
rect 564114 241454 564734 241538
rect 564114 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 564734 241454
rect 564114 205774 564734 241218
rect 564114 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 564734 205774
rect 564114 205454 564734 205538
rect 564114 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 564734 205454
rect 564114 169774 564734 205218
rect 564114 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 564734 169774
rect 564114 169454 564734 169538
rect 564114 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 564734 169454
rect 564114 133774 564734 169218
rect 564114 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 564734 133774
rect 564114 133454 564734 133538
rect 564114 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 564734 133454
rect 564114 97774 564734 133218
rect 564114 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 564734 97774
rect 564114 97454 564734 97538
rect 564114 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 564734 97454
rect 564114 61774 564734 97218
rect 564114 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 564734 61774
rect 564114 61454 564734 61538
rect 564114 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 564734 61454
rect 560723 43174 561043 43206
rect 560723 42938 560765 43174
rect 561001 42938 561043 43174
rect 560723 42854 561043 42938
rect 560723 42618 560765 42854
rect 561001 42618 561043 42854
rect 560723 42586 561043 42618
rect 558251 39454 558571 39486
rect 558251 39218 558293 39454
rect 558529 39218 558571 39454
rect 558251 39134 558571 39218
rect 558251 38898 558293 39134
rect 558529 38898 558571 39134
rect 558251 38866 558571 38898
rect 556674 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 557294 18334
rect 556674 18014 557294 18098
rect 556674 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 557294 18014
rect 556674 -4186 557294 17778
rect 556674 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 557294 -4186
rect 556674 -4506 557294 -4422
rect 556674 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 557294 -4506
rect 556674 -7654 557294 -4742
rect 560394 22054 561014 30068
rect 560394 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 561014 22054
rect 560394 21734 561014 21818
rect 560394 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 561014 21734
rect 560394 -5146 561014 21498
rect 560394 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 561014 -5146
rect 560394 -5466 561014 -5382
rect 560394 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 561014 -5466
rect 560394 -7654 561014 -5702
rect 564114 25774 564734 61218
rect 564114 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 564734 25774
rect 564114 25454 564734 25538
rect 564114 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 564734 25454
rect 564114 -6106 564734 25218
rect 564114 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 564734 -6106
rect 564114 -6426 564734 -6342
rect 564114 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 564734 -6426
rect 564114 -7654 564734 -6662
rect 567834 353494 568454 388938
rect 567834 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 568454 353494
rect 567834 353174 568454 353258
rect 567834 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 568454 353174
rect 567834 317494 568454 352938
rect 567834 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 568454 317494
rect 567834 317174 568454 317258
rect 567834 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 568454 317174
rect 567834 281494 568454 316938
rect 567834 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 568454 281494
rect 567834 281174 568454 281258
rect 567834 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 568454 281174
rect 567834 245494 568454 280938
rect 567834 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 568454 245494
rect 567834 245174 568454 245258
rect 567834 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 568454 245174
rect 567834 209494 568454 244938
rect 567834 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 568454 209494
rect 567834 209174 568454 209258
rect 567834 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 568454 209174
rect 567834 173494 568454 208938
rect 567834 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 568454 173494
rect 567834 173174 568454 173258
rect 567834 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 568454 173174
rect 567834 137494 568454 172938
rect 567834 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 568454 137494
rect 567834 137174 568454 137258
rect 567834 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 568454 137174
rect 567834 101494 568454 136938
rect 567834 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 568454 101494
rect 567834 101174 568454 101258
rect 567834 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 568454 101174
rect 567834 65494 568454 100938
rect 567834 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 568454 65494
rect 567834 65174 568454 65258
rect 567834 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 568454 65174
rect 567834 29494 568454 64938
rect 567834 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 568454 29494
rect 567834 29174 568454 29258
rect 567834 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 568454 29174
rect 567834 -7066 568454 28938
rect 567834 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 568454 -7066
rect 567834 -7386 568454 -7302
rect 567834 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 568454 -7386
rect 567834 -7654 568454 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 581514 705798 582134 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 581514 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 582134 705798
rect 581514 705478 582134 705562
rect 581514 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 582134 705478
rect 581514 691174 582134 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -1306 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691174 586890 705242
rect 586270 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 586890 691174
rect 586270 690854 586890 690938
rect 586270 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 586890 690854
rect 586270 655174 586890 690618
rect 586270 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 586890 655174
rect 586270 654854 586890 654938
rect 586270 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 586890 654854
rect 586270 619174 586890 654618
rect 586270 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 586890 619174
rect 586270 618854 586890 618938
rect 586270 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 586890 618854
rect 586270 583174 586890 618618
rect 586270 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 586890 583174
rect 586270 582854 586890 582938
rect 586270 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 586890 582854
rect 586270 547174 586890 582618
rect 586270 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 586890 547174
rect 586270 546854 586890 546938
rect 586270 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 586890 546854
rect 586270 511174 586890 546618
rect 586270 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 586890 511174
rect 586270 510854 586890 510938
rect 586270 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 586890 510854
rect 586270 475174 586890 510618
rect 586270 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 586890 475174
rect 586270 474854 586890 474938
rect 586270 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 586890 474854
rect 586270 439174 586890 474618
rect 586270 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 586890 439174
rect 586270 438854 586890 438938
rect 586270 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 586890 438854
rect 586270 403174 586890 438618
rect 586270 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 586890 403174
rect 586270 402854 586890 402938
rect 586270 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 586890 402854
rect 586270 367174 586890 402618
rect 586270 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 586890 367174
rect 586270 366854 586890 366938
rect 586270 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 586890 366854
rect 586270 331174 586890 366618
rect 586270 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 586890 331174
rect 586270 330854 586890 330938
rect 586270 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 586890 330854
rect 586270 295174 586890 330618
rect 586270 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 586890 295174
rect 586270 294854 586890 294938
rect 586270 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 586890 294854
rect 586270 259174 586890 294618
rect 586270 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 586890 259174
rect 586270 258854 586890 258938
rect 586270 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 586890 258854
rect 586270 223174 586890 258618
rect 586270 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 586890 223174
rect 586270 222854 586890 222938
rect 586270 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 586890 222854
rect 586270 187174 586890 222618
rect 586270 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 586890 187174
rect 586270 186854 586890 186938
rect 586270 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 586890 186854
rect 586270 151174 586890 186618
rect 586270 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 586890 151174
rect 586270 150854 586890 150938
rect 586270 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 586890 150854
rect 586270 115174 586890 150618
rect 586270 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 586890 115174
rect 586270 114854 586890 114938
rect 586270 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 586890 114854
rect 586270 79174 586890 114618
rect 586270 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 586890 79174
rect 586270 78854 586890 78938
rect 586270 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 586890 78854
rect 586270 43174 586890 78618
rect 586270 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 586890 43174
rect 586270 42854 586890 42938
rect 586270 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 586890 42854
rect 586270 7174 586890 42618
rect 586270 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 586890 7174
rect 586270 6854 586890 6938
rect 586270 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 586890 6854
rect 581514 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 582134 -1306
rect 581514 -1626 582134 -1542
rect 581514 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 582134 -1626
rect 581514 -7654 582134 -1862
rect 586270 -1306 586890 6618
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 694894 587850 706202
rect 587230 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 587850 694894
rect 587230 694574 587850 694658
rect 587230 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 587850 694574
rect 587230 658894 587850 694338
rect 587230 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 587850 658894
rect 587230 658574 587850 658658
rect 587230 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 587850 658574
rect 587230 622894 587850 658338
rect 587230 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 587850 622894
rect 587230 622574 587850 622658
rect 587230 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 587850 622574
rect 587230 586894 587850 622338
rect 587230 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 587850 586894
rect 587230 586574 587850 586658
rect 587230 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 587850 586574
rect 587230 550894 587850 586338
rect 587230 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 587850 550894
rect 587230 550574 587850 550658
rect 587230 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 587850 550574
rect 587230 514894 587850 550338
rect 587230 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 587850 514894
rect 587230 514574 587850 514658
rect 587230 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 587850 514574
rect 587230 478894 587850 514338
rect 587230 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 587850 478894
rect 587230 478574 587850 478658
rect 587230 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 587850 478574
rect 587230 442894 587850 478338
rect 587230 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 587850 442894
rect 587230 442574 587850 442658
rect 587230 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 587850 442574
rect 587230 406894 587850 442338
rect 587230 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 587850 406894
rect 587230 406574 587850 406658
rect 587230 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 587850 406574
rect 587230 370894 587850 406338
rect 587230 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 587850 370894
rect 587230 370574 587850 370658
rect 587230 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 587850 370574
rect 587230 334894 587850 370338
rect 587230 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 587850 334894
rect 587230 334574 587850 334658
rect 587230 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 587850 334574
rect 587230 298894 587850 334338
rect 587230 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 587850 298894
rect 587230 298574 587850 298658
rect 587230 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 587850 298574
rect 587230 262894 587850 298338
rect 587230 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 587850 262894
rect 587230 262574 587850 262658
rect 587230 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 587850 262574
rect 587230 226894 587850 262338
rect 587230 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 587850 226894
rect 587230 226574 587850 226658
rect 587230 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 587850 226574
rect 587230 190894 587850 226338
rect 587230 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 587850 190894
rect 587230 190574 587850 190658
rect 587230 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 587850 190574
rect 587230 154894 587850 190338
rect 587230 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 587850 154894
rect 587230 154574 587850 154658
rect 587230 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 587850 154574
rect 587230 118894 587850 154338
rect 587230 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 587850 118894
rect 587230 118574 587850 118658
rect 587230 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 587850 118574
rect 587230 82894 587850 118338
rect 587230 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 587850 82894
rect 587230 82574 587850 82658
rect 587230 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 587850 82574
rect 587230 46894 587850 82338
rect 587230 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 587850 46894
rect 587230 46574 587850 46658
rect 587230 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 587850 46574
rect 587230 10894 587850 46338
rect 587230 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 587850 10894
rect 587230 10574 587850 10658
rect 587230 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 587850 10574
rect 587230 -2266 587850 10338
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 698614 588810 707162
rect 588190 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 588810 698614
rect 588190 698294 588810 698378
rect 588190 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 588810 698294
rect 588190 662614 588810 698058
rect 588190 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 588810 662614
rect 588190 662294 588810 662378
rect 588190 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 588810 662294
rect 588190 626614 588810 662058
rect 588190 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 588810 626614
rect 588190 626294 588810 626378
rect 588190 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 588810 626294
rect 588190 590614 588810 626058
rect 588190 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 588810 590614
rect 588190 590294 588810 590378
rect 588190 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 588810 590294
rect 588190 554614 588810 590058
rect 588190 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 588810 554614
rect 588190 554294 588810 554378
rect 588190 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 588810 554294
rect 588190 518614 588810 554058
rect 588190 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 588810 518614
rect 588190 518294 588810 518378
rect 588190 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 588810 518294
rect 588190 482614 588810 518058
rect 588190 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 588810 482614
rect 588190 482294 588810 482378
rect 588190 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 588810 482294
rect 588190 446614 588810 482058
rect 588190 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 588810 446614
rect 588190 446294 588810 446378
rect 588190 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 588810 446294
rect 588190 410614 588810 446058
rect 588190 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 588810 410614
rect 588190 410294 588810 410378
rect 588190 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 588810 410294
rect 588190 374614 588810 410058
rect 588190 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 588810 374614
rect 588190 374294 588810 374378
rect 588190 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 588810 374294
rect 588190 338614 588810 374058
rect 588190 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 588810 338614
rect 588190 338294 588810 338378
rect 588190 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 588810 338294
rect 588190 302614 588810 338058
rect 588190 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 588810 302614
rect 588190 302294 588810 302378
rect 588190 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 588810 302294
rect 588190 266614 588810 302058
rect 588190 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 588810 266614
rect 588190 266294 588810 266378
rect 588190 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 588810 266294
rect 588190 230614 588810 266058
rect 588190 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 588810 230614
rect 588190 230294 588810 230378
rect 588190 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 588810 230294
rect 588190 194614 588810 230058
rect 588190 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 588810 194614
rect 588190 194294 588810 194378
rect 588190 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 588810 194294
rect 588190 158614 588810 194058
rect 588190 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 588810 158614
rect 588190 158294 588810 158378
rect 588190 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 588810 158294
rect 588190 122614 588810 158058
rect 588190 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 588810 122614
rect 588190 122294 588810 122378
rect 588190 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 588810 122294
rect 588190 86614 588810 122058
rect 588190 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 588810 86614
rect 588190 86294 588810 86378
rect 588190 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 588810 86294
rect 588190 50614 588810 86058
rect 588190 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 588810 50614
rect 588190 50294 588810 50378
rect 588190 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 588810 50294
rect 588190 14614 588810 50058
rect 588190 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 588810 14614
rect 588190 14294 588810 14378
rect 588190 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 588810 14294
rect 588190 -3226 588810 14058
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 666334 589770 708122
rect 589150 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 589770 666334
rect 589150 666014 589770 666098
rect 589150 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 589770 666014
rect 589150 630334 589770 665778
rect 589150 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 589770 630334
rect 589150 630014 589770 630098
rect 589150 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 589770 630014
rect 589150 594334 589770 629778
rect 589150 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 589770 594334
rect 589150 594014 589770 594098
rect 589150 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 589770 594014
rect 589150 558334 589770 593778
rect 589150 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 589770 558334
rect 589150 558014 589770 558098
rect 589150 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 589770 558014
rect 589150 522334 589770 557778
rect 589150 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 589770 522334
rect 589150 522014 589770 522098
rect 589150 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 589770 522014
rect 589150 486334 589770 521778
rect 589150 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 589770 486334
rect 589150 486014 589770 486098
rect 589150 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 589770 486014
rect 589150 450334 589770 485778
rect 589150 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 589770 450334
rect 589150 450014 589770 450098
rect 589150 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 589770 450014
rect 589150 414334 589770 449778
rect 589150 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 589770 414334
rect 589150 414014 589770 414098
rect 589150 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 589770 414014
rect 589150 378334 589770 413778
rect 589150 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 589770 378334
rect 589150 378014 589770 378098
rect 589150 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 589770 378014
rect 589150 342334 589770 377778
rect 589150 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 589770 342334
rect 589150 342014 589770 342098
rect 589150 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 589770 342014
rect 589150 306334 589770 341778
rect 589150 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 589770 306334
rect 589150 306014 589770 306098
rect 589150 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 589770 306014
rect 589150 270334 589770 305778
rect 589150 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 589770 270334
rect 589150 270014 589770 270098
rect 589150 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 589770 270014
rect 589150 234334 589770 269778
rect 589150 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 589770 234334
rect 589150 234014 589770 234098
rect 589150 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 589770 234014
rect 589150 198334 589770 233778
rect 589150 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 589770 198334
rect 589150 198014 589770 198098
rect 589150 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 589770 198014
rect 589150 162334 589770 197778
rect 589150 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 589770 162334
rect 589150 162014 589770 162098
rect 589150 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 589770 162014
rect 589150 126334 589770 161778
rect 589150 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 589770 126334
rect 589150 126014 589770 126098
rect 589150 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 589770 126014
rect 589150 90334 589770 125778
rect 589150 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 589770 90334
rect 589150 90014 589770 90098
rect 589150 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 589770 90014
rect 589150 54334 589770 89778
rect 589150 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 589770 54334
rect 589150 54014 589770 54098
rect 589150 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 589770 54014
rect 589150 18334 589770 53778
rect 589150 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 589770 18334
rect 589150 18014 589770 18098
rect 589150 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 589770 18014
rect 589150 -4186 589770 17778
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 670054 590730 709082
rect 590110 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 590730 670054
rect 590110 669734 590730 669818
rect 590110 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 590730 669734
rect 590110 634054 590730 669498
rect 590110 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 590730 634054
rect 590110 633734 590730 633818
rect 590110 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 590730 633734
rect 590110 598054 590730 633498
rect 590110 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 590730 598054
rect 590110 597734 590730 597818
rect 590110 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 590730 597734
rect 590110 562054 590730 597498
rect 590110 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 590730 562054
rect 590110 561734 590730 561818
rect 590110 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 590730 561734
rect 590110 526054 590730 561498
rect 590110 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 590730 526054
rect 590110 525734 590730 525818
rect 590110 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 590730 525734
rect 590110 490054 590730 525498
rect 590110 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 590730 490054
rect 590110 489734 590730 489818
rect 590110 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 590730 489734
rect 590110 454054 590730 489498
rect 590110 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 590730 454054
rect 590110 453734 590730 453818
rect 590110 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 590730 453734
rect 590110 418054 590730 453498
rect 590110 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 590730 418054
rect 590110 417734 590730 417818
rect 590110 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 590730 417734
rect 590110 382054 590730 417498
rect 590110 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 590730 382054
rect 590110 381734 590730 381818
rect 590110 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 590730 381734
rect 590110 346054 590730 381498
rect 590110 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 590730 346054
rect 590110 345734 590730 345818
rect 590110 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 590730 345734
rect 590110 310054 590730 345498
rect 590110 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 590730 310054
rect 590110 309734 590730 309818
rect 590110 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 590730 309734
rect 590110 274054 590730 309498
rect 590110 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 590730 274054
rect 590110 273734 590730 273818
rect 590110 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 590730 273734
rect 590110 238054 590730 273498
rect 590110 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 590730 238054
rect 590110 237734 590730 237818
rect 590110 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 590730 237734
rect 590110 202054 590730 237498
rect 590110 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 590730 202054
rect 590110 201734 590730 201818
rect 590110 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 590730 201734
rect 590110 166054 590730 201498
rect 590110 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 590730 166054
rect 590110 165734 590730 165818
rect 590110 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 590730 165734
rect 590110 130054 590730 165498
rect 590110 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 590730 130054
rect 590110 129734 590730 129818
rect 590110 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 590730 129734
rect 590110 94054 590730 129498
rect 590110 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 590730 94054
rect 590110 93734 590730 93818
rect 590110 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 590730 93734
rect 590110 58054 590730 93498
rect 590110 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 590730 58054
rect 590110 57734 590730 57818
rect 590110 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 590730 57734
rect 590110 22054 590730 57498
rect 590110 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 590730 22054
rect 590110 21734 590730 21818
rect 590110 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 590730 21734
rect 590110 -5146 590730 21498
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 673774 591690 710042
rect 591070 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 591690 673774
rect 591070 673454 591690 673538
rect 591070 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 591690 673454
rect 591070 637774 591690 673218
rect 591070 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 591690 637774
rect 591070 637454 591690 637538
rect 591070 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 591690 637454
rect 591070 601774 591690 637218
rect 591070 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 591690 601774
rect 591070 601454 591690 601538
rect 591070 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 591690 601454
rect 591070 565774 591690 601218
rect 591070 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 591690 565774
rect 591070 565454 591690 565538
rect 591070 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 591690 565454
rect 591070 529774 591690 565218
rect 591070 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 591690 529774
rect 591070 529454 591690 529538
rect 591070 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 591690 529454
rect 591070 493774 591690 529218
rect 591070 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 591690 493774
rect 591070 493454 591690 493538
rect 591070 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 591690 493454
rect 591070 457774 591690 493218
rect 591070 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 591690 457774
rect 591070 457454 591690 457538
rect 591070 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 591690 457454
rect 591070 421774 591690 457218
rect 591070 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 591690 421774
rect 591070 421454 591690 421538
rect 591070 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 591690 421454
rect 591070 385774 591690 421218
rect 591070 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 591690 385774
rect 591070 385454 591690 385538
rect 591070 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 591690 385454
rect 591070 349774 591690 385218
rect 591070 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 591690 349774
rect 591070 349454 591690 349538
rect 591070 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 591690 349454
rect 591070 313774 591690 349218
rect 591070 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 591690 313774
rect 591070 313454 591690 313538
rect 591070 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 591690 313454
rect 591070 277774 591690 313218
rect 591070 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 591690 277774
rect 591070 277454 591690 277538
rect 591070 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 591690 277454
rect 591070 241774 591690 277218
rect 591070 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 591690 241774
rect 591070 241454 591690 241538
rect 591070 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 591690 241454
rect 591070 205774 591690 241218
rect 591070 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 591690 205774
rect 591070 205454 591690 205538
rect 591070 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 591690 205454
rect 591070 169774 591690 205218
rect 591070 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 591690 169774
rect 591070 169454 591690 169538
rect 591070 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 591690 169454
rect 591070 133774 591690 169218
rect 591070 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 591690 133774
rect 591070 133454 591690 133538
rect 591070 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 591690 133454
rect 591070 97774 591690 133218
rect 591070 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 591690 97774
rect 591070 97454 591690 97538
rect 591070 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 591690 97454
rect 591070 61774 591690 97218
rect 591070 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 591690 61774
rect 591070 61454 591690 61538
rect 591070 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 591690 61454
rect 591070 25774 591690 61218
rect 591070 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 591690 25774
rect 591070 25454 591690 25538
rect 591070 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 591690 25454
rect 591070 -6106 591690 25218
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 677494 592650 711002
rect 592030 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect 592030 677174 592650 677258
rect 592030 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect 592030 641494 592650 676938
rect 592030 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect 592030 641174 592650 641258
rect 592030 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect 592030 605494 592650 640938
rect 592030 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect 592030 605174 592650 605258
rect 592030 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect 592030 569494 592650 604938
rect 592030 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect 592030 569174 592650 569258
rect 592030 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect 592030 533494 592650 568938
rect 592030 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect 592030 533174 592650 533258
rect 592030 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect 592030 497494 592650 532938
rect 592030 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect 592030 497174 592650 497258
rect 592030 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect 592030 461494 592650 496938
rect 592030 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect 592030 461174 592650 461258
rect 592030 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect 592030 425494 592650 460938
rect 592030 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect 592030 425174 592650 425258
rect 592030 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect 592030 389494 592650 424938
rect 592030 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect 592030 389174 592650 389258
rect 592030 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect 592030 353494 592650 388938
rect 592030 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect 592030 353174 592650 353258
rect 592030 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect 592030 317494 592650 352938
rect 592030 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect 592030 317174 592650 317258
rect 592030 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect 592030 281494 592650 316938
rect 592030 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect 592030 281174 592650 281258
rect 592030 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect 592030 245494 592650 280938
rect 592030 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect 592030 245174 592650 245258
rect 592030 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect 592030 209494 592650 244938
rect 592030 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect 592030 209174 592650 209258
rect 592030 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect 592030 173494 592650 208938
rect 592030 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect 592030 173174 592650 173258
rect 592030 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect 592030 137494 592650 172938
rect 592030 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect 592030 137174 592650 137258
rect 592030 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect 592030 101494 592650 136938
rect 592030 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect 592030 101174 592650 101258
rect 592030 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect 592030 65494 592650 100938
rect 592030 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect 592030 65174 592650 65258
rect 592030 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect 592030 29494 592650 64938
rect 592030 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect 592030 29174 592650 29258
rect 592030 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect 592030 -7066 592650 28938
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 677258 -8458 677494
rect -8374 677258 -8138 677494
rect -8694 676938 -8458 677174
rect -8374 676938 -8138 677174
rect -8694 641258 -8458 641494
rect -8374 641258 -8138 641494
rect -8694 640938 -8458 641174
rect -8374 640938 -8138 641174
rect -8694 605258 -8458 605494
rect -8374 605258 -8138 605494
rect -8694 604938 -8458 605174
rect -8374 604938 -8138 605174
rect -8694 569258 -8458 569494
rect -8374 569258 -8138 569494
rect -8694 568938 -8458 569174
rect -8374 568938 -8138 569174
rect -8694 533258 -8458 533494
rect -8374 533258 -8138 533494
rect -8694 532938 -8458 533174
rect -8374 532938 -8138 533174
rect -8694 497258 -8458 497494
rect -8374 497258 -8138 497494
rect -8694 496938 -8458 497174
rect -8374 496938 -8138 497174
rect -8694 461258 -8458 461494
rect -8374 461258 -8138 461494
rect -8694 460938 -8458 461174
rect -8374 460938 -8138 461174
rect -8694 425258 -8458 425494
rect -8374 425258 -8138 425494
rect -8694 424938 -8458 425174
rect -8374 424938 -8138 425174
rect -8694 389258 -8458 389494
rect -8374 389258 -8138 389494
rect -8694 388938 -8458 389174
rect -8374 388938 -8138 389174
rect -8694 353258 -8458 353494
rect -8374 353258 -8138 353494
rect -8694 352938 -8458 353174
rect -8374 352938 -8138 353174
rect -8694 317258 -8458 317494
rect -8374 317258 -8138 317494
rect -8694 316938 -8458 317174
rect -8374 316938 -8138 317174
rect -8694 281258 -8458 281494
rect -8374 281258 -8138 281494
rect -8694 280938 -8458 281174
rect -8374 280938 -8138 281174
rect -8694 245258 -8458 245494
rect -8374 245258 -8138 245494
rect -8694 244938 -8458 245174
rect -8374 244938 -8138 245174
rect -8694 209258 -8458 209494
rect -8374 209258 -8138 209494
rect -8694 208938 -8458 209174
rect -8374 208938 -8138 209174
rect -8694 173258 -8458 173494
rect -8374 173258 -8138 173494
rect -8694 172938 -8458 173174
rect -8374 172938 -8138 173174
rect -8694 137258 -8458 137494
rect -8374 137258 -8138 137494
rect -8694 136938 -8458 137174
rect -8374 136938 -8138 137174
rect -8694 101258 -8458 101494
rect -8374 101258 -8138 101494
rect -8694 100938 -8458 101174
rect -8374 100938 -8138 101174
rect -8694 65258 -8458 65494
rect -8374 65258 -8138 65494
rect -8694 64938 -8458 65174
rect -8374 64938 -8138 65174
rect -8694 29258 -8458 29494
rect -8374 29258 -8138 29494
rect -8694 28938 -8458 29174
rect -8374 28938 -8138 29174
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 673538 -7498 673774
rect -7414 673538 -7178 673774
rect -7734 673218 -7498 673454
rect -7414 673218 -7178 673454
rect -7734 637538 -7498 637774
rect -7414 637538 -7178 637774
rect -7734 637218 -7498 637454
rect -7414 637218 -7178 637454
rect -7734 601538 -7498 601774
rect -7414 601538 -7178 601774
rect -7734 601218 -7498 601454
rect -7414 601218 -7178 601454
rect -7734 565538 -7498 565774
rect -7414 565538 -7178 565774
rect -7734 565218 -7498 565454
rect -7414 565218 -7178 565454
rect -7734 529538 -7498 529774
rect -7414 529538 -7178 529774
rect -7734 529218 -7498 529454
rect -7414 529218 -7178 529454
rect -7734 493538 -7498 493774
rect -7414 493538 -7178 493774
rect -7734 493218 -7498 493454
rect -7414 493218 -7178 493454
rect -7734 457538 -7498 457774
rect -7414 457538 -7178 457774
rect -7734 457218 -7498 457454
rect -7414 457218 -7178 457454
rect -7734 421538 -7498 421774
rect -7414 421538 -7178 421774
rect -7734 421218 -7498 421454
rect -7414 421218 -7178 421454
rect -7734 385538 -7498 385774
rect -7414 385538 -7178 385774
rect -7734 385218 -7498 385454
rect -7414 385218 -7178 385454
rect -7734 349538 -7498 349774
rect -7414 349538 -7178 349774
rect -7734 349218 -7498 349454
rect -7414 349218 -7178 349454
rect -7734 313538 -7498 313774
rect -7414 313538 -7178 313774
rect -7734 313218 -7498 313454
rect -7414 313218 -7178 313454
rect -7734 277538 -7498 277774
rect -7414 277538 -7178 277774
rect -7734 277218 -7498 277454
rect -7414 277218 -7178 277454
rect -7734 241538 -7498 241774
rect -7414 241538 -7178 241774
rect -7734 241218 -7498 241454
rect -7414 241218 -7178 241454
rect -7734 205538 -7498 205774
rect -7414 205538 -7178 205774
rect -7734 205218 -7498 205454
rect -7414 205218 -7178 205454
rect -7734 169538 -7498 169774
rect -7414 169538 -7178 169774
rect -7734 169218 -7498 169454
rect -7414 169218 -7178 169454
rect -7734 133538 -7498 133774
rect -7414 133538 -7178 133774
rect -7734 133218 -7498 133454
rect -7414 133218 -7178 133454
rect -7734 97538 -7498 97774
rect -7414 97538 -7178 97774
rect -7734 97218 -7498 97454
rect -7414 97218 -7178 97454
rect -7734 61538 -7498 61774
rect -7414 61538 -7178 61774
rect -7734 61218 -7498 61454
rect -7414 61218 -7178 61454
rect -7734 25538 -7498 25774
rect -7414 25538 -7178 25774
rect -7734 25218 -7498 25454
rect -7414 25218 -7178 25454
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 669818 -6538 670054
rect -6454 669818 -6218 670054
rect -6774 669498 -6538 669734
rect -6454 669498 -6218 669734
rect -6774 633818 -6538 634054
rect -6454 633818 -6218 634054
rect -6774 633498 -6538 633734
rect -6454 633498 -6218 633734
rect -6774 597818 -6538 598054
rect -6454 597818 -6218 598054
rect -6774 597498 -6538 597734
rect -6454 597498 -6218 597734
rect -6774 561818 -6538 562054
rect -6454 561818 -6218 562054
rect -6774 561498 -6538 561734
rect -6454 561498 -6218 561734
rect -6774 525818 -6538 526054
rect -6454 525818 -6218 526054
rect -6774 525498 -6538 525734
rect -6454 525498 -6218 525734
rect -6774 489818 -6538 490054
rect -6454 489818 -6218 490054
rect -6774 489498 -6538 489734
rect -6454 489498 -6218 489734
rect -6774 453818 -6538 454054
rect -6454 453818 -6218 454054
rect -6774 453498 -6538 453734
rect -6454 453498 -6218 453734
rect -6774 417818 -6538 418054
rect -6454 417818 -6218 418054
rect -6774 417498 -6538 417734
rect -6454 417498 -6218 417734
rect -6774 381818 -6538 382054
rect -6454 381818 -6218 382054
rect -6774 381498 -6538 381734
rect -6454 381498 -6218 381734
rect -6774 345818 -6538 346054
rect -6454 345818 -6218 346054
rect -6774 345498 -6538 345734
rect -6454 345498 -6218 345734
rect -6774 309818 -6538 310054
rect -6454 309818 -6218 310054
rect -6774 309498 -6538 309734
rect -6454 309498 -6218 309734
rect -6774 273818 -6538 274054
rect -6454 273818 -6218 274054
rect -6774 273498 -6538 273734
rect -6454 273498 -6218 273734
rect -6774 237818 -6538 238054
rect -6454 237818 -6218 238054
rect -6774 237498 -6538 237734
rect -6454 237498 -6218 237734
rect -6774 201818 -6538 202054
rect -6454 201818 -6218 202054
rect -6774 201498 -6538 201734
rect -6454 201498 -6218 201734
rect -6774 165818 -6538 166054
rect -6454 165818 -6218 166054
rect -6774 165498 -6538 165734
rect -6454 165498 -6218 165734
rect -6774 129818 -6538 130054
rect -6454 129818 -6218 130054
rect -6774 129498 -6538 129734
rect -6454 129498 -6218 129734
rect -6774 93818 -6538 94054
rect -6454 93818 -6218 94054
rect -6774 93498 -6538 93734
rect -6454 93498 -6218 93734
rect -6774 57818 -6538 58054
rect -6454 57818 -6218 58054
rect -6774 57498 -6538 57734
rect -6454 57498 -6218 57734
rect -6774 21818 -6538 22054
rect -6454 21818 -6218 22054
rect -6774 21498 -6538 21734
rect -6454 21498 -6218 21734
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 666098 -5578 666334
rect -5494 666098 -5258 666334
rect -5814 665778 -5578 666014
rect -5494 665778 -5258 666014
rect -5814 630098 -5578 630334
rect -5494 630098 -5258 630334
rect -5814 629778 -5578 630014
rect -5494 629778 -5258 630014
rect -5814 594098 -5578 594334
rect -5494 594098 -5258 594334
rect -5814 593778 -5578 594014
rect -5494 593778 -5258 594014
rect -5814 558098 -5578 558334
rect -5494 558098 -5258 558334
rect -5814 557778 -5578 558014
rect -5494 557778 -5258 558014
rect -5814 522098 -5578 522334
rect -5494 522098 -5258 522334
rect -5814 521778 -5578 522014
rect -5494 521778 -5258 522014
rect -5814 486098 -5578 486334
rect -5494 486098 -5258 486334
rect -5814 485778 -5578 486014
rect -5494 485778 -5258 486014
rect -5814 450098 -5578 450334
rect -5494 450098 -5258 450334
rect -5814 449778 -5578 450014
rect -5494 449778 -5258 450014
rect -5814 414098 -5578 414334
rect -5494 414098 -5258 414334
rect -5814 413778 -5578 414014
rect -5494 413778 -5258 414014
rect -5814 378098 -5578 378334
rect -5494 378098 -5258 378334
rect -5814 377778 -5578 378014
rect -5494 377778 -5258 378014
rect -5814 342098 -5578 342334
rect -5494 342098 -5258 342334
rect -5814 341778 -5578 342014
rect -5494 341778 -5258 342014
rect -5814 306098 -5578 306334
rect -5494 306098 -5258 306334
rect -5814 305778 -5578 306014
rect -5494 305778 -5258 306014
rect -5814 270098 -5578 270334
rect -5494 270098 -5258 270334
rect -5814 269778 -5578 270014
rect -5494 269778 -5258 270014
rect -5814 234098 -5578 234334
rect -5494 234098 -5258 234334
rect -5814 233778 -5578 234014
rect -5494 233778 -5258 234014
rect -5814 198098 -5578 198334
rect -5494 198098 -5258 198334
rect -5814 197778 -5578 198014
rect -5494 197778 -5258 198014
rect -5814 162098 -5578 162334
rect -5494 162098 -5258 162334
rect -5814 161778 -5578 162014
rect -5494 161778 -5258 162014
rect -5814 126098 -5578 126334
rect -5494 126098 -5258 126334
rect -5814 125778 -5578 126014
rect -5494 125778 -5258 126014
rect -5814 90098 -5578 90334
rect -5494 90098 -5258 90334
rect -5814 89778 -5578 90014
rect -5494 89778 -5258 90014
rect -5814 54098 -5578 54334
rect -5494 54098 -5258 54334
rect -5814 53778 -5578 54014
rect -5494 53778 -5258 54014
rect -5814 18098 -5578 18334
rect -5494 18098 -5258 18334
rect -5814 17778 -5578 18014
rect -5494 17778 -5258 18014
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 698378 -4618 698614
rect -4534 698378 -4298 698614
rect -4854 698058 -4618 698294
rect -4534 698058 -4298 698294
rect -4854 662378 -4618 662614
rect -4534 662378 -4298 662614
rect -4854 662058 -4618 662294
rect -4534 662058 -4298 662294
rect -4854 626378 -4618 626614
rect -4534 626378 -4298 626614
rect -4854 626058 -4618 626294
rect -4534 626058 -4298 626294
rect -4854 590378 -4618 590614
rect -4534 590378 -4298 590614
rect -4854 590058 -4618 590294
rect -4534 590058 -4298 590294
rect -4854 554378 -4618 554614
rect -4534 554378 -4298 554614
rect -4854 554058 -4618 554294
rect -4534 554058 -4298 554294
rect -4854 518378 -4618 518614
rect -4534 518378 -4298 518614
rect -4854 518058 -4618 518294
rect -4534 518058 -4298 518294
rect -4854 482378 -4618 482614
rect -4534 482378 -4298 482614
rect -4854 482058 -4618 482294
rect -4534 482058 -4298 482294
rect -4854 446378 -4618 446614
rect -4534 446378 -4298 446614
rect -4854 446058 -4618 446294
rect -4534 446058 -4298 446294
rect -4854 410378 -4618 410614
rect -4534 410378 -4298 410614
rect -4854 410058 -4618 410294
rect -4534 410058 -4298 410294
rect -4854 374378 -4618 374614
rect -4534 374378 -4298 374614
rect -4854 374058 -4618 374294
rect -4534 374058 -4298 374294
rect -4854 338378 -4618 338614
rect -4534 338378 -4298 338614
rect -4854 338058 -4618 338294
rect -4534 338058 -4298 338294
rect -4854 302378 -4618 302614
rect -4534 302378 -4298 302614
rect -4854 302058 -4618 302294
rect -4534 302058 -4298 302294
rect -4854 266378 -4618 266614
rect -4534 266378 -4298 266614
rect -4854 266058 -4618 266294
rect -4534 266058 -4298 266294
rect -4854 230378 -4618 230614
rect -4534 230378 -4298 230614
rect -4854 230058 -4618 230294
rect -4534 230058 -4298 230294
rect -4854 194378 -4618 194614
rect -4534 194378 -4298 194614
rect -4854 194058 -4618 194294
rect -4534 194058 -4298 194294
rect -4854 158378 -4618 158614
rect -4534 158378 -4298 158614
rect -4854 158058 -4618 158294
rect -4534 158058 -4298 158294
rect -4854 122378 -4618 122614
rect -4534 122378 -4298 122614
rect -4854 122058 -4618 122294
rect -4534 122058 -4298 122294
rect -4854 86378 -4618 86614
rect -4534 86378 -4298 86614
rect -4854 86058 -4618 86294
rect -4534 86058 -4298 86294
rect -4854 50378 -4618 50614
rect -4534 50378 -4298 50614
rect -4854 50058 -4618 50294
rect -4534 50058 -4298 50294
rect -4854 14378 -4618 14614
rect -4534 14378 -4298 14614
rect -4854 14058 -4618 14294
rect -4534 14058 -4298 14294
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 694658 -3658 694894
rect -3574 694658 -3338 694894
rect -3894 694338 -3658 694574
rect -3574 694338 -3338 694574
rect -3894 658658 -3658 658894
rect -3574 658658 -3338 658894
rect -3894 658338 -3658 658574
rect -3574 658338 -3338 658574
rect -3894 622658 -3658 622894
rect -3574 622658 -3338 622894
rect -3894 622338 -3658 622574
rect -3574 622338 -3338 622574
rect -3894 586658 -3658 586894
rect -3574 586658 -3338 586894
rect -3894 586338 -3658 586574
rect -3574 586338 -3338 586574
rect -3894 550658 -3658 550894
rect -3574 550658 -3338 550894
rect -3894 550338 -3658 550574
rect -3574 550338 -3338 550574
rect -3894 514658 -3658 514894
rect -3574 514658 -3338 514894
rect -3894 514338 -3658 514574
rect -3574 514338 -3338 514574
rect -3894 478658 -3658 478894
rect -3574 478658 -3338 478894
rect -3894 478338 -3658 478574
rect -3574 478338 -3338 478574
rect -3894 442658 -3658 442894
rect -3574 442658 -3338 442894
rect -3894 442338 -3658 442574
rect -3574 442338 -3338 442574
rect -3894 406658 -3658 406894
rect -3574 406658 -3338 406894
rect -3894 406338 -3658 406574
rect -3574 406338 -3338 406574
rect -3894 370658 -3658 370894
rect -3574 370658 -3338 370894
rect -3894 370338 -3658 370574
rect -3574 370338 -3338 370574
rect -3894 334658 -3658 334894
rect -3574 334658 -3338 334894
rect -3894 334338 -3658 334574
rect -3574 334338 -3338 334574
rect -3894 298658 -3658 298894
rect -3574 298658 -3338 298894
rect -3894 298338 -3658 298574
rect -3574 298338 -3338 298574
rect -3894 262658 -3658 262894
rect -3574 262658 -3338 262894
rect -3894 262338 -3658 262574
rect -3574 262338 -3338 262574
rect -3894 226658 -3658 226894
rect -3574 226658 -3338 226894
rect -3894 226338 -3658 226574
rect -3574 226338 -3338 226574
rect -3894 190658 -3658 190894
rect -3574 190658 -3338 190894
rect -3894 190338 -3658 190574
rect -3574 190338 -3338 190574
rect -3894 154658 -3658 154894
rect -3574 154658 -3338 154894
rect -3894 154338 -3658 154574
rect -3574 154338 -3338 154574
rect -3894 118658 -3658 118894
rect -3574 118658 -3338 118894
rect -3894 118338 -3658 118574
rect -3574 118338 -3338 118574
rect -3894 82658 -3658 82894
rect -3574 82658 -3338 82894
rect -3894 82338 -3658 82574
rect -3574 82338 -3338 82574
rect -3894 46658 -3658 46894
rect -3574 46658 -3338 46894
rect -3894 46338 -3658 46574
rect -3574 46338 -3338 46574
rect -3894 10658 -3658 10894
rect -3574 10658 -3338 10894
rect -3894 10338 -3658 10574
rect -3574 10338 -3338 10574
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 690938 -2698 691174
rect -2614 690938 -2378 691174
rect -2934 690618 -2698 690854
rect -2614 690618 -2378 690854
rect -2934 654938 -2698 655174
rect -2614 654938 -2378 655174
rect -2934 654618 -2698 654854
rect -2614 654618 -2378 654854
rect -2934 618938 -2698 619174
rect -2614 618938 -2378 619174
rect -2934 618618 -2698 618854
rect -2614 618618 -2378 618854
rect -2934 582938 -2698 583174
rect -2614 582938 -2378 583174
rect -2934 582618 -2698 582854
rect -2614 582618 -2378 582854
rect -2934 546938 -2698 547174
rect -2614 546938 -2378 547174
rect -2934 546618 -2698 546854
rect -2614 546618 -2378 546854
rect -2934 510938 -2698 511174
rect -2614 510938 -2378 511174
rect -2934 510618 -2698 510854
rect -2614 510618 -2378 510854
rect -2934 474938 -2698 475174
rect -2614 474938 -2378 475174
rect -2934 474618 -2698 474854
rect -2614 474618 -2378 474854
rect -2934 438938 -2698 439174
rect -2614 438938 -2378 439174
rect -2934 438618 -2698 438854
rect -2614 438618 -2378 438854
rect -2934 402938 -2698 403174
rect -2614 402938 -2378 403174
rect -2934 402618 -2698 402854
rect -2614 402618 -2378 402854
rect -2934 366938 -2698 367174
rect -2614 366938 -2378 367174
rect -2934 366618 -2698 366854
rect -2614 366618 -2378 366854
rect -2934 330938 -2698 331174
rect -2614 330938 -2378 331174
rect -2934 330618 -2698 330854
rect -2614 330618 -2378 330854
rect -2934 294938 -2698 295174
rect -2614 294938 -2378 295174
rect -2934 294618 -2698 294854
rect -2614 294618 -2378 294854
rect -2934 258938 -2698 259174
rect -2614 258938 -2378 259174
rect -2934 258618 -2698 258854
rect -2614 258618 -2378 258854
rect -2934 222938 -2698 223174
rect -2614 222938 -2378 223174
rect -2934 222618 -2698 222854
rect -2614 222618 -2378 222854
rect -2934 186938 -2698 187174
rect -2614 186938 -2378 187174
rect -2934 186618 -2698 186854
rect -2614 186618 -2378 186854
rect -2934 150938 -2698 151174
rect -2614 150938 -2378 151174
rect -2934 150618 -2698 150854
rect -2614 150618 -2378 150854
rect -2934 114938 -2698 115174
rect -2614 114938 -2378 115174
rect -2934 114618 -2698 114854
rect -2614 114618 -2378 114854
rect -2934 78938 -2698 79174
rect -2614 78938 -2378 79174
rect -2934 78618 -2698 78854
rect -2614 78618 -2378 78854
rect -2934 42938 -2698 43174
rect -2614 42938 -2378 43174
rect -2934 42618 -2698 42854
rect -2614 42618 -2378 42854
rect -2934 6938 -2698 7174
rect -2614 6938 -2378 7174
rect -2934 6618 -2698 6854
rect -2614 6618 -2378 6854
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 5546 705562 5782 705798
rect 5866 705562 6102 705798
rect 5546 705242 5782 705478
rect 5866 705242 6102 705478
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect 5546 -1542 5782 -1306
rect 5866 -1542 6102 -1306
rect 5546 -1862 5782 -1626
rect 5866 -1862 6102 -1626
rect 9266 706522 9502 706758
rect 9586 706522 9822 706758
rect 9266 706202 9502 706438
rect 9586 706202 9822 706438
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect 9266 -2502 9502 -2266
rect 9586 -2502 9822 -2266
rect 9266 -2822 9502 -2586
rect 9586 -2822 9822 -2586
rect 12986 707482 13222 707718
rect 13306 707482 13542 707718
rect 12986 707162 13222 707398
rect 13306 707162 13542 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect 12986 -3462 13222 -3226
rect 13306 -3462 13542 -3226
rect 12986 -3782 13222 -3546
rect 13306 -3782 13542 -3546
rect 16706 708442 16942 708678
rect 17026 708442 17262 708678
rect 16706 708122 16942 708358
rect 17026 708122 17262 708358
rect 16706 666098 16942 666334
rect 17026 666098 17262 666334
rect 16706 665778 16942 666014
rect 17026 665778 17262 666014
rect 16706 630098 16942 630334
rect 17026 630098 17262 630334
rect 16706 629778 16942 630014
rect 17026 629778 17262 630014
rect 16706 594098 16942 594334
rect 17026 594098 17262 594334
rect 16706 593778 16942 594014
rect 17026 593778 17262 594014
rect 16706 558098 16942 558334
rect 17026 558098 17262 558334
rect 16706 557778 16942 558014
rect 17026 557778 17262 558014
rect 16706 522098 16942 522334
rect 17026 522098 17262 522334
rect 16706 521778 16942 522014
rect 17026 521778 17262 522014
rect 16706 486098 16942 486334
rect 17026 486098 17262 486334
rect 16706 485778 16942 486014
rect 17026 485778 17262 486014
rect 16706 450098 16942 450334
rect 17026 450098 17262 450334
rect 16706 449778 16942 450014
rect 17026 449778 17262 450014
rect 16706 414098 16942 414334
rect 17026 414098 17262 414334
rect 16706 413778 16942 414014
rect 17026 413778 17262 414014
rect 16706 378098 16942 378334
rect 17026 378098 17262 378334
rect 16706 377778 16942 378014
rect 17026 377778 17262 378014
rect 16706 342098 16942 342334
rect 17026 342098 17262 342334
rect 16706 341778 16942 342014
rect 17026 341778 17262 342014
rect 16706 306098 16942 306334
rect 17026 306098 17262 306334
rect 16706 305778 16942 306014
rect 17026 305778 17262 306014
rect 16706 270098 16942 270334
rect 17026 270098 17262 270334
rect 16706 269778 16942 270014
rect 17026 269778 17262 270014
rect 16706 234098 16942 234334
rect 17026 234098 17262 234334
rect 16706 233778 16942 234014
rect 17026 233778 17262 234014
rect 16706 198098 16942 198334
rect 17026 198098 17262 198334
rect 16706 197778 16942 198014
rect 17026 197778 17262 198014
rect 16706 162098 16942 162334
rect 17026 162098 17262 162334
rect 16706 161778 16942 162014
rect 17026 161778 17262 162014
rect 16706 126098 16942 126334
rect 17026 126098 17262 126334
rect 16706 125778 16942 126014
rect 17026 125778 17262 126014
rect 16706 90098 16942 90334
rect 17026 90098 17262 90334
rect 16706 89778 16942 90014
rect 17026 89778 17262 90014
rect 16706 54098 16942 54334
rect 17026 54098 17262 54334
rect 16706 53778 16942 54014
rect 17026 53778 17262 54014
rect 16706 18098 16942 18334
rect 17026 18098 17262 18334
rect 16706 17778 16942 18014
rect 17026 17778 17262 18014
rect 16706 -4422 16942 -4186
rect 17026 -4422 17262 -4186
rect 16706 -4742 16942 -4506
rect 17026 -4742 17262 -4506
rect 20426 709402 20662 709638
rect 20746 709402 20982 709638
rect 20426 709082 20662 709318
rect 20746 709082 20982 709318
rect 20426 669818 20662 670054
rect 20746 669818 20982 670054
rect 20426 669498 20662 669734
rect 20746 669498 20982 669734
rect 27866 711322 28102 711558
rect 28186 711322 28422 711558
rect 27866 711002 28102 711238
rect 28186 711002 28422 711238
rect 27866 677258 28102 677494
rect 28186 677258 28422 677494
rect 27866 676938 28102 677174
rect 28186 676938 28422 677174
rect 24250 651218 24486 651454
rect 24250 650898 24486 651134
rect 20426 633818 20662 634054
rect 20746 633818 20982 634054
rect 20426 633498 20662 633734
rect 20746 633498 20982 633734
rect 27866 641258 28102 641494
rect 28186 641258 28422 641494
rect 27866 640938 28102 641174
rect 28186 640938 28422 641174
rect 24250 615218 24486 615454
rect 24250 614898 24486 615134
rect 20426 597818 20662 598054
rect 20746 597818 20982 598054
rect 20426 597498 20662 597734
rect 20746 597498 20982 597734
rect 27866 605258 28102 605494
rect 28186 605258 28422 605494
rect 27866 604938 28102 605174
rect 28186 604938 28422 605174
rect 24250 579218 24486 579454
rect 24250 578898 24486 579134
rect 20426 561818 20662 562054
rect 20746 561818 20982 562054
rect 20426 561498 20662 561734
rect 20746 561498 20982 561734
rect 27866 569258 28102 569494
rect 28186 569258 28422 569494
rect 27866 568938 28102 569174
rect 28186 568938 28422 569174
rect 24250 543218 24486 543454
rect 24250 542898 24486 543134
rect 20426 525818 20662 526054
rect 20746 525818 20982 526054
rect 20426 525498 20662 525734
rect 20746 525498 20982 525734
rect 27866 533258 28102 533494
rect 28186 533258 28422 533494
rect 27866 532938 28102 533174
rect 28186 532938 28422 533174
rect 24250 507218 24486 507454
rect 24250 506898 24486 507134
rect 20426 489818 20662 490054
rect 20746 489818 20982 490054
rect 20426 489498 20662 489734
rect 20746 489498 20982 489734
rect 27866 497258 28102 497494
rect 28186 497258 28422 497494
rect 27866 496938 28102 497174
rect 28186 496938 28422 497174
rect 24250 471218 24486 471454
rect 24250 470898 24486 471134
rect 20426 453818 20662 454054
rect 20746 453818 20982 454054
rect 20426 453498 20662 453734
rect 20746 453498 20982 453734
rect 27866 461258 28102 461494
rect 28186 461258 28422 461494
rect 27866 460938 28102 461174
rect 28186 460938 28422 461174
rect 24250 435218 24486 435454
rect 24250 434898 24486 435134
rect 20426 417818 20662 418054
rect 20746 417818 20982 418054
rect 20426 417498 20662 417734
rect 20746 417498 20982 417734
rect 27866 425258 28102 425494
rect 28186 425258 28422 425494
rect 27866 424938 28102 425174
rect 28186 424938 28422 425174
rect 24250 399218 24486 399454
rect 24250 398898 24486 399134
rect 20426 381818 20662 382054
rect 20746 381818 20982 382054
rect 20426 381498 20662 381734
rect 20746 381498 20982 381734
rect 27866 389258 28102 389494
rect 28186 389258 28422 389494
rect 27866 388938 28102 389174
rect 28186 388938 28422 389174
rect 24250 363218 24486 363454
rect 24250 362898 24486 363134
rect 20426 345818 20662 346054
rect 20746 345818 20982 346054
rect 20426 345498 20662 345734
rect 20746 345498 20982 345734
rect 27866 353258 28102 353494
rect 28186 353258 28422 353494
rect 27866 352938 28102 353174
rect 28186 352938 28422 353174
rect 24250 327218 24486 327454
rect 24250 326898 24486 327134
rect 20426 309818 20662 310054
rect 20746 309818 20982 310054
rect 20426 309498 20662 309734
rect 20746 309498 20982 309734
rect 27866 317258 28102 317494
rect 28186 317258 28422 317494
rect 27866 316938 28102 317174
rect 28186 316938 28422 317174
rect 24250 291218 24486 291454
rect 24250 290898 24486 291134
rect 20426 273818 20662 274054
rect 20746 273818 20982 274054
rect 20426 273498 20662 273734
rect 20746 273498 20982 273734
rect 27866 281258 28102 281494
rect 28186 281258 28422 281494
rect 27866 280938 28102 281174
rect 28186 280938 28422 281174
rect 24250 255218 24486 255454
rect 24250 254898 24486 255134
rect 20426 237818 20662 238054
rect 20746 237818 20982 238054
rect 20426 237498 20662 237734
rect 20746 237498 20982 237734
rect 27866 245258 28102 245494
rect 28186 245258 28422 245494
rect 27866 244938 28102 245174
rect 28186 244938 28422 245174
rect 24250 219218 24486 219454
rect 24250 218898 24486 219134
rect 20426 201818 20662 202054
rect 20746 201818 20982 202054
rect 20426 201498 20662 201734
rect 20746 201498 20982 201734
rect 27866 209258 28102 209494
rect 28186 209258 28422 209494
rect 27866 208938 28102 209174
rect 28186 208938 28422 209174
rect 24250 183218 24486 183454
rect 24250 182898 24486 183134
rect 20426 165818 20662 166054
rect 20746 165818 20982 166054
rect 20426 165498 20662 165734
rect 20746 165498 20982 165734
rect 27866 173258 28102 173494
rect 28186 173258 28422 173494
rect 27866 172938 28102 173174
rect 28186 172938 28422 173174
rect 24250 147218 24486 147454
rect 24250 146898 24486 147134
rect 20426 129818 20662 130054
rect 20746 129818 20982 130054
rect 20426 129498 20662 129734
rect 20746 129498 20982 129734
rect 27866 137258 28102 137494
rect 28186 137258 28422 137494
rect 27866 136938 28102 137174
rect 28186 136938 28422 137174
rect 24250 111218 24486 111454
rect 24250 110898 24486 111134
rect 20426 93818 20662 94054
rect 20746 93818 20982 94054
rect 20426 93498 20662 93734
rect 20746 93498 20982 93734
rect 27866 101258 28102 101494
rect 28186 101258 28422 101494
rect 27866 100938 28102 101174
rect 28186 100938 28422 101174
rect 24250 75218 24486 75454
rect 24250 74898 24486 75134
rect 27866 65258 28102 65494
rect 28186 65258 28422 65494
rect 27866 64938 28102 65174
rect 28186 64938 28422 65174
rect 20426 57818 20662 58054
rect 20746 57818 20982 58054
rect 20426 57498 20662 57734
rect 20746 57498 20982 57734
rect 20426 21818 20662 22054
rect 20746 21818 20982 22054
rect 20426 21498 20662 21734
rect 20746 21498 20982 21734
rect 20426 -5382 20662 -5146
rect 20746 -5382 20982 -5146
rect 20426 -5702 20662 -5466
rect 20746 -5702 20982 -5466
rect 24146 25538 24382 25774
rect 24466 25538 24702 25774
rect 24146 25218 24382 25454
rect 24466 25218 24702 25454
rect 24146 -6342 24382 -6106
rect 24466 -6342 24702 -6106
rect 24146 -6662 24382 -6426
rect 24466 -6662 24702 -6426
rect 27866 29258 28102 29494
rect 28186 29258 28422 29494
rect 27866 28938 28102 29174
rect 28186 28938 28422 29174
rect 27866 -7302 28102 -7066
rect 28186 -7302 28422 -7066
rect 27866 -7622 28102 -7386
rect 28186 -7622 28422 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 41546 705562 41782 705798
rect 41866 705562 42102 705798
rect 41546 705242 41782 705478
rect 41866 705242 42102 705478
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 39610 654938 39846 655174
rect 39610 654618 39846 654854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 39610 618938 39846 619174
rect 39610 618618 39846 618854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 39610 582938 39846 583174
rect 39610 582618 39846 582854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 39610 546938 39846 547174
rect 39610 546618 39846 546854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 39610 510938 39846 511174
rect 39610 510618 39846 510854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 39610 474938 39846 475174
rect 39610 474618 39846 474854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 39610 438938 39846 439174
rect 39610 438618 39846 438854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 39610 402938 39846 403174
rect 39610 402618 39846 402854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 39610 366938 39846 367174
rect 39610 366618 39846 366854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 39610 330938 39846 331174
rect 39610 330618 39846 330854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 39610 294938 39846 295174
rect 39610 294618 39846 294854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 39610 258938 39846 259174
rect 39610 258618 39846 258854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 39610 222938 39846 223174
rect 39610 222618 39846 222854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 39610 186938 39846 187174
rect 39610 186618 39846 186854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 39610 150938 39846 151174
rect 39610 150618 39846 150854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 39610 114938 39846 115174
rect 39610 114618 39846 114854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 39610 78938 39846 79174
rect 39610 78618 39846 78854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -1542 41782 -1306
rect 41866 -1542 42102 -1306
rect 41546 -1862 41782 -1626
rect 41866 -1862 42102 -1626
rect 45266 706522 45502 706758
rect 45586 706522 45822 706758
rect 45266 706202 45502 706438
rect 45586 706202 45822 706438
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -2502 45502 -2266
rect 45586 -2502 45822 -2266
rect 45266 -2822 45502 -2586
rect 45586 -2822 45822 -2586
rect 48986 707482 49222 707718
rect 49306 707482 49542 707718
rect 48986 707162 49222 707398
rect 49306 707162 49542 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 77546 705562 77782 705798
rect 77866 705562 78102 705798
rect 77546 705242 77782 705478
rect 77866 705242 78102 705478
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 81266 706522 81502 706758
rect 81586 706522 81822 706758
rect 81266 706202 81502 706438
rect 81586 706202 81822 706438
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 84986 707482 85222 707718
rect 85306 707482 85542 707718
rect 84986 707162 85222 707398
rect 85306 707162 85542 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 113546 705562 113782 705798
rect 113866 705562 114102 705798
rect 113546 705242 113782 705478
rect 113866 705242 114102 705478
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 117266 706522 117502 706758
rect 117586 706522 117822 706758
rect 117266 706202 117502 706438
rect 117586 706202 117822 706438
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 120986 707482 121222 707718
rect 121306 707482 121542 707718
rect 120986 707162 121222 707398
rect 121306 707162 121542 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 149546 705562 149782 705798
rect 149866 705562 150102 705798
rect 149546 705242 149782 705478
rect 149866 705242 150102 705478
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 153266 706522 153502 706758
rect 153586 706522 153822 706758
rect 153266 706202 153502 706438
rect 153586 706202 153822 706438
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 156986 707482 157222 707718
rect 157306 707482 157542 707718
rect 156986 707162 157222 707398
rect 157306 707162 157542 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 185546 705562 185782 705798
rect 185866 705562 186102 705798
rect 185546 705242 185782 705478
rect 185866 705242 186102 705478
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 189266 706522 189502 706758
rect 189586 706522 189822 706758
rect 189266 706202 189502 706438
rect 189586 706202 189822 706438
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 192986 707482 193222 707718
rect 193306 707482 193542 707718
rect 192986 707162 193222 707398
rect 193306 707162 193542 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 221546 705562 221782 705798
rect 221866 705562 222102 705798
rect 221546 705242 221782 705478
rect 221866 705242 222102 705478
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 225266 706522 225502 706758
rect 225586 706522 225822 706758
rect 225266 706202 225502 706438
rect 225586 706202 225822 706438
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 228986 707482 229222 707718
rect 229306 707482 229542 707718
rect 228986 707162 229222 707398
rect 229306 707162 229542 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 257546 705562 257782 705798
rect 257866 705562 258102 705798
rect 257546 705242 257782 705478
rect 257866 705242 258102 705478
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 261266 706522 261502 706758
rect 261586 706522 261822 706758
rect 261266 706202 261502 706438
rect 261586 706202 261822 706438
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 264986 707482 265222 707718
rect 265306 707482 265542 707718
rect 264986 707162 265222 707398
rect 265306 707162 265542 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 293546 705562 293782 705798
rect 293866 705562 294102 705798
rect 293546 705242 293782 705478
rect 293866 705242 294102 705478
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 297266 706522 297502 706758
rect 297586 706522 297822 706758
rect 297266 706202 297502 706438
rect 297586 706202 297822 706438
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 300986 707482 301222 707718
rect 301306 707482 301542 707718
rect 300986 707162 301222 707398
rect 301306 707162 301542 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 329546 705562 329782 705798
rect 329866 705562 330102 705798
rect 329546 705242 329782 705478
rect 329866 705242 330102 705478
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 333266 706522 333502 706758
rect 333586 706522 333822 706758
rect 333266 706202 333502 706438
rect 333586 706202 333822 706438
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 336986 707482 337222 707718
rect 337306 707482 337542 707718
rect 336986 707162 337222 707398
rect 337306 707162 337542 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 344426 709402 344662 709638
rect 344746 709402 344982 709638
rect 344426 709082 344662 709318
rect 344746 709082 344982 709318
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 344426 669818 344662 670054
rect 344746 669818 344982 670054
rect 344426 669498 344662 669734
rect 344746 669498 344982 669734
rect 70330 654938 70566 655174
rect 70330 654618 70566 654854
rect 101050 654938 101286 655174
rect 101050 654618 101286 654854
rect 131770 654938 132006 655174
rect 131770 654618 132006 654854
rect 162490 654938 162726 655174
rect 162490 654618 162726 654854
rect 193210 654938 193446 655174
rect 193210 654618 193446 654854
rect 223930 654938 224166 655174
rect 223930 654618 224166 654854
rect 254650 654938 254886 655174
rect 254650 654618 254886 654854
rect 285370 654938 285606 655174
rect 285370 654618 285606 654854
rect 316090 654938 316326 655174
rect 316090 654618 316326 654854
rect 54970 651218 55206 651454
rect 54970 650898 55206 651134
rect 85690 651218 85926 651454
rect 85690 650898 85926 651134
rect 116410 651218 116646 651454
rect 116410 650898 116646 651134
rect 147130 651218 147366 651454
rect 147130 650898 147366 651134
rect 177850 651218 178086 651454
rect 177850 650898 178086 651134
rect 208570 651218 208806 651454
rect 208570 650898 208806 651134
rect 239290 651218 239526 651454
rect 239290 650898 239526 651134
rect 270010 651218 270246 651454
rect 270010 650898 270246 651134
rect 300730 651218 300966 651454
rect 300730 650898 300966 651134
rect 331450 651218 331686 651454
rect 331450 650898 331686 651134
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 348146 710362 348382 710598
rect 348466 710362 348702 710598
rect 348146 710042 348382 710278
rect 348466 710042 348702 710278
rect 348146 673538 348382 673774
rect 348466 673538 348702 673774
rect 348146 673218 348382 673454
rect 348466 673218 348702 673454
rect 346810 654938 347046 655174
rect 346810 654618 347046 654854
rect 344426 633818 344662 634054
rect 344746 633818 344982 634054
rect 344426 633498 344662 633734
rect 344746 633498 344982 633734
rect 70330 618938 70566 619174
rect 70330 618618 70566 618854
rect 101050 618938 101286 619174
rect 101050 618618 101286 618854
rect 131770 618938 132006 619174
rect 131770 618618 132006 618854
rect 162490 618938 162726 619174
rect 162490 618618 162726 618854
rect 193210 618938 193446 619174
rect 193210 618618 193446 618854
rect 223930 618938 224166 619174
rect 223930 618618 224166 618854
rect 254650 618938 254886 619174
rect 254650 618618 254886 618854
rect 285370 618938 285606 619174
rect 285370 618618 285606 618854
rect 316090 618938 316326 619174
rect 316090 618618 316326 618854
rect 54970 615218 55206 615454
rect 54970 614898 55206 615134
rect 85690 615218 85926 615454
rect 85690 614898 85926 615134
rect 116410 615218 116646 615454
rect 116410 614898 116646 615134
rect 147130 615218 147366 615454
rect 147130 614898 147366 615134
rect 177850 615218 178086 615454
rect 177850 614898 178086 615134
rect 208570 615218 208806 615454
rect 208570 614898 208806 615134
rect 239290 615218 239526 615454
rect 239290 614898 239526 615134
rect 270010 615218 270246 615454
rect 270010 614898 270246 615134
rect 300730 615218 300966 615454
rect 300730 614898 300966 615134
rect 331450 615218 331686 615454
rect 331450 614898 331686 615134
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 348146 637538 348382 637774
rect 348466 637538 348702 637774
rect 348146 637218 348382 637454
rect 348466 637218 348702 637454
rect 346810 618938 347046 619174
rect 346810 618618 347046 618854
rect 344426 597818 344662 598054
rect 344746 597818 344982 598054
rect 344426 597498 344662 597734
rect 344746 597498 344982 597734
rect 70330 582938 70566 583174
rect 70330 582618 70566 582854
rect 101050 582938 101286 583174
rect 101050 582618 101286 582854
rect 131770 582938 132006 583174
rect 131770 582618 132006 582854
rect 162490 582938 162726 583174
rect 162490 582618 162726 582854
rect 193210 582938 193446 583174
rect 193210 582618 193446 582854
rect 223930 582938 224166 583174
rect 223930 582618 224166 582854
rect 254650 582938 254886 583174
rect 254650 582618 254886 582854
rect 285370 582938 285606 583174
rect 285370 582618 285606 582854
rect 316090 582938 316326 583174
rect 316090 582618 316326 582854
rect 54970 579218 55206 579454
rect 54970 578898 55206 579134
rect 85690 579218 85926 579454
rect 85690 578898 85926 579134
rect 116410 579218 116646 579454
rect 116410 578898 116646 579134
rect 147130 579218 147366 579454
rect 147130 578898 147366 579134
rect 177850 579218 178086 579454
rect 177850 578898 178086 579134
rect 208570 579218 208806 579454
rect 208570 578898 208806 579134
rect 239290 579218 239526 579454
rect 239290 578898 239526 579134
rect 270010 579218 270246 579454
rect 270010 578898 270246 579134
rect 300730 579218 300966 579454
rect 300730 578898 300966 579134
rect 331450 579218 331686 579454
rect 331450 578898 331686 579134
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 348146 601538 348382 601774
rect 348466 601538 348702 601774
rect 348146 601218 348382 601454
rect 348466 601218 348702 601454
rect 346810 582938 347046 583174
rect 346810 582618 347046 582854
rect 344426 561818 344662 562054
rect 344746 561818 344982 562054
rect 344426 561498 344662 561734
rect 344746 561498 344982 561734
rect 70330 546938 70566 547174
rect 70330 546618 70566 546854
rect 101050 546938 101286 547174
rect 101050 546618 101286 546854
rect 131770 546938 132006 547174
rect 131770 546618 132006 546854
rect 162490 546938 162726 547174
rect 162490 546618 162726 546854
rect 193210 546938 193446 547174
rect 193210 546618 193446 546854
rect 223930 546938 224166 547174
rect 223930 546618 224166 546854
rect 254650 546938 254886 547174
rect 254650 546618 254886 546854
rect 285370 546938 285606 547174
rect 285370 546618 285606 546854
rect 316090 546938 316326 547174
rect 316090 546618 316326 546854
rect 54970 543218 55206 543454
rect 54970 542898 55206 543134
rect 85690 543218 85926 543454
rect 85690 542898 85926 543134
rect 116410 543218 116646 543454
rect 116410 542898 116646 543134
rect 147130 543218 147366 543454
rect 147130 542898 147366 543134
rect 177850 543218 178086 543454
rect 177850 542898 178086 543134
rect 208570 543218 208806 543454
rect 208570 542898 208806 543134
rect 239290 543218 239526 543454
rect 239290 542898 239526 543134
rect 270010 543218 270246 543454
rect 270010 542898 270246 543134
rect 300730 543218 300966 543454
rect 300730 542898 300966 543134
rect 331450 543218 331686 543454
rect 331450 542898 331686 543134
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 348146 565538 348382 565774
rect 348466 565538 348702 565774
rect 348146 565218 348382 565454
rect 348466 565218 348702 565454
rect 346810 546938 347046 547174
rect 346810 546618 347046 546854
rect 344426 525818 344662 526054
rect 344746 525818 344982 526054
rect 344426 525498 344662 525734
rect 344746 525498 344982 525734
rect 70330 510938 70566 511174
rect 70330 510618 70566 510854
rect 101050 510938 101286 511174
rect 101050 510618 101286 510854
rect 131770 510938 132006 511174
rect 131770 510618 132006 510854
rect 162490 510938 162726 511174
rect 162490 510618 162726 510854
rect 193210 510938 193446 511174
rect 193210 510618 193446 510854
rect 223930 510938 224166 511174
rect 223930 510618 224166 510854
rect 254650 510938 254886 511174
rect 254650 510618 254886 510854
rect 285370 510938 285606 511174
rect 285370 510618 285606 510854
rect 316090 510938 316326 511174
rect 316090 510618 316326 510854
rect 54970 507218 55206 507454
rect 54970 506898 55206 507134
rect 85690 507218 85926 507454
rect 85690 506898 85926 507134
rect 116410 507218 116646 507454
rect 116410 506898 116646 507134
rect 147130 507218 147366 507454
rect 147130 506898 147366 507134
rect 177850 507218 178086 507454
rect 177850 506898 178086 507134
rect 208570 507218 208806 507454
rect 208570 506898 208806 507134
rect 239290 507218 239526 507454
rect 239290 506898 239526 507134
rect 270010 507218 270246 507454
rect 270010 506898 270246 507134
rect 300730 507218 300966 507454
rect 300730 506898 300966 507134
rect 331450 507218 331686 507454
rect 331450 506898 331686 507134
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 348146 529538 348382 529774
rect 348466 529538 348702 529774
rect 348146 529218 348382 529454
rect 348466 529218 348702 529454
rect 346810 510938 347046 511174
rect 346810 510618 347046 510854
rect 344426 489818 344662 490054
rect 344746 489818 344982 490054
rect 344426 489498 344662 489734
rect 344746 489498 344982 489734
rect 70330 474938 70566 475174
rect 70330 474618 70566 474854
rect 101050 474938 101286 475174
rect 101050 474618 101286 474854
rect 131770 474938 132006 475174
rect 131770 474618 132006 474854
rect 162490 474938 162726 475174
rect 162490 474618 162726 474854
rect 193210 474938 193446 475174
rect 193210 474618 193446 474854
rect 223930 474938 224166 475174
rect 223930 474618 224166 474854
rect 254650 474938 254886 475174
rect 254650 474618 254886 474854
rect 285370 474938 285606 475174
rect 285370 474618 285606 474854
rect 316090 474938 316326 475174
rect 316090 474618 316326 474854
rect 54970 471218 55206 471454
rect 54970 470898 55206 471134
rect 85690 471218 85926 471454
rect 85690 470898 85926 471134
rect 116410 471218 116646 471454
rect 116410 470898 116646 471134
rect 147130 471218 147366 471454
rect 147130 470898 147366 471134
rect 177850 471218 178086 471454
rect 177850 470898 178086 471134
rect 208570 471218 208806 471454
rect 208570 470898 208806 471134
rect 239290 471218 239526 471454
rect 239290 470898 239526 471134
rect 270010 471218 270246 471454
rect 270010 470898 270246 471134
rect 300730 471218 300966 471454
rect 300730 470898 300966 471134
rect 331450 471218 331686 471454
rect 331450 470898 331686 471134
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 348146 493538 348382 493774
rect 348466 493538 348702 493774
rect 348146 493218 348382 493454
rect 348466 493218 348702 493454
rect 346810 474938 347046 475174
rect 346810 474618 347046 474854
rect 344426 453818 344662 454054
rect 344746 453818 344982 454054
rect 344426 453498 344662 453734
rect 344746 453498 344982 453734
rect 70330 438938 70566 439174
rect 70330 438618 70566 438854
rect 101050 438938 101286 439174
rect 101050 438618 101286 438854
rect 131770 438938 132006 439174
rect 131770 438618 132006 438854
rect 162490 438938 162726 439174
rect 162490 438618 162726 438854
rect 193210 438938 193446 439174
rect 193210 438618 193446 438854
rect 223930 438938 224166 439174
rect 223930 438618 224166 438854
rect 254650 438938 254886 439174
rect 254650 438618 254886 438854
rect 285370 438938 285606 439174
rect 285370 438618 285606 438854
rect 316090 438938 316326 439174
rect 316090 438618 316326 438854
rect 54970 435218 55206 435454
rect 54970 434898 55206 435134
rect 85690 435218 85926 435454
rect 85690 434898 85926 435134
rect 116410 435218 116646 435454
rect 116410 434898 116646 435134
rect 147130 435218 147366 435454
rect 147130 434898 147366 435134
rect 177850 435218 178086 435454
rect 177850 434898 178086 435134
rect 208570 435218 208806 435454
rect 208570 434898 208806 435134
rect 239290 435218 239526 435454
rect 239290 434898 239526 435134
rect 270010 435218 270246 435454
rect 270010 434898 270246 435134
rect 300730 435218 300966 435454
rect 300730 434898 300966 435134
rect 331450 435218 331686 435454
rect 331450 434898 331686 435134
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 348146 457538 348382 457774
rect 348466 457538 348702 457774
rect 348146 457218 348382 457454
rect 348466 457218 348702 457454
rect 346810 438938 347046 439174
rect 346810 438618 347046 438854
rect 344426 417818 344662 418054
rect 344746 417818 344982 418054
rect 344426 417498 344662 417734
rect 344746 417498 344982 417734
rect 70330 402938 70566 403174
rect 70330 402618 70566 402854
rect 101050 402938 101286 403174
rect 101050 402618 101286 402854
rect 131770 402938 132006 403174
rect 131770 402618 132006 402854
rect 162490 402938 162726 403174
rect 162490 402618 162726 402854
rect 193210 402938 193446 403174
rect 193210 402618 193446 402854
rect 223930 402938 224166 403174
rect 223930 402618 224166 402854
rect 254650 402938 254886 403174
rect 254650 402618 254886 402854
rect 285370 402938 285606 403174
rect 285370 402618 285606 402854
rect 316090 402938 316326 403174
rect 316090 402618 316326 402854
rect 54970 399218 55206 399454
rect 54970 398898 55206 399134
rect 85690 399218 85926 399454
rect 85690 398898 85926 399134
rect 116410 399218 116646 399454
rect 116410 398898 116646 399134
rect 147130 399218 147366 399454
rect 147130 398898 147366 399134
rect 177850 399218 178086 399454
rect 177850 398898 178086 399134
rect 208570 399218 208806 399454
rect 208570 398898 208806 399134
rect 239290 399218 239526 399454
rect 239290 398898 239526 399134
rect 270010 399218 270246 399454
rect 270010 398898 270246 399134
rect 300730 399218 300966 399454
rect 300730 398898 300966 399134
rect 331450 399218 331686 399454
rect 331450 398898 331686 399134
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 348146 421538 348382 421774
rect 348466 421538 348702 421774
rect 348146 421218 348382 421454
rect 348466 421218 348702 421454
rect 346810 402938 347046 403174
rect 346810 402618 347046 402854
rect 344426 381818 344662 382054
rect 344746 381818 344982 382054
rect 344426 381498 344662 381734
rect 344746 381498 344982 381734
rect 70330 366938 70566 367174
rect 70330 366618 70566 366854
rect 101050 366938 101286 367174
rect 101050 366618 101286 366854
rect 131770 366938 132006 367174
rect 131770 366618 132006 366854
rect 162490 366938 162726 367174
rect 162490 366618 162726 366854
rect 193210 366938 193446 367174
rect 193210 366618 193446 366854
rect 223930 366938 224166 367174
rect 223930 366618 224166 366854
rect 254650 366938 254886 367174
rect 254650 366618 254886 366854
rect 285370 366938 285606 367174
rect 285370 366618 285606 366854
rect 316090 366938 316326 367174
rect 316090 366618 316326 366854
rect 54970 363218 55206 363454
rect 54970 362898 55206 363134
rect 85690 363218 85926 363454
rect 85690 362898 85926 363134
rect 116410 363218 116646 363454
rect 116410 362898 116646 363134
rect 147130 363218 147366 363454
rect 147130 362898 147366 363134
rect 177850 363218 178086 363454
rect 177850 362898 178086 363134
rect 208570 363218 208806 363454
rect 208570 362898 208806 363134
rect 239290 363218 239526 363454
rect 239290 362898 239526 363134
rect 270010 363218 270246 363454
rect 270010 362898 270246 363134
rect 300730 363218 300966 363454
rect 300730 362898 300966 363134
rect 331450 363218 331686 363454
rect 331450 362898 331686 363134
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 348146 385538 348382 385774
rect 348466 385538 348702 385774
rect 348146 385218 348382 385454
rect 348466 385218 348702 385454
rect 346810 366938 347046 367174
rect 346810 366618 347046 366854
rect 344426 345818 344662 346054
rect 344746 345818 344982 346054
rect 344426 345498 344662 345734
rect 344746 345498 344982 345734
rect 70330 330938 70566 331174
rect 70330 330618 70566 330854
rect 101050 330938 101286 331174
rect 101050 330618 101286 330854
rect 131770 330938 132006 331174
rect 131770 330618 132006 330854
rect 162490 330938 162726 331174
rect 162490 330618 162726 330854
rect 193210 330938 193446 331174
rect 193210 330618 193446 330854
rect 223930 330938 224166 331174
rect 223930 330618 224166 330854
rect 254650 330938 254886 331174
rect 254650 330618 254886 330854
rect 285370 330938 285606 331174
rect 285370 330618 285606 330854
rect 316090 330938 316326 331174
rect 316090 330618 316326 330854
rect 54970 327218 55206 327454
rect 54970 326898 55206 327134
rect 85690 327218 85926 327454
rect 85690 326898 85926 327134
rect 116410 327218 116646 327454
rect 116410 326898 116646 327134
rect 147130 327218 147366 327454
rect 147130 326898 147366 327134
rect 177850 327218 178086 327454
rect 177850 326898 178086 327134
rect 208570 327218 208806 327454
rect 208570 326898 208806 327134
rect 239290 327218 239526 327454
rect 239290 326898 239526 327134
rect 270010 327218 270246 327454
rect 270010 326898 270246 327134
rect 300730 327218 300966 327454
rect 300730 326898 300966 327134
rect 331450 327218 331686 327454
rect 331450 326898 331686 327134
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 348146 349538 348382 349774
rect 348466 349538 348702 349774
rect 348146 349218 348382 349454
rect 348466 349218 348702 349454
rect 346810 330938 347046 331174
rect 346810 330618 347046 330854
rect 344426 309818 344662 310054
rect 344746 309818 344982 310054
rect 344426 309498 344662 309734
rect 344746 309498 344982 309734
rect 70330 294938 70566 295174
rect 70330 294618 70566 294854
rect 101050 294938 101286 295174
rect 101050 294618 101286 294854
rect 131770 294938 132006 295174
rect 131770 294618 132006 294854
rect 162490 294938 162726 295174
rect 162490 294618 162726 294854
rect 193210 294938 193446 295174
rect 193210 294618 193446 294854
rect 223930 294938 224166 295174
rect 223930 294618 224166 294854
rect 254650 294938 254886 295174
rect 254650 294618 254886 294854
rect 285370 294938 285606 295174
rect 285370 294618 285606 294854
rect 316090 294938 316326 295174
rect 316090 294618 316326 294854
rect 54970 291218 55206 291454
rect 54970 290898 55206 291134
rect 85690 291218 85926 291454
rect 85690 290898 85926 291134
rect 116410 291218 116646 291454
rect 116410 290898 116646 291134
rect 147130 291218 147366 291454
rect 147130 290898 147366 291134
rect 177850 291218 178086 291454
rect 177850 290898 178086 291134
rect 208570 291218 208806 291454
rect 208570 290898 208806 291134
rect 239290 291218 239526 291454
rect 239290 290898 239526 291134
rect 270010 291218 270246 291454
rect 270010 290898 270246 291134
rect 300730 291218 300966 291454
rect 300730 290898 300966 291134
rect 331450 291218 331686 291454
rect 331450 290898 331686 291134
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 348146 313538 348382 313774
rect 348466 313538 348702 313774
rect 348146 313218 348382 313454
rect 348466 313218 348702 313454
rect 346810 294938 347046 295174
rect 346810 294618 347046 294854
rect 344426 273818 344662 274054
rect 344746 273818 344982 274054
rect 344426 273498 344662 273734
rect 344746 273498 344982 273734
rect 70330 258938 70566 259174
rect 70330 258618 70566 258854
rect 101050 258938 101286 259174
rect 101050 258618 101286 258854
rect 131770 258938 132006 259174
rect 131770 258618 132006 258854
rect 162490 258938 162726 259174
rect 162490 258618 162726 258854
rect 193210 258938 193446 259174
rect 193210 258618 193446 258854
rect 223930 258938 224166 259174
rect 223930 258618 224166 258854
rect 254650 258938 254886 259174
rect 254650 258618 254886 258854
rect 285370 258938 285606 259174
rect 285370 258618 285606 258854
rect 316090 258938 316326 259174
rect 316090 258618 316326 258854
rect 54970 255218 55206 255454
rect 54970 254898 55206 255134
rect 85690 255218 85926 255454
rect 85690 254898 85926 255134
rect 116410 255218 116646 255454
rect 116410 254898 116646 255134
rect 147130 255218 147366 255454
rect 147130 254898 147366 255134
rect 177850 255218 178086 255454
rect 177850 254898 178086 255134
rect 208570 255218 208806 255454
rect 208570 254898 208806 255134
rect 239290 255218 239526 255454
rect 239290 254898 239526 255134
rect 270010 255218 270246 255454
rect 270010 254898 270246 255134
rect 300730 255218 300966 255454
rect 300730 254898 300966 255134
rect 331450 255218 331686 255454
rect 331450 254898 331686 255134
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 348146 277538 348382 277774
rect 348466 277538 348702 277774
rect 348146 277218 348382 277454
rect 348466 277218 348702 277454
rect 346810 258938 347046 259174
rect 346810 258618 347046 258854
rect 344426 237818 344662 238054
rect 344746 237818 344982 238054
rect 344426 237498 344662 237734
rect 344746 237498 344982 237734
rect 70330 222938 70566 223174
rect 70330 222618 70566 222854
rect 101050 222938 101286 223174
rect 101050 222618 101286 222854
rect 131770 222938 132006 223174
rect 131770 222618 132006 222854
rect 162490 222938 162726 223174
rect 162490 222618 162726 222854
rect 193210 222938 193446 223174
rect 193210 222618 193446 222854
rect 223930 222938 224166 223174
rect 223930 222618 224166 222854
rect 254650 222938 254886 223174
rect 254650 222618 254886 222854
rect 285370 222938 285606 223174
rect 285370 222618 285606 222854
rect 316090 222938 316326 223174
rect 316090 222618 316326 222854
rect 54970 219218 55206 219454
rect 54970 218898 55206 219134
rect 85690 219218 85926 219454
rect 85690 218898 85926 219134
rect 116410 219218 116646 219454
rect 116410 218898 116646 219134
rect 147130 219218 147366 219454
rect 147130 218898 147366 219134
rect 177850 219218 178086 219454
rect 177850 218898 178086 219134
rect 208570 219218 208806 219454
rect 208570 218898 208806 219134
rect 239290 219218 239526 219454
rect 239290 218898 239526 219134
rect 270010 219218 270246 219454
rect 270010 218898 270246 219134
rect 300730 219218 300966 219454
rect 300730 218898 300966 219134
rect 331450 219218 331686 219454
rect 331450 218898 331686 219134
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 348146 241538 348382 241774
rect 348466 241538 348702 241774
rect 348146 241218 348382 241454
rect 348466 241218 348702 241454
rect 346810 222938 347046 223174
rect 346810 222618 347046 222854
rect 344426 201818 344662 202054
rect 344746 201818 344982 202054
rect 344426 201498 344662 201734
rect 344746 201498 344982 201734
rect 70330 186938 70566 187174
rect 70330 186618 70566 186854
rect 101050 186938 101286 187174
rect 101050 186618 101286 186854
rect 131770 186938 132006 187174
rect 131770 186618 132006 186854
rect 162490 186938 162726 187174
rect 162490 186618 162726 186854
rect 193210 186938 193446 187174
rect 193210 186618 193446 186854
rect 223930 186938 224166 187174
rect 223930 186618 224166 186854
rect 254650 186938 254886 187174
rect 254650 186618 254886 186854
rect 285370 186938 285606 187174
rect 285370 186618 285606 186854
rect 316090 186938 316326 187174
rect 316090 186618 316326 186854
rect 54970 183218 55206 183454
rect 54970 182898 55206 183134
rect 85690 183218 85926 183454
rect 85690 182898 85926 183134
rect 116410 183218 116646 183454
rect 116410 182898 116646 183134
rect 147130 183218 147366 183454
rect 147130 182898 147366 183134
rect 177850 183218 178086 183454
rect 177850 182898 178086 183134
rect 208570 183218 208806 183454
rect 208570 182898 208806 183134
rect 239290 183218 239526 183454
rect 239290 182898 239526 183134
rect 270010 183218 270246 183454
rect 270010 182898 270246 183134
rect 300730 183218 300966 183454
rect 300730 182898 300966 183134
rect 331450 183218 331686 183454
rect 331450 182898 331686 183134
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 348146 205538 348382 205774
rect 348466 205538 348702 205774
rect 348146 205218 348382 205454
rect 348466 205218 348702 205454
rect 346810 186938 347046 187174
rect 346810 186618 347046 186854
rect 344426 165818 344662 166054
rect 344746 165818 344982 166054
rect 344426 165498 344662 165734
rect 344746 165498 344982 165734
rect 70330 150938 70566 151174
rect 70330 150618 70566 150854
rect 101050 150938 101286 151174
rect 101050 150618 101286 150854
rect 131770 150938 132006 151174
rect 131770 150618 132006 150854
rect 162490 150938 162726 151174
rect 162490 150618 162726 150854
rect 193210 150938 193446 151174
rect 193210 150618 193446 150854
rect 223930 150938 224166 151174
rect 223930 150618 224166 150854
rect 254650 150938 254886 151174
rect 254650 150618 254886 150854
rect 285370 150938 285606 151174
rect 285370 150618 285606 150854
rect 316090 150938 316326 151174
rect 316090 150618 316326 150854
rect 54970 147218 55206 147454
rect 54970 146898 55206 147134
rect 85690 147218 85926 147454
rect 85690 146898 85926 147134
rect 116410 147218 116646 147454
rect 116410 146898 116646 147134
rect 147130 147218 147366 147454
rect 147130 146898 147366 147134
rect 177850 147218 178086 147454
rect 177850 146898 178086 147134
rect 208570 147218 208806 147454
rect 208570 146898 208806 147134
rect 239290 147218 239526 147454
rect 239290 146898 239526 147134
rect 270010 147218 270246 147454
rect 270010 146898 270246 147134
rect 300730 147218 300966 147454
rect 300730 146898 300966 147134
rect 331450 147218 331686 147454
rect 331450 146898 331686 147134
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 348146 169538 348382 169774
rect 348466 169538 348702 169774
rect 348146 169218 348382 169454
rect 348466 169218 348702 169454
rect 346810 150938 347046 151174
rect 346810 150618 347046 150854
rect 344426 129818 344662 130054
rect 344746 129818 344982 130054
rect 344426 129498 344662 129734
rect 344746 129498 344982 129734
rect 70330 114938 70566 115174
rect 70330 114618 70566 114854
rect 101050 114938 101286 115174
rect 101050 114618 101286 114854
rect 131770 114938 132006 115174
rect 131770 114618 132006 114854
rect 162490 114938 162726 115174
rect 162490 114618 162726 114854
rect 193210 114938 193446 115174
rect 193210 114618 193446 114854
rect 223930 114938 224166 115174
rect 223930 114618 224166 114854
rect 254650 114938 254886 115174
rect 254650 114618 254886 114854
rect 285370 114938 285606 115174
rect 285370 114618 285606 114854
rect 316090 114938 316326 115174
rect 316090 114618 316326 114854
rect 54970 111218 55206 111454
rect 54970 110898 55206 111134
rect 85690 111218 85926 111454
rect 85690 110898 85926 111134
rect 116410 111218 116646 111454
rect 116410 110898 116646 111134
rect 147130 111218 147366 111454
rect 147130 110898 147366 111134
rect 177850 111218 178086 111454
rect 177850 110898 178086 111134
rect 208570 111218 208806 111454
rect 208570 110898 208806 111134
rect 239290 111218 239526 111454
rect 239290 110898 239526 111134
rect 270010 111218 270246 111454
rect 270010 110898 270246 111134
rect 300730 111218 300966 111454
rect 300730 110898 300966 111134
rect 331450 111218 331686 111454
rect 331450 110898 331686 111134
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 348146 133538 348382 133774
rect 348466 133538 348702 133774
rect 348146 133218 348382 133454
rect 348466 133218 348702 133454
rect 346810 114938 347046 115174
rect 346810 114618 347046 114854
rect 344426 93818 344662 94054
rect 344746 93818 344982 94054
rect 344426 93498 344662 93734
rect 344746 93498 344982 93734
rect 70330 78938 70566 79174
rect 70330 78618 70566 78854
rect 101050 78938 101286 79174
rect 101050 78618 101286 78854
rect 131770 78938 132006 79174
rect 131770 78618 132006 78854
rect 162490 78938 162726 79174
rect 162490 78618 162726 78854
rect 193210 78938 193446 79174
rect 193210 78618 193446 78854
rect 223930 78938 224166 79174
rect 223930 78618 224166 78854
rect 254650 78938 254886 79174
rect 254650 78618 254886 78854
rect 285370 78938 285606 79174
rect 285370 78618 285606 78854
rect 316090 78938 316326 79174
rect 316090 78618 316326 78854
rect 54970 75218 55206 75454
rect 54970 74898 55206 75134
rect 85690 75218 85926 75454
rect 85690 74898 85926 75134
rect 116410 75218 116646 75454
rect 116410 74898 116646 75134
rect 147130 75218 147366 75454
rect 147130 74898 147366 75134
rect 177850 75218 178086 75454
rect 177850 74898 178086 75134
rect 208570 75218 208806 75454
rect 208570 74898 208806 75134
rect 239290 75218 239526 75454
rect 239290 74898 239526 75134
rect 270010 75218 270246 75454
rect 270010 74898 270246 75134
rect 300730 75218 300966 75454
rect 300730 74898 300966 75134
rect 331450 75218 331686 75454
rect 331450 74898 331686 75134
rect 348146 97538 348382 97774
rect 348466 97538 348702 97774
rect 348146 97218 348382 97454
rect 348466 97218 348702 97454
rect 346810 78938 347046 79174
rect 346810 78618 347046 78854
rect 344426 57818 344662 58054
rect 344746 57818 344982 58054
rect 344426 57498 344662 57734
rect 344746 57498 344982 57734
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 48986 -3462 49222 -3226
rect 49306 -3462 49542 -3226
rect 48986 -3782 49222 -3546
rect 49306 -3782 49542 -3546
rect 52706 54098 52942 54334
rect 53026 54098 53262 54334
rect 52706 53778 52942 54014
rect 53026 53778 53262 54014
rect 52706 18098 52942 18334
rect 53026 18098 53262 18334
rect 52706 17778 52942 18014
rect 53026 17778 53262 18014
rect 52706 -4422 52942 -4186
rect 53026 -4422 53262 -4186
rect 52706 -4742 52942 -4506
rect 53026 -4742 53262 -4506
rect 56426 21818 56662 22054
rect 56746 21818 56982 22054
rect 56426 21498 56662 21734
rect 56746 21498 56982 21734
rect 56426 -5382 56662 -5146
rect 56746 -5382 56982 -5146
rect 56426 -5702 56662 -5466
rect 56746 -5702 56982 -5466
rect 60146 25538 60382 25774
rect 60466 25538 60702 25774
rect 60146 25218 60382 25454
rect 60466 25218 60702 25454
rect 60146 -6342 60382 -6106
rect 60466 -6342 60702 -6106
rect 60146 -6662 60382 -6426
rect 60466 -6662 60702 -6426
rect 63866 29258 64102 29494
rect 64186 29258 64422 29494
rect 63866 28938 64102 29174
rect 64186 28938 64422 29174
rect 63866 -7302 64102 -7066
rect 64186 -7302 64422 -7066
rect 63866 -7622 64102 -7386
rect 64186 -7622 64422 -7386
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -1542 77782 -1306
rect 77866 -1542 78102 -1306
rect 77546 -1862 77782 -1626
rect 77866 -1862 78102 -1626
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -2502 81502 -2266
rect 81586 -2502 81822 -2266
rect 81266 -2822 81502 -2586
rect 81586 -2822 81822 -2586
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 84986 -3462 85222 -3226
rect 85306 -3462 85542 -3226
rect 84986 -3782 85222 -3546
rect 85306 -3782 85542 -3546
rect 88706 54098 88942 54334
rect 89026 54098 89262 54334
rect 88706 53778 88942 54014
rect 89026 53778 89262 54014
rect 88706 18098 88942 18334
rect 89026 18098 89262 18334
rect 88706 17778 88942 18014
rect 89026 17778 89262 18014
rect 88706 -4422 88942 -4186
rect 89026 -4422 89262 -4186
rect 88706 -4742 88942 -4506
rect 89026 -4742 89262 -4506
rect 92426 21818 92662 22054
rect 92746 21818 92982 22054
rect 92426 21498 92662 21734
rect 92746 21498 92982 21734
rect 92426 -5382 92662 -5146
rect 92746 -5382 92982 -5146
rect 92426 -5702 92662 -5466
rect 92746 -5702 92982 -5466
rect 96146 25538 96382 25774
rect 96466 25538 96702 25774
rect 96146 25218 96382 25454
rect 96466 25218 96702 25454
rect 96146 -6342 96382 -6106
rect 96466 -6342 96702 -6106
rect 96146 -6662 96382 -6426
rect 96466 -6662 96702 -6426
rect 99866 29258 100102 29494
rect 100186 29258 100422 29494
rect 99866 28938 100102 29174
rect 100186 28938 100422 29174
rect 99866 -7302 100102 -7066
rect 100186 -7302 100422 -7066
rect 99866 -7622 100102 -7386
rect 100186 -7622 100422 -7386
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -1542 113782 -1306
rect 113866 -1542 114102 -1306
rect 113546 -1862 113782 -1626
rect 113866 -1862 114102 -1626
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -2502 117502 -2266
rect 117586 -2502 117822 -2266
rect 117266 -2822 117502 -2586
rect 117586 -2822 117822 -2586
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 120986 -3462 121222 -3226
rect 121306 -3462 121542 -3226
rect 120986 -3782 121222 -3546
rect 121306 -3782 121542 -3546
rect 124706 54098 124942 54334
rect 125026 54098 125262 54334
rect 124706 53778 124942 54014
rect 125026 53778 125262 54014
rect 124706 18098 124942 18334
rect 125026 18098 125262 18334
rect 124706 17778 124942 18014
rect 125026 17778 125262 18014
rect 124706 -4422 124942 -4186
rect 125026 -4422 125262 -4186
rect 124706 -4742 124942 -4506
rect 125026 -4742 125262 -4506
rect 128426 21818 128662 22054
rect 128746 21818 128982 22054
rect 128426 21498 128662 21734
rect 128746 21498 128982 21734
rect 128426 -5382 128662 -5146
rect 128746 -5382 128982 -5146
rect 128426 -5702 128662 -5466
rect 128746 -5702 128982 -5466
rect 132146 25538 132382 25774
rect 132466 25538 132702 25774
rect 132146 25218 132382 25454
rect 132466 25218 132702 25454
rect 132146 -6342 132382 -6106
rect 132466 -6342 132702 -6106
rect 132146 -6662 132382 -6426
rect 132466 -6662 132702 -6426
rect 135866 29258 136102 29494
rect 136186 29258 136422 29494
rect 135866 28938 136102 29174
rect 136186 28938 136422 29174
rect 135866 -7302 136102 -7066
rect 136186 -7302 136422 -7066
rect 135866 -7622 136102 -7386
rect 136186 -7622 136422 -7386
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -1542 149782 -1306
rect 149866 -1542 150102 -1306
rect 149546 -1862 149782 -1626
rect 149866 -1862 150102 -1626
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -2502 153502 -2266
rect 153586 -2502 153822 -2266
rect 153266 -2822 153502 -2586
rect 153586 -2822 153822 -2586
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 156986 -3462 157222 -3226
rect 157306 -3462 157542 -3226
rect 156986 -3782 157222 -3546
rect 157306 -3782 157542 -3546
rect 160706 54098 160942 54334
rect 161026 54098 161262 54334
rect 160706 53778 160942 54014
rect 161026 53778 161262 54014
rect 160706 18098 160942 18334
rect 161026 18098 161262 18334
rect 160706 17778 160942 18014
rect 161026 17778 161262 18014
rect 160706 -4422 160942 -4186
rect 161026 -4422 161262 -4186
rect 160706 -4742 160942 -4506
rect 161026 -4742 161262 -4506
rect 164426 21818 164662 22054
rect 164746 21818 164982 22054
rect 164426 21498 164662 21734
rect 164746 21498 164982 21734
rect 164426 -5382 164662 -5146
rect 164746 -5382 164982 -5146
rect 164426 -5702 164662 -5466
rect 164746 -5702 164982 -5466
rect 168146 25538 168382 25774
rect 168466 25538 168702 25774
rect 168146 25218 168382 25454
rect 168466 25218 168702 25454
rect 168146 -6342 168382 -6106
rect 168466 -6342 168702 -6106
rect 168146 -6662 168382 -6426
rect 168466 -6662 168702 -6426
rect 171866 29258 172102 29494
rect 172186 29258 172422 29494
rect 171866 28938 172102 29174
rect 172186 28938 172422 29174
rect 171866 -7302 172102 -7066
rect 172186 -7302 172422 -7066
rect 171866 -7622 172102 -7386
rect 172186 -7622 172422 -7386
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -1542 185782 -1306
rect 185866 -1542 186102 -1306
rect 185546 -1862 185782 -1626
rect 185866 -1862 186102 -1626
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 196706 54098 196942 54334
rect 197026 54098 197262 54334
rect 196706 53778 196942 54014
rect 197026 53778 197262 54014
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -2502 189502 -2266
rect 189586 -2502 189822 -2266
rect 189266 -2822 189502 -2586
rect 189586 -2822 189822 -2586
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 192986 -3462 193222 -3226
rect 193306 -3462 193542 -3226
rect 192986 -3782 193222 -3546
rect 193306 -3782 193542 -3546
rect 196706 18098 196942 18334
rect 197026 18098 197262 18334
rect 196706 17778 196942 18014
rect 197026 17778 197262 18014
rect 196706 -4422 196942 -4186
rect 197026 -4422 197262 -4186
rect 196706 -4742 196942 -4506
rect 197026 -4742 197262 -4506
rect 200426 21818 200662 22054
rect 200746 21818 200982 22054
rect 200426 21498 200662 21734
rect 200746 21498 200982 21734
rect 200426 -5382 200662 -5146
rect 200746 -5382 200982 -5146
rect 200426 -5702 200662 -5466
rect 200746 -5702 200982 -5466
rect 204146 25538 204382 25774
rect 204466 25538 204702 25774
rect 204146 25218 204382 25454
rect 204466 25218 204702 25454
rect 204146 -6342 204382 -6106
rect 204466 -6342 204702 -6106
rect 204146 -6662 204382 -6426
rect 204466 -6662 204702 -6426
rect 207866 29258 208102 29494
rect 208186 29258 208422 29494
rect 207866 28938 208102 29174
rect 208186 28938 208422 29174
rect 207866 -7302 208102 -7066
rect 208186 -7302 208422 -7066
rect 207866 -7622 208102 -7386
rect 208186 -7622 208422 -7386
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -1542 221782 -1306
rect 221866 -1542 222102 -1306
rect 221546 -1862 221782 -1626
rect 221866 -1862 222102 -1626
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -2502 225502 -2266
rect 225586 -2502 225822 -2266
rect 225266 -2822 225502 -2586
rect 225586 -2822 225822 -2586
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 228986 -3462 229222 -3226
rect 229306 -3462 229542 -3226
rect 228986 -3782 229222 -3546
rect 229306 -3782 229542 -3546
rect 232706 54098 232942 54334
rect 233026 54098 233262 54334
rect 232706 53778 232942 54014
rect 233026 53778 233262 54014
rect 232706 18098 232942 18334
rect 233026 18098 233262 18334
rect 232706 17778 232942 18014
rect 233026 17778 233262 18014
rect 232706 -4422 232942 -4186
rect 233026 -4422 233262 -4186
rect 232706 -4742 232942 -4506
rect 233026 -4742 233262 -4506
rect 236426 21818 236662 22054
rect 236746 21818 236982 22054
rect 236426 21498 236662 21734
rect 236746 21498 236982 21734
rect 236426 -5382 236662 -5146
rect 236746 -5382 236982 -5146
rect 236426 -5702 236662 -5466
rect 236746 -5702 236982 -5466
rect 240146 25538 240382 25774
rect 240466 25538 240702 25774
rect 240146 25218 240382 25454
rect 240466 25218 240702 25454
rect 240146 -6342 240382 -6106
rect 240466 -6342 240702 -6106
rect 240146 -6662 240382 -6426
rect 240466 -6662 240702 -6426
rect 243866 29258 244102 29494
rect 244186 29258 244422 29494
rect 243866 28938 244102 29174
rect 244186 28938 244422 29174
rect 243866 -7302 244102 -7066
rect 244186 -7302 244422 -7066
rect 243866 -7622 244102 -7386
rect 244186 -7622 244422 -7386
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -1542 257782 -1306
rect 257866 -1542 258102 -1306
rect 257546 -1862 257782 -1626
rect 257866 -1862 258102 -1626
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -2502 261502 -2266
rect 261586 -2502 261822 -2266
rect 261266 -2822 261502 -2586
rect 261586 -2822 261822 -2586
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 264986 -3462 265222 -3226
rect 265306 -3462 265542 -3226
rect 264986 -3782 265222 -3546
rect 265306 -3782 265542 -3546
rect 268706 54098 268942 54334
rect 269026 54098 269262 54334
rect 268706 53778 268942 54014
rect 269026 53778 269262 54014
rect 268706 18098 268942 18334
rect 269026 18098 269262 18334
rect 268706 17778 268942 18014
rect 269026 17778 269262 18014
rect 268706 -4422 268942 -4186
rect 269026 -4422 269262 -4186
rect 268706 -4742 268942 -4506
rect 269026 -4742 269262 -4506
rect 272426 21818 272662 22054
rect 272746 21818 272982 22054
rect 272426 21498 272662 21734
rect 272746 21498 272982 21734
rect 272426 -5382 272662 -5146
rect 272746 -5382 272982 -5146
rect 272426 -5702 272662 -5466
rect 272746 -5702 272982 -5466
rect 276146 25538 276382 25774
rect 276466 25538 276702 25774
rect 276146 25218 276382 25454
rect 276466 25218 276702 25454
rect 276146 -6342 276382 -6106
rect 276466 -6342 276702 -6106
rect 276146 -6662 276382 -6426
rect 276466 -6662 276702 -6426
rect 279866 29258 280102 29494
rect 280186 29258 280422 29494
rect 279866 28938 280102 29174
rect 280186 28938 280422 29174
rect 279866 -7302 280102 -7066
rect 280186 -7302 280422 -7066
rect 279866 -7622 280102 -7386
rect 280186 -7622 280422 -7386
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -1542 293782 -1306
rect 293866 -1542 294102 -1306
rect 293546 -1862 293782 -1626
rect 293866 -1862 294102 -1626
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 304706 54098 304942 54334
rect 305026 54098 305262 54334
rect 304706 53778 304942 54014
rect 305026 53778 305262 54014
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -2502 297502 -2266
rect 297586 -2502 297822 -2266
rect 297266 -2822 297502 -2586
rect 297586 -2822 297822 -2586
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 300986 -3462 301222 -3226
rect 301306 -3462 301542 -3226
rect 300986 -3782 301222 -3546
rect 301306 -3782 301542 -3546
rect 304706 18098 304942 18334
rect 305026 18098 305262 18334
rect 304706 17778 304942 18014
rect 305026 17778 305262 18014
rect 304706 -4422 304942 -4186
rect 305026 -4422 305262 -4186
rect 304706 -4742 304942 -4506
rect 305026 -4742 305262 -4506
rect 308426 21818 308662 22054
rect 308746 21818 308982 22054
rect 308426 21498 308662 21734
rect 308746 21498 308982 21734
rect 308426 -5382 308662 -5146
rect 308746 -5382 308982 -5146
rect 308426 -5702 308662 -5466
rect 308746 -5702 308982 -5466
rect 312146 25538 312382 25774
rect 312466 25538 312702 25774
rect 312146 25218 312382 25454
rect 312466 25218 312702 25454
rect 312146 -6342 312382 -6106
rect 312466 -6342 312702 -6106
rect 312146 -6662 312382 -6426
rect 312466 -6662 312702 -6426
rect 315866 29258 316102 29494
rect 316186 29258 316422 29494
rect 315866 28938 316102 29174
rect 316186 28938 316422 29174
rect 315866 -7302 316102 -7066
rect 316186 -7302 316422 -7066
rect 315866 -7622 316102 -7386
rect 316186 -7622 316422 -7386
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -1542 329782 -1306
rect 329866 -1542 330102 -1306
rect 329546 -1862 329782 -1626
rect 329866 -1862 330102 -1626
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -2502 333502 -2266
rect 333586 -2502 333822 -2266
rect 333266 -2822 333502 -2586
rect 333586 -2822 333822 -2586
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 336986 -3462 337222 -3226
rect 337306 -3462 337542 -3226
rect 336986 -3782 337222 -3546
rect 337306 -3782 337542 -3546
rect 340706 54098 340942 54334
rect 341026 54098 341262 54334
rect 340706 53778 340942 54014
rect 341026 53778 341262 54014
rect 340706 18098 340942 18334
rect 341026 18098 341262 18334
rect 340706 17778 340942 18014
rect 341026 17778 341262 18014
rect 340706 -4422 340942 -4186
rect 341026 -4422 341262 -4186
rect 340706 -4742 340942 -4506
rect 341026 -4742 341262 -4506
rect 344426 21818 344662 22054
rect 344746 21818 344982 22054
rect 344426 21498 344662 21734
rect 344746 21498 344982 21734
rect 344426 -5382 344662 -5146
rect 344746 -5382 344982 -5146
rect 344426 -5702 344662 -5466
rect 344746 -5702 344982 -5466
rect 348146 61538 348382 61774
rect 348466 61538 348702 61774
rect 348146 61218 348382 61454
rect 348466 61218 348702 61454
rect 348146 25538 348382 25774
rect 348466 25538 348702 25774
rect 348146 25218 348382 25454
rect 348466 25218 348702 25454
rect 348146 -6342 348382 -6106
rect 348466 -6342 348702 -6106
rect 348146 -6662 348382 -6426
rect 348466 -6662 348702 -6426
rect 351866 711322 352102 711558
rect 352186 711322 352422 711558
rect 351866 711002 352102 711238
rect 352186 711002 352422 711238
rect 351866 677258 352102 677494
rect 352186 677258 352422 677494
rect 351866 676938 352102 677174
rect 352186 676938 352422 677174
rect 351866 641258 352102 641494
rect 352186 641258 352422 641494
rect 351866 640938 352102 641174
rect 352186 640938 352422 641174
rect 351866 605258 352102 605494
rect 352186 605258 352422 605494
rect 351866 604938 352102 605174
rect 352186 604938 352422 605174
rect 351866 569258 352102 569494
rect 352186 569258 352422 569494
rect 351866 568938 352102 569174
rect 352186 568938 352422 569174
rect 351866 533258 352102 533494
rect 352186 533258 352422 533494
rect 351866 532938 352102 533174
rect 352186 532938 352422 533174
rect 351866 497258 352102 497494
rect 352186 497258 352422 497494
rect 351866 496938 352102 497174
rect 352186 496938 352422 497174
rect 351866 461258 352102 461494
rect 352186 461258 352422 461494
rect 351866 460938 352102 461174
rect 352186 460938 352422 461174
rect 351866 425258 352102 425494
rect 352186 425258 352422 425494
rect 351866 424938 352102 425174
rect 352186 424938 352422 425174
rect 351866 389258 352102 389494
rect 352186 389258 352422 389494
rect 351866 388938 352102 389174
rect 352186 388938 352422 389174
rect 351866 353258 352102 353494
rect 352186 353258 352422 353494
rect 351866 352938 352102 353174
rect 352186 352938 352422 353174
rect 351866 317258 352102 317494
rect 352186 317258 352422 317494
rect 351866 316938 352102 317174
rect 352186 316938 352422 317174
rect 351866 281258 352102 281494
rect 352186 281258 352422 281494
rect 351866 280938 352102 281174
rect 352186 280938 352422 281174
rect 351866 245258 352102 245494
rect 352186 245258 352422 245494
rect 351866 244938 352102 245174
rect 352186 244938 352422 245174
rect 351866 209258 352102 209494
rect 352186 209258 352422 209494
rect 351866 208938 352102 209174
rect 352186 208938 352422 209174
rect 351866 173258 352102 173494
rect 352186 173258 352422 173494
rect 351866 172938 352102 173174
rect 352186 172938 352422 173174
rect 351866 137258 352102 137494
rect 352186 137258 352422 137494
rect 351866 136938 352102 137174
rect 352186 136938 352422 137174
rect 351866 101258 352102 101494
rect 352186 101258 352422 101494
rect 351866 100938 352102 101174
rect 352186 100938 352422 101174
rect 351866 65258 352102 65494
rect 352186 65258 352422 65494
rect 351866 64938 352102 65174
rect 352186 64938 352422 65174
rect 351866 29258 352102 29494
rect 352186 29258 352422 29494
rect 351866 28938 352102 29174
rect 352186 28938 352422 29174
rect 351866 -7302 352102 -7066
rect 352186 -7302 352422 -7066
rect 351866 -7622 352102 -7386
rect 352186 -7622 352422 -7386
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 705562 365782 705798
rect 365866 705562 366102 705798
rect 365546 705242 365782 705478
rect 365866 705242 366102 705478
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -1542 365782 -1306
rect 365866 -1542 366102 -1306
rect 365546 -1862 365782 -1626
rect 365866 -1862 366102 -1626
rect 369266 706522 369502 706758
rect 369586 706522 369822 706758
rect 369266 706202 369502 706438
rect 369586 706202 369822 706438
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -2502 369502 -2266
rect 369586 -2502 369822 -2266
rect 369266 -2822 369502 -2586
rect 369586 -2822 369822 -2586
rect 372986 707482 373222 707718
rect 373306 707482 373542 707718
rect 372986 707162 373222 707398
rect 373306 707162 373542 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 372986 -3462 373222 -3226
rect 373306 -3462 373542 -3226
rect 372986 -3782 373222 -3546
rect 373306 -3782 373542 -3546
rect 376706 708442 376942 708678
rect 377026 708442 377262 708678
rect 376706 708122 376942 708358
rect 377026 708122 377262 708358
rect 376706 666098 376942 666334
rect 377026 666098 377262 666334
rect 376706 665778 376942 666014
rect 377026 665778 377262 666014
rect 376706 630098 376942 630334
rect 377026 630098 377262 630334
rect 376706 629778 376942 630014
rect 377026 629778 377262 630014
rect 376706 594098 376942 594334
rect 377026 594098 377262 594334
rect 376706 593778 376942 594014
rect 377026 593778 377262 594014
rect 376706 558098 376942 558334
rect 377026 558098 377262 558334
rect 376706 557778 376942 558014
rect 377026 557778 377262 558014
rect 376706 522098 376942 522334
rect 377026 522098 377262 522334
rect 376706 521778 376942 522014
rect 377026 521778 377262 522014
rect 376706 486098 376942 486334
rect 377026 486098 377262 486334
rect 376706 485778 376942 486014
rect 377026 485778 377262 486014
rect 376706 450098 376942 450334
rect 377026 450098 377262 450334
rect 376706 449778 376942 450014
rect 377026 449778 377262 450014
rect 376706 414098 376942 414334
rect 377026 414098 377262 414334
rect 376706 413778 376942 414014
rect 377026 413778 377262 414014
rect 376706 378098 376942 378334
rect 377026 378098 377262 378334
rect 376706 377778 376942 378014
rect 377026 377778 377262 378014
rect 376706 342098 376942 342334
rect 377026 342098 377262 342334
rect 376706 341778 376942 342014
rect 377026 341778 377262 342014
rect 376706 306098 376942 306334
rect 377026 306098 377262 306334
rect 376706 305778 376942 306014
rect 377026 305778 377262 306014
rect 376706 270098 376942 270334
rect 377026 270098 377262 270334
rect 376706 269778 376942 270014
rect 377026 269778 377262 270014
rect 376706 234098 376942 234334
rect 377026 234098 377262 234334
rect 376706 233778 376942 234014
rect 377026 233778 377262 234014
rect 376706 198098 376942 198334
rect 377026 198098 377262 198334
rect 376706 197778 376942 198014
rect 377026 197778 377262 198014
rect 376706 162098 376942 162334
rect 377026 162098 377262 162334
rect 376706 161778 376942 162014
rect 377026 161778 377262 162014
rect 376706 126098 376942 126334
rect 377026 126098 377262 126334
rect 376706 125778 376942 126014
rect 377026 125778 377262 126014
rect 376706 90098 376942 90334
rect 377026 90098 377262 90334
rect 376706 89778 376942 90014
rect 377026 89778 377262 90014
rect 376706 54098 376942 54334
rect 377026 54098 377262 54334
rect 376706 53778 376942 54014
rect 377026 53778 377262 54014
rect 376706 18098 376942 18334
rect 377026 18098 377262 18334
rect 376706 17778 376942 18014
rect 377026 17778 377262 18014
rect 376706 -4422 376942 -4186
rect 377026 -4422 377262 -4186
rect 376706 -4742 376942 -4506
rect 377026 -4742 377262 -4506
rect 380426 709402 380662 709638
rect 380746 709402 380982 709638
rect 380426 709082 380662 709318
rect 380746 709082 380982 709318
rect 380426 669818 380662 670054
rect 380746 669818 380982 670054
rect 380426 669498 380662 669734
rect 380746 669498 380982 669734
rect 380426 633818 380662 634054
rect 380746 633818 380982 634054
rect 380426 633498 380662 633734
rect 380746 633498 380982 633734
rect 380426 597818 380662 598054
rect 380746 597818 380982 598054
rect 380426 597498 380662 597734
rect 380746 597498 380982 597734
rect 380426 561818 380662 562054
rect 380746 561818 380982 562054
rect 380426 561498 380662 561734
rect 380746 561498 380982 561734
rect 380426 525818 380662 526054
rect 380746 525818 380982 526054
rect 380426 525498 380662 525734
rect 380746 525498 380982 525734
rect 380426 489818 380662 490054
rect 380746 489818 380982 490054
rect 380426 489498 380662 489734
rect 380746 489498 380982 489734
rect 380426 453818 380662 454054
rect 380746 453818 380982 454054
rect 380426 453498 380662 453734
rect 380746 453498 380982 453734
rect 380426 417818 380662 418054
rect 380746 417818 380982 418054
rect 380426 417498 380662 417734
rect 380746 417498 380982 417734
rect 380426 381818 380662 382054
rect 380746 381818 380982 382054
rect 380426 381498 380662 381734
rect 380746 381498 380982 381734
rect 380426 345818 380662 346054
rect 380746 345818 380982 346054
rect 380426 345498 380662 345734
rect 380746 345498 380982 345734
rect 380426 309818 380662 310054
rect 380746 309818 380982 310054
rect 380426 309498 380662 309734
rect 380746 309498 380982 309734
rect 384146 710362 384382 710598
rect 384466 710362 384702 710598
rect 384146 710042 384382 710278
rect 384466 710042 384702 710278
rect 384146 673538 384382 673774
rect 384466 673538 384702 673774
rect 384146 673218 384382 673454
rect 384466 673218 384702 673454
rect 384146 637538 384382 637774
rect 384466 637538 384702 637774
rect 384146 637218 384382 637454
rect 384466 637218 384702 637454
rect 384146 601538 384382 601774
rect 384466 601538 384702 601774
rect 384146 601218 384382 601454
rect 384466 601218 384702 601454
rect 384146 565538 384382 565774
rect 384466 565538 384702 565774
rect 384146 565218 384382 565454
rect 384466 565218 384702 565454
rect 384146 529538 384382 529774
rect 384466 529538 384702 529774
rect 384146 529218 384382 529454
rect 384466 529218 384702 529454
rect 384146 493538 384382 493774
rect 384466 493538 384702 493774
rect 384146 493218 384382 493454
rect 384466 493218 384702 493454
rect 384146 457538 384382 457774
rect 384466 457538 384702 457774
rect 384146 457218 384382 457454
rect 384466 457218 384702 457454
rect 384146 421538 384382 421774
rect 384466 421538 384702 421774
rect 384146 421218 384382 421454
rect 384466 421218 384702 421454
rect 384146 385538 384382 385774
rect 384466 385538 384702 385774
rect 384146 385218 384382 385454
rect 384466 385218 384702 385454
rect 384146 349538 384382 349774
rect 384466 349538 384702 349774
rect 384146 349218 384382 349454
rect 384466 349218 384702 349454
rect 384146 313538 384382 313774
rect 384466 313538 384702 313774
rect 384146 313218 384382 313454
rect 384466 313218 384702 313454
rect 380426 273818 380662 274054
rect 380746 273818 380982 274054
rect 380426 273498 380662 273734
rect 380746 273498 380982 273734
rect 380426 237818 380662 238054
rect 380746 237818 380982 238054
rect 380426 237498 380662 237734
rect 380746 237498 380982 237734
rect 380426 201818 380662 202054
rect 380746 201818 380982 202054
rect 380426 201498 380662 201734
rect 380746 201498 380982 201734
rect 380426 165818 380662 166054
rect 380746 165818 380982 166054
rect 380426 165498 380662 165734
rect 380746 165498 380982 165734
rect 380426 129818 380662 130054
rect 380746 129818 380982 130054
rect 380426 129498 380662 129734
rect 380746 129498 380982 129734
rect 380426 93818 380662 94054
rect 380746 93818 380982 94054
rect 380426 93498 380662 93734
rect 380746 93498 380982 93734
rect 380426 57818 380662 58054
rect 380746 57818 380982 58054
rect 380426 57498 380662 57734
rect 380746 57498 380982 57734
rect 384146 277538 384382 277774
rect 384466 277538 384702 277774
rect 384146 277218 384382 277454
rect 384466 277218 384702 277454
rect 384146 241538 384382 241774
rect 384466 241538 384702 241774
rect 384146 241218 384382 241454
rect 384466 241218 384702 241454
rect 384146 205538 384382 205774
rect 384466 205538 384702 205774
rect 384146 205218 384382 205454
rect 384466 205218 384702 205454
rect 384146 169538 384382 169774
rect 384466 169538 384702 169774
rect 384146 169218 384382 169454
rect 384466 169218 384702 169454
rect 384146 133538 384382 133774
rect 384466 133538 384702 133774
rect 384146 133218 384382 133454
rect 384466 133218 384702 133454
rect 384146 97538 384382 97774
rect 384466 97538 384702 97774
rect 384146 97218 384382 97454
rect 384466 97218 384702 97454
rect 387866 711322 388102 711558
rect 388186 711322 388422 711558
rect 387866 711002 388102 711238
rect 388186 711002 388422 711238
rect 387866 677258 388102 677494
rect 388186 677258 388422 677494
rect 387866 676938 388102 677174
rect 388186 676938 388422 677174
rect 387866 641258 388102 641494
rect 388186 641258 388422 641494
rect 387866 640938 388102 641174
rect 388186 640938 388422 641174
rect 387866 605258 388102 605494
rect 388186 605258 388422 605494
rect 387866 604938 388102 605174
rect 388186 604938 388422 605174
rect 387866 569258 388102 569494
rect 388186 569258 388422 569494
rect 387866 568938 388102 569174
rect 388186 568938 388422 569174
rect 387866 533258 388102 533494
rect 388186 533258 388422 533494
rect 387866 532938 388102 533174
rect 388186 532938 388422 533174
rect 387866 497258 388102 497494
rect 388186 497258 388422 497494
rect 387866 496938 388102 497174
rect 388186 496938 388422 497174
rect 387866 461258 388102 461494
rect 388186 461258 388422 461494
rect 387866 460938 388102 461174
rect 388186 460938 388422 461174
rect 387866 425258 388102 425494
rect 388186 425258 388422 425494
rect 387866 424938 388102 425174
rect 388186 424938 388422 425174
rect 387866 389258 388102 389494
rect 388186 389258 388422 389494
rect 387866 388938 388102 389174
rect 388186 388938 388422 389174
rect 387866 353258 388102 353494
rect 388186 353258 388422 353494
rect 387866 352938 388102 353174
rect 388186 352938 388422 353174
rect 387866 317258 388102 317494
rect 388186 317258 388422 317494
rect 387866 316938 388102 317174
rect 388186 316938 388422 317174
rect 387866 281258 388102 281494
rect 388186 281258 388422 281494
rect 387866 280938 388102 281174
rect 388186 280938 388422 281174
rect 387866 245258 388102 245494
rect 388186 245258 388422 245494
rect 387866 244938 388102 245174
rect 388186 244938 388422 245174
rect 387866 209258 388102 209494
rect 388186 209258 388422 209494
rect 387866 208938 388102 209174
rect 388186 208938 388422 209174
rect 387866 173258 388102 173494
rect 388186 173258 388422 173494
rect 387866 172938 388102 173174
rect 388186 172938 388422 173174
rect 387866 137258 388102 137494
rect 388186 137258 388422 137494
rect 387866 136938 388102 137174
rect 388186 136938 388422 137174
rect 387866 101258 388102 101494
rect 388186 101258 388422 101494
rect 387866 100938 388102 101174
rect 388186 100938 388422 101174
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 401546 705562 401782 705798
rect 401866 705562 402102 705798
rect 401546 705242 401782 705478
rect 401866 705242 402102 705478
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 405266 706522 405502 706758
rect 405586 706522 405822 706758
rect 405266 706202 405502 706438
rect 405586 706202 405822 706438
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 404459 327218 404695 327454
rect 404459 326898 404695 327134
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 408986 707482 409222 707718
rect 409306 707482 409542 707718
rect 408986 707162 409222 707398
rect 409306 707162 409542 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 407932 330938 408168 331174
rect 407932 330618 408168 330854
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 412706 708442 412942 708678
rect 413026 708442 413262 708678
rect 412706 708122 412942 708358
rect 413026 708122 413262 708358
rect 412706 666098 412942 666334
rect 413026 666098 413262 666334
rect 412706 665778 412942 666014
rect 413026 665778 413262 666014
rect 412706 630098 412942 630334
rect 413026 630098 413262 630334
rect 412706 629778 412942 630014
rect 413026 629778 413262 630014
rect 412706 594098 412942 594334
rect 413026 594098 413262 594334
rect 412706 593778 412942 594014
rect 413026 593778 413262 594014
rect 412706 558098 412942 558334
rect 413026 558098 413262 558334
rect 412706 557778 412942 558014
rect 413026 557778 413262 558014
rect 412706 522098 412942 522334
rect 413026 522098 413262 522334
rect 412706 521778 412942 522014
rect 413026 521778 413262 522014
rect 412706 486098 412942 486334
rect 413026 486098 413262 486334
rect 412706 485778 412942 486014
rect 413026 485778 413262 486014
rect 412706 450098 412942 450334
rect 413026 450098 413262 450334
rect 412706 449778 412942 450014
rect 413026 449778 413262 450014
rect 412706 414098 412942 414334
rect 413026 414098 413262 414334
rect 412706 413778 412942 414014
rect 413026 413778 413262 414014
rect 412706 378098 412942 378334
rect 413026 378098 413262 378334
rect 412706 377778 412942 378014
rect 413026 377778 413262 378014
rect 412706 342098 412942 342334
rect 413026 342098 413262 342334
rect 412706 341778 412942 342014
rect 413026 341778 413262 342014
rect 411405 327218 411641 327454
rect 411405 326898 411641 327134
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 416426 709402 416662 709638
rect 416746 709402 416982 709638
rect 416426 709082 416662 709318
rect 416746 709082 416982 709318
rect 416426 669818 416662 670054
rect 416746 669818 416982 670054
rect 416426 669498 416662 669734
rect 416746 669498 416982 669734
rect 416426 633818 416662 634054
rect 416746 633818 416982 634054
rect 416426 633498 416662 633734
rect 416746 633498 416982 633734
rect 416426 597818 416662 598054
rect 416746 597818 416982 598054
rect 416426 597498 416662 597734
rect 416746 597498 416982 597734
rect 416426 561818 416662 562054
rect 416746 561818 416982 562054
rect 416426 561498 416662 561734
rect 416746 561498 416982 561734
rect 416426 525818 416662 526054
rect 416746 525818 416982 526054
rect 416426 525498 416662 525734
rect 416746 525498 416982 525734
rect 416426 489818 416662 490054
rect 416746 489818 416982 490054
rect 416426 489498 416662 489734
rect 416746 489498 416982 489734
rect 416426 453818 416662 454054
rect 416746 453818 416982 454054
rect 416426 453498 416662 453734
rect 416746 453498 416982 453734
rect 416426 417818 416662 418054
rect 416746 417818 416982 418054
rect 416426 417498 416662 417734
rect 416746 417498 416982 417734
rect 416426 381818 416662 382054
rect 416746 381818 416982 382054
rect 416426 381498 416662 381734
rect 416746 381498 416982 381734
rect 416426 345818 416662 346054
rect 416746 345818 416982 346054
rect 416426 345498 416662 345734
rect 416746 345498 416982 345734
rect 414878 330938 415114 331174
rect 414878 330618 415114 330854
rect 412706 306098 412942 306334
rect 413026 306098 413262 306334
rect 412706 305778 412942 306014
rect 413026 305778 413262 306014
rect 412706 270098 412942 270334
rect 413026 270098 413262 270334
rect 412706 269778 412942 270014
rect 413026 269778 413262 270014
rect 412706 234098 412942 234334
rect 413026 234098 413262 234334
rect 412706 233778 412942 234014
rect 413026 233778 413262 234014
rect 412706 198098 412942 198334
rect 413026 198098 413262 198334
rect 412706 197778 412942 198014
rect 413026 197778 413262 198014
rect 412706 162098 412942 162334
rect 413026 162098 413262 162334
rect 412706 161778 412942 162014
rect 413026 161778 413262 162014
rect 420146 710362 420382 710598
rect 420466 710362 420702 710598
rect 420146 710042 420382 710278
rect 420466 710042 420702 710278
rect 420146 673538 420382 673774
rect 420466 673538 420702 673774
rect 420146 673218 420382 673454
rect 420466 673218 420702 673454
rect 420146 637538 420382 637774
rect 420466 637538 420702 637774
rect 420146 637218 420382 637454
rect 420466 637218 420702 637454
rect 420146 601538 420382 601774
rect 420466 601538 420702 601774
rect 420146 601218 420382 601454
rect 420466 601218 420702 601454
rect 420146 565538 420382 565774
rect 420466 565538 420702 565774
rect 420146 565218 420382 565454
rect 420466 565218 420702 565454
rect 420146 529538 420382 529774
rect 420466 529538 420702 529774
rect 420146 529218 420382 529454
rect 420466 529218 420702 529454
rect 420146 493538 420382 493774
rect 420466 493538 420702 493774
rect 420146 493218 420382 493454
rect 420466 493218 420702 493454
rect 420146 457538 420382 457774
rect 420466 457538 420702 457774
rect 420146 457218 420382 457454
rect 420466 457218 420702 457454
rect 423866 711322 424102 711558
rect 424186 711322 424422 711558
rect 423866 711002 424102 711238
rect 424186 711002 424422 711238
rect 423866 677258 424102 677494
rect 424186 677258 424422 677494
rect 423866 676938 424102 677174
rect 424186 676938 424422 677174
rect 423866 641258 424102 641494
rect 424186 641258 424422 641494
rect 423866 640938 424102 641174
rect 424186 640938 424422 641174
rect 423866 605258 424102 605494
rect 424186 605258 424422 605494
rect 423866 604938 424102 605174
rect 424186 604938 424422 605174
rect 423866 569258 424102 569494
rect 424186 569258 424422 569494
rect 423866 568938 424102 569174
rect 424186 568938 424422 569174
rect 423866 533258 424102 533494
rect 424186 533258 424422 533494
rect 423866 532938 424102 533174
rect 424186 532938 424422 533174
rect 423866 497258 424102 497494
rect 424186 497258 424422 497494
rect 423866 496938 424102 497174
rect 424186 496938 424422 497174
rect 423866 461258 424102 461494
rect 424186 461258 424422 461494
rect 423866 460938 424102 461174
rect 424186 460938 424422 461174
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 437546 705562 437782 705798
rect 437866 705562 438102 705798
rect 437546 705242 437782 705478
rect 437866 705242 438102 705478
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 441266 706522 441502 706758
rect 441586 706522 441822 706758
rect 441266 706202 441502 706438
rect 441586 706202 441822 706438
rect 444986 707482 445222 707718
rect 445306 707482 445542 707718
rect 444986 707162 445222 707398
rect 445306 707162 445542 707398
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 426666 438938 426902 439174
rect 426666 438618 426902 438854
rect 432347 438938 432583 439174
rect 432347 438618 432583 438854
rect 438028 438938 438264 439174
rect 438028 438618 438264 438854
rect 443709 438938 443945 439174
rect 443709 438618 443945 438854
rect 423826 435218 424062 435454
rect 423826 434898 424062 435134
rect 429507 435218 429743 435454
rect 429507 434898 429743 435134
rect 435188 435218 435424 435454
rect 435188 434898 435424 435134
rect 440869 435218 441105 435454
rect 440869 434898 441105 435134
rect 420146 421538 420382 421774
rect 420466 421538 420702 421774
rect 420146 421218 420382 421454
rect 420466 421218 420702 421454
rect 420146 385538 420382 385774
rect 420466 385538 420702 385774
rect 420146 385218 420382 385454
rect 420466 385218 420702 385454
rect 420146 349538 420382 349774
rect 420466 349538 420702 349774
rect 420146 349218 420382 349454
rect 420466 349218 420702 349454
rect 418351 327218 418587 327454
rect 418351 326898 418587 327134
rect 416426 309818 416662 310054
rect 416746 309818 416982 310054
rect 416426 309498 416662 309734
rect 416746 309498 416982 309734
rect 416426 273818 416662 274054
rect 416746 273818 416982 274054
rect 416426 273498 416662 273734
rect 416746 273498 416982 273734
rect 416426 237818 416662 238054
rect 416746 237818 416982 238054
rect 416426 237498 416662 237734
rect 416746 237498 416982 237734
rect 416426 201818 416662 202054
rect 416746 201818 416982 202054
rect 416426 201498 416662 201734
rect 416746 201498 416982 201734
rect 416426 165818 416662 166054
rect 416746 165818 416982 166054
rect 416426 165498 416662 165734
rect 416746 165498 416982 165734
rect 423866 389258 424102 389494
rect 424186 389258 424422 389494
rect 423866 388938 424102 389174
rect 424186 388938 424422 389174
rect 423866 353258 424102 353494
rect 424186 353258 424422 353494
rect 423866 352938 424102 353174
rect 424186 352938 424422 353174
rect 420146 313538 420382 313774
rect 420466 313538 420702 313774
rect 420146 313218 420382 313454
rect 420466 313218 420702 313454
rect 420146 277538 420382 277774
rect 420466 277538 420702 277774
rect 420146 277218 420382 277454
rect 420466 277218 420702 277454
rect 420146 241538 420382 241774
rect 420466 241538 420702 241774
rect 420146 241218 420382 241454
rect 420466 241218 420702 241454
rect 420146 205538 420382 205774
rect 420466 205538 420702 205774
rect 420146 205218 420382 205454
rect 420466 205218 420702 205454
rect 420146 169538 420382 169774
rect 420466 169538 420702 169774
rect 420146 169218 420382 169454
rect 420466 169218 420702 169454
rect 421824 330938 422060 331174
rect 421824 330618 422060 330854
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 425297 327218 425533 327454
rect 425297 326898 425533 327134
rect 423866 317258 424102 317494
rect 424186 317258 424422 317494
rect 423866 316938 424102 317174
rect 424186 316938 424422 317174
rect 423866 281258 424102 281494
rect 424186 281258 424422 281494
rect 423866 280938 424102 281174
rect 424186 280938 424422 281174
rect 423866 245258 424102 245494
rect 424186 245258 424422 245494
rect 423866 244938 424102 245174
rect 424186 244938 424422 245174
rect 423866 209258 424102 209494
rect 424186 209258 424422 209494
rect 423866 208938 424102 209174
rect 424186 208938 424422 209174
rect 423866 173258 424102 173494
rect 424186 173258 424422 173494
rect 423866 172938 424102 173174
rect 424186 172938 424422 173174
rect 428770 330938 429006 331174
rect 428770 330618 429006 330854
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 448706 708442 448942 708678
rect 449026 708442 449262 708678
rect 448706 708122 448942 708358
rect 449026 708122 449262 708358
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 452426 709402 452662 709638
rect 452746 709402 452982 709638
rect 452426 709082 452662 709318
rect 452746 709082 452982 709318
rect 448706 666098 448942 666334
rect 449026 666098 449262 666334
rect 448706 665778 448942 666014
rect 449026 665778 449262 666014
rect 448706 630098 448942 630334
rect 449026 630098 449262 630334
rect 448706 629778 448942 630014
rect 449026 629778 449262 630014
rect 448706 594098 448942 594334
rect 449026 594098 449262 594334
rect 448706 593778 448942 594014
rect 449026 593778 449262 594014
rect 448706 558098 448942 558334
rect 449026 558098 449262 558334
rect 448706 557778 448942 558014
rect 449026 557778 449262 558014
rect 448706 522098 448942 522334
rect 449026 522098 449262 522334
rect 448706 521778 448942 522014
rect 449026 521778 449262 522014
rect 448706 486098 448942 486334
rect 449026 486098 449262 486334
rect 448706 485778 448942 486014
rect 449026 485778 449262 486014
rect 448706 450098 448942 450334
rect 449026 450098 449262 450334
rect 448706 449778 448942 450014
rect 449026 449778 449262 450014
rect 448706 414098 448942 414334
rect 449026 414098 449262 414334
rect 448706 413778 448942 414014
rect 449026 413778 449262 414014
rect 448706 378098 448942 378334
rect 449026 378098 449262 378334
rect 448706 377778 448942 378014
rect 449026 377778 449262 378014
rect 448706 342098 448942 342334
rect 449026 342098 449262 342334
rect 448706 341778 448942 342014
rect 449026 341778 449262 342014
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 452426 669818 452662 670054
rect 452746 669818 452982 670054
rect 452426 669498 452662 669734
rect 452746 669498 452982 669734
rect 452426 633818 452662 634054
rect 452746 633818 452982 634054
rect 452426 633498 452662 633734
rect 452746 633498 452982 633734
rect 452426 597818 452662 598054
rect 452746 597818 452982 598054
rect 452426 597498 452662 597734
rect 452746 597498 452982 597734
rect 452426 561818 452662 562054
rect 452746 561818 452982 562054
rect 452426 561498 452662 561734
rect 452746 561498 452982 561734
rect 452426 525818 452662 526054
rect 452746 525818 452982 526054
rect 452426 525498 452662 525734
rect 452746 525498 452982 525734
rect 456146 710362 456382 710598
rect 456466 710362 456702 710598
rect 456146 710042 456382 710278
rect 456466 710042 456702 710278
rect 456146 673538 456382 673774
rect 456466 673538 456702 673774
rect 456146 673218 456382 673454
rect 456466 673218 456702 673454
rect 459866 711322 460102 711558
rect 460186 711322 460422 711558
rect 459866 711002 460102 711238
rect 460186 711002 460422 711238
rect 459866 677258 460102 677494
rect 460186 677258 460422 677494
rect 459866 676938 460102 677174
rect 460186 676938 460422 677174
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 473546 705562 473782 705798
rect 473866 705562 474102 705798
rect 473546 705242 473782 705478
rect 473866 705242 474102 705478
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 477266 706522 477502 706758
rect 477586 706522 477822 706758
rect 477266 706202 477502 706438
rect 477586 706202 477822 706438
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 480986 707482 481222 707718
rect 481306 707482 481542 707718
rect 480986 707162 481222 707398
rect 481306 707162 481542 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 488426 709402 488662 709638
rect 488746 709402 488982 709638
rect 488426 709082 488662 709318
rect 488746 709082 488982 709318
rect 488426 669818 488662 670054
rect 488746 669818 488982 670054
rect 488426 669498 488662 669734
rect 488746 669498 488982 669734
rect 492146 710362 492382 710598
rect 492466 710362 492702 710598
rect 492146 710042 492382 710278
rect 492466 710042 492702 710278
rect 492146 673538 492382 673774
rect 492466 673538 492702 673774
rect 492146 673218 492382 673454
rect 492466 673218 492702 673454
rect 495866 711322 496102 711558
rect 496186 711322 496422 711558
rect 495866 711002 496102 711238
rect 496186 711002 496422 711238
rect 495866 677258 496102 677494
rect 496186 677258 496422 677494
rect 495866 676938 496102 677174
rect 496186 676938 496422 677174
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 509546 705562 509782 705798
rect 509866 705562 510102 705798
rect 509546 705242 509782 705478
rect 509866 705242 510102 705478
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 513266 706522 513502 706758
rect 513586 706522 513822 706758
rect 513266 706202 513502 706438
rect 513586 706202 513822 706438
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 516986 707482 517222 707718
rect 517306 707482 517542 707718
rect 516986 707162 517222 707398
rect 517306 707162 517542 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 520706 708442 520942 708678
rect 521026 708442 521262 708678
rect 520706 708122 520942 708358
rect 521026 708122 521262 708358
rect 520706 666098 520942 666334
rect 521026 666098 521262 666334
rect 520706 665778 520942 666014
rect 521026 665778 521262 666014
rect 456146 637538 456382 637774
rect 456466 637538 456702 637774
rect 456146 637218 456382 637454
rect 456466 637218 456702 637454
rect 456146 601538 456382 601774
rect 456466 601538 456702 601774
rect 456146 601218 456382 601454
rect 456466 601218 456702 601454
rect 456146 565538 456382 565774
rect 456466 565538 456702 565774
rect 456146 565218 456382 565454
rect 456466 565218 456702 565454
rect 456146 529538 456382 529774
rect 456466 529538 456702 529774
rect 456146 529218 456382 529454
rect 456466 529218 456702 529454
rect 479610 654938 479846 655174
rect 479610 654618 479846 654854
rect 510330 654938 510566 655174
rect 510330 654618 510566 654854
rect 464250 651218 464486 651454
rect 464250 650898 464486 651134
rect 494970 651218 495206 651454
rect 494970 650898 495206 651134
rect 453424 510938 453660 511174
rect 453424 510618 453660 510854
rect 455862 510938 456098 511174
rect 455862 510618 456098 510854
rect 458300 510938 458536 511174
rect 458300 510618 458536 510854
rect 452205 507218 452441 507454
rect 452205 506898 452441 507134
rect 454643 507218 454879 507454
rect 454643 506898 454879 507134
rect 457081 507218 457317 507454
rect 457081 506898 457317 507134
rect 452426 489818 452662 490054
rect 452746 489818 452982 490054
rect 452426 489498 452662 489734
rect 452746 489498 452982 489734
rect 452426 453818 452662 454054
rect 452746 453818 452982 454054
rect 452426 453498 452662 453734
rect 452746 453498 452982 453734
rect 452426 417818 452662 418054
rect 452746 417818 452982 418054
rect 452426 417498 452662 417734
rect 452746 417498 452982 417734
rect 452426 381818 452662 382054
rect 452746 381818 452982 382054
rect 452426 381498 452662 381734
rect 452746 381498 452982 381734
rect 456146 493538 456382 493774
rect 456466 493538 456702 493774
rect 456146 493218 456382 493454
rect 456466 493218 456702 493454
rect 456146 457538 456382 457774
rect 456466 457538 456702 457774
rect 456146 457218 456382 457454
rect 456466 457218 456702 457454
rect 456146 421538 456382 421774
rect 456466 421538 456702 421774
rect 456146 421218 456382 421454
rect 456466 421218 456702 421454
rect 520706 630098 520942 630334
rect 521026 630098 521262 630334
rect 520706 629778 520942 630014
rect 521026 629778 521262 630014
rect 479610 618938 479846 619174
rect 479610 618618 479846 618854
rect 510330 618938 510566 619174
rect 510330 618618 510566 618854
rect 464250 615218 464486 615454
rect 464250 614898 464486 615134
rect 494970 615218 495206 615454
rect 494970 614898 495206 615134
rect 459866 569258 460102 569494
rect 460186 569258 460422 569494
rect 459866 568938 460102 569174
rect 460186 568938 460422 569174
rect 459866 533258 460102 533494
rect 460186 533258 460422 533494
rect 459866 532938 460102 533174
rect 460186 532938 460422 533174
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 460738 510938 460974 511174
rect 460738 510618 460974 510854
rect 459519 507218 459755 507454
rect 459519 506898 459755 507134
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 459866 497258 460102 497494
rect 460186 497258 460422 497494
rect 459866 496938 460102 497174
rect 460186 496938 460422 497174
rect 459866 461258 460102 461494
rect 460186 461258 460422 461494
rect 459866 460938 460102 461174
rect 460186 460938 460422 461174
rect 459866 425258 460102 425494
rect 460186 425258 460422 425494
rect 459866 424938 460102 425174
rect 460186 424938 460422 425174
rect 456146 385538 456382 385774
rect 456466 385538 456702 385774
rect 456146 385218 456382 385454
rect 456466 385218 456702 385454
rect 454250 363218 454486 363454
rect 454250 362898 454486 363134
rect 452426 345818 452662 346054
rect 452746 345818 452982 346054
rect 452426 345498 452662 345734
rect 452746 345498 452982 345734
rect 448706 306098 448942 306334
rect 449026 306098 449262 306334
rect 448706 305778 448942 306014
rect 449026 305778 449262 306014
rect 448706 270098 448942 270334
rect 449026 270098 449262 270334
rect 448706 269778 448942 270014
rect 449026 269778 449262 270014
rect 448706 234098 448942 234334
rect 449026 234098 449262 234334
rect 448706 233778 448942 234014
rect 449026 233778 449262 234014
rect 448706 198098 448942 198334
rect 449026 198098 449262 198334
rect 448706 197778 448942 198014
rect 449026 197778 449262 198014
rect 448706 162098 448942 162334
rect 449026 162098 449262 162334
rect 448706 161778 448942 162014
rect 449026 161778 449262 162014
rect 456146 349538 456382 349774
rect 456466 349538 456702 349774
rect 456146 349218 456382 349454
rect 456466 349218 456702 349454
rect 454250 327218 454486 327454
rect 454250 326898 454486 327134
rect 452426 309818 452662 310054
rect 452746 309818 452982 310054
rect 452426 309498 452662 309734
rect 452746 309498 452982 309734
rect 452426 273818 452662 274054
rect 452746 273818 452982 274054
rect 452426 273498 452662 273734
rect 452746 273498 452982 273734
rect 452426 237818 452662 238054
rect 452746 237818 452982 238054
rect 452426 237498 452662 237734
rect 452746 237498 452982 237734
rect 452426 201818 452662 202054
rect 452746 201818 452982 202054
rect 452426 201498 452662 201734
rect 452746 201498 452982 201734
rect 452426 165818 452662 166054
rect 452746 165818 452982 166054
rect 452426 165498 452662 165734
rect 452746 165498 452982 165734
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 429610 150938 429846 151174
rect 429610 150618 429846 150854
rect 414250 147218 414486 147454
rect 414250 146898 414486 147134
rect 444970 147218 445206 147454
rect 444970 146898 445206 147134
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 452426 129818 452662 130054
rect 452746 129818 452982 130054
rect 452426 129498 452662 129734
rect 452746 129498 452982 129734
rect 416426 93818 416662 94054
rect 416746 93818 416982 94054
rect 416426 93498 416662 93734
rect 416746 93498 416982 93734
rect 420146 97538 420382 97774
rect 420466 97538 420702 97774
rect 420146 97218 420382 97454
rect 420466 97218 420702 97454
rect 423866 101258 424102 101494
rect 424186 101258 424422 101494
rect 423866 100938 424102 101174
rect 424186 100938 424422 101174
rect 452426 93818 452662 94054
rect 452746 93818 452982 94054
rect 452426 93498 452662 93734
rect 452746 93498 452982 93734
rect 456146 313538 456382 313774
rect 456466 313538 456702 313774
rect 456146 313218 456382 313454
rect 456466 313218 456702 313454
rect 456146 277538 456382 277774
rect 456466 277538 456702 277774
rect 456146 277218 456382 277454
rect 456466 277218 456702 277454
rect 456146 241538 456382 241774
rect 456466 241538 456702 241774
rect 456146 241218 456382 241454
rect 456466 241218 456702 241454
rect 456146 205538 456382 205774
rect 456466 205538 456702 205774
rect 456146 205218 456382 205454
rect 456466 205218 456702 205454
rect 456146 169538 456382 169774
rect 456466 169538 456702 169774
rect 456146 169218 456382 169454
rect 456466 169218 456702 169454
rect 456146 133538 456382 133774
rect 456466 133538 456702 133774
rect 456146 133218 456382 133454
rect 456466 133218 456702 133454
rect 456146 97538 456382 97774
rect 456466 97538 456702 97774
rect 456146 97218 456382 97454
rect 456466 97218 456702 97454
rect 459866 389258 460102 389494
rect 460186 389258 460422 389494
rect 459866 388938 460102 389174
rect 460186 388938 460422 389174
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473458 435218 473694 435454
rect 473458 434898 473694 435134
rect 475930 438938 476166 439174
rect 475930 438618 476166 438854
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 478403 435218 478639 435454
rect 478403 434898 478639 435134
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 484706 594098 484942 594334
rect 485026 594098 485262 594334
rect 484706 593778 484942 594014
rect 485026 593778 485262 594014
rect 484706 558098 484942 558334
rect 485026 558098 485262 558334
rect 484706 557778 484942 558014
rect 485026 557778 485262 558014
rect 484706 522098 484942 522334
rect 485026 522098 485262 522334
rect 484706 521778 484942 522014
rect 485026 521778 485262 522014
rect 488426 597818 488662 598054
rect 488746 597818 488982 598054
rect 488426 597498 488662 597734
rect 488746 597498 488982 597734
rect 488426 561818 488662 562054
rect 488746 561818 488982 562054
rect 488426 561498 488662 561734
rect 488746 561498 488982 561734
rect 488426 525818 488662 526054
rect 488746 525818 488982 526054
rect 488426 525498 488662 525734
rect 488746 525498 488982 525734
rect 492146 565538 492382 565774
rect 492466 565538 492702 565774
rect 492146 565218 492382 565454
rect 492466 565218 492702 565454
rect 492146 529538 492382 529774
rect 492466 529538 492702 529774
rect 492146 529218 492382 529454
rect 492466 529218 492702 529454
rect 483424 510938 483660 511174
rect 483424 510618 483660 510854
rect 485862 510938 486098 511174
rect 485862 510618 486098 510854
rect 488300 510938 488536 511174
rect 488300 510618 488536 510854
rect 490738 510938 490974 511174
rect 490738 510618 490974 510854
rect 482205 507218 482441 507454
rect 482205 506898 482441 507134
rect 484643 507218 484879 507454
rect 484643 506898 484879 507134
rect 487081 507218 487317 507454
rect 487081 506898 487317 507134
rect 489519 507218 489755 507454
rect 489519 506898 489755 507134
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 484706 486098 484942 486334
rect 485026 486098 485262 486334
rect 484706 485778 484942 486014
rect 485026 485778 485262 486014
rect 488426 489818 488662 490054
rect 488746 489818 488982 490054
rect 488426 489498 488662 489734
rect 488746 489498 488982 489734
rect 484706 450098 484942 450334
rect 485026 450098 485262 450334
rect 484706 449778 484942 450014
rect 485026 449778 485262 450014
rect 480875 438938 481111 439174
rect 480875 438618 481111 438854
rect 483348 435218 483584 435454
rect 483348 434898 483584 435134
rect 485820 438938 486056 439174
rect 485820 438618 486056 438854
rect 484706 414098 484942 414334
rect 485026 414098 485262 414334
rect 484706 413778 484942 414014
rect 485026 413778 485262 414014
rect 488426 453771 488662 454007
rect 488746 453771 488982 454007
rect 492146 493538 492382 493774
rect 492466 493538 492702 493774
rect 492146 493218 492382 493454
rect 492466 493218 492702 493454
rect 492146 457538 492382 457774
rect 492466 457538 492702 457774
rect 492146 457218 492382 457454
rect 492466 457218 492702 457454
rect 490765 438938 491001 439174
rect 490765 438618 491001 438854
rect 488293 435218 488529 435454
rect 488293 434898 488529 435134
rect 492146 421538 492382 421774
rect 492466 421538 492702 421774
rect 492146 421218 492382 421454
rect 492466 421218 492702 421454
rect 495866 569258 496102 569494
rect 496186 569258 496422 569494
rect 495866 568938 496102 569174
rect 496186 568938 496422 569174
rect 495866 533258 496102 533494
rect 496186 533258 496422 533494
rect 495866 532938 496102 533174
rect 496186 532938 496422 533174
rect 495866 497258 496102 497494
rect 496186 497258 496422 497494
rect 495866 496938 496102 497174
rect 496186 496938 496422 497174
rect 495866 461258 496102 461494
rect 496186 461258 496422 461494
rect 495866 460938 496102 461174
rect 496186 460938 496422 461174
rect 495866 425258 496102 425494
rect 496186 425258 496422 425494
rect 495866 424938 496102 425174
rect 496186 424938 496422 425174
rect 495866 389258 496102 389494
rect 496186 389258 496422 389494
rect 495866 388938 496102 389174
rect 496186 388938 496422 389174
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 469610 366938 469846 367174
rect 469610 366618 469846 366854
rect 500330 366938 500566 367174
rect 500330 366618 500566 366854
rect 484970 363218 485206 363454
rect 484970 362898 485206 363134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 459866 353258 460102 353494
rect 460186 353258 460422 353494
rect 459866 352938 460102 353174
rect 460186 352938 460422 353174
rect 469610 330938 469846 331174
rect 469610 330618 469846 330854
rect 500330 330938 500566 331174
rect 500330 330618 500566 330854
rect 484970 327218 485206 327454
rect 484970 326898 485206 327134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 459866 317258 460102 317494
rect 460186 317258 460422 317494
rect 459866 316938 460102 317174
rect 460186 316938 460422 317174
rect 459866 281258 460102 281494
rect 460186 281258 460422 281494
rect 459866 280938 460102 281174
rect 460186 280938 460422 281174
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 484706 306098 484942 306334
rect 485026 306098 485262 306334
rect 484706 305778 484942 306014
rect 485026 305778 485262 306014
rect 484706 270098 484942 270334
rect 485026 270098 485262 270334
rect 484706 269778 484942 270014
rect 485026 269778 485262 270014
rect 488426 309818 488662 310054
rect 488746 309818 488982 310054
rect 488426 309498 488662 309734
rect 488746 309498 488982 309734
rect 488426 273818 488662 274054
rect 488746 273818 488982 274054
rect 488426 273498 488662 273734
rect 488746 273498 488982 273734
rect 492146 313538 492382 313774
rect 492466 313538 492702 313774
rect 492146 313218 492382 313454
rect 492466 313218 492702 313454
rect 492146 277538 492382 277774
rect 492466 277538 492702 277774
rect 492146 277218 492382 277454
rect 492466 277218 492702 277454
rect 495866 317258 496102 317494
rect 496186 317258 496422 317494
rect 495866 316938 496102 317174
rect 496186 316938 496422 317174
rect 495866 281258 496102 281494
rect 496186 281258 496422 281494
rect 495866 280938 496102 281174
rect 496186 280938 496422 281174
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 520706 594098 520942 594334
rect 521026 594098 521262 594334
rect 520706 593778 520942 594014
rect 521026 593778 521262 594014
rect 520706 558098 520942 558334
rect 521026 558098 521262 558334
rect 520706 557778 520942 558014
rect 521026 557778 521262 558014
rect 520706 522098 520942 522334
rect 521026 522098 521262 522334
rect 520706 521778 520942 522014
rect 521026 521778 521262 522014
rect 520706 486098 520942 486334
rect 521026 486098 521262 486334
rect 520706 485778 520942 486014
rect 521026 485778 521262 486014
rect 520706 450098 520942 450334
rect 521026 450098 521262 450334
rect 520706 449778 520942 450014
rect 521026 449778 521262 450014
rect 520706 414098 520942 414334
rect 521026 414098 521262 414334
rect 520706 413778 520942 414014
rect 521026 413778 521262 414014
rect 520706 378098 520942 378334
rect 521026 378098 521262 378334
rect 520706 377778 520942 378014
rect 521026 377778 521262 378014
rect 520706 342098 520942 342334
rect 521026 342098 521262 342334
rect 520706 341778 520942 342014
rect 521026 341778 521262 342014
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 520706 306098 520942 306334
rect 521026 306098 521262 306334
rect 520706 305778 520942 306014
rect 521026 305778 521262 306014
rect 520706 270098 520942 270334
rect 521026 270098 521262 270334
rect 520706 269778 520942 270014
rect 521026 269778 521262 270014
rect 524426 709402 524662 709638
rect 524746 709402 524982 709638
rect 524426 709082 524662 709318
rect 524746 709082 524982 709318
rect 528146 710362 528382 710598
rect 528466 710362 528702 710598
rect 528146 710042 528382 710278
rect 528466 710042 528702 710278
rect 524426 669818 524662 670054
rect 524746 669818 524982 670054
rect 524426 669498 524662 669734
rect 524746 669498 524982 669734
rect 525690 651218 525926 651454
rect 525690 650898 525926 651134
rect 524426 633818 524662 634054
rect 524746 633818 524982 634054
rect 524426 633498 524662 633734
rect 524746 633498 524982 633734
rect 525690 615218 525926 615454
rect 525690 614898 525926 615134
rect 524426 597818 524662 598054
rect 524746 597818 524982 598054
rect 524426 597498 524662 597734
rect 524746 597498 524982 597734
rect 524426 561818 524662 562054
rect 524746 561818 524982 562054
rect 524426 561498 524662 561734
rect 524746 561498 524982 561734
rect 524426 525818 524662 526054
rect 524746 525818 524982 526054
rect 524426 525498 524662 525734
rect 524746 525498 524982 525734
rect 524426 489818 524662 490054
rect 524746 489818 524982 490054
rect 524426 489498 524662 489734
rect 524746 489498 524982 489734
rect 524426 453818 524662 454054
rect 524746 453818 524982 454054
rect 524426 453498 524662 453734
rect 524746 453498 524982 453734
rect 525206 435218 525442 435454
rect 525206 434898 525442 435134
rect 524426 417818 524662 418054
rect 524746 417818 524982 418054
rect 524426 417498 524662 417734
rect 524746 417498 524982 417734
rect 524426 381818 524662 382054
rect 524746 381818 524982 382054
rect 524426 381498 524662 381734
rect 524746 381498 524982 381734
rect 524426 345818 524662 346054
rect 524746 345818 524982 346054
rect 524426 345498 524662 345734
rect 524746 345498 524982 345734
rect 528146 673538 528382 673774
rect 528466 673538 528702 673774
rect 528146 673218 528382 673454
rect 528466 673218 528702 673454
rect 528146 637538 528382 637774
rect 528466 637538 528702 637774
rect 528146 637218 528382 637454
rect 528466 637218 528702 637454
rect 528146 601538 528382 601774
rect 528466 601538 528702 601774
rect 528146 601218 528382 601454
rect 528466 601218 528702 601454
rect 528146 565538 528382 565774
rect 528466 565538 528702 565774
rect 528146 565218 528382 565454
rect 528466 565218 528702 565454
rect 528146 529538 528382 529774
rect 528466 529538 528702 529774
rect 528146 529218 528382 529454
rect 528466 529218 528702 529454
rect 528146 493538 528382 493774
rect 528466 493538 528702 493774
rect 528146 493218 528382 493454
rect 528466 493218 528702 493454
rect 528146 457538 528382 457774
rect 528466 457538 528702 457774
rect 528146 457218 528382 457454
rect 528466 457218 528702 457454
rect 531866 711322 532102 711558
rect 532186 711322 532422 711558
rect 531866 711002 532102 711238
rect 532186 711002 532422 711238
rect 531866 677258 532102 677494
rect 532186 677258 532422 677494
rect 531866 676938 532102 677174
rect 532186 676938 532422 677174
rect 531866 641258 532102 641494
rect 532186 641258 532422 641494
rect 531866 640938 532102 641174
rect 532186 640938 532422 641174
rect 531866 605258 532102 605494
rect 532186 605258 532422 605494
rect 531866 604938 532102 605174
rect 532186 604938 532422 605174
rect 531866 569258 532102 569494
rect 532186 569258 532422 569494
rect 531866 568938 532102 569174
rect 532186 568938 532422 569174
rect 531866 533258 532102 533494
rect 532186 533258 532422 533494
rect 531866 532938 532102 533174
rect 532186 532938 532422 533174
rect 531866 497258 532102 497494
rect 532186 497258 532422 497494
rect 531866 496938 532102 497174
rect 532186 496938 532422 497174
rect 531866 461258 532102 461494
rect 532186 461258 532422 461494
rect 531866 460938 532102 461174
rect 532186 460938 532422 461174
rect 529426 438938 529662 439174
rect 529426 438618 529662 438854
rect 528146 421538 528382 421774
rect 528466 421538 528702 421774
rect 528146 421218 528382 421454
rect 528466 421218 528702 421454
rect 528146 385538 528382 385774
rect 528466 385538 528702 385774
rect 528146 385218 528382 385454
rect 528466 385218 528702 385454
rect 528146 349538 528382 349774
rect 528466 349538 528702 349774
rect 528146 349218 528382 349454
rect 528466 349218 528702 349454
rect 524426 309818 524662 310054
rect 524746 309818 524982 310054
rect 524426 309498 524662 309734
rect 524746 309498 524982 309734
rect 524426 273818 524662 274054
rect 524746 273818 524982 274054
rect 524426 273498 524662 273734
rect 524746 273498 524982 273734
rect 528146 313538 528382 313774
rect 528466 313538 528702 313774
rect 528146 313218 528382 313454
rect 528466 313218 528702 313454
rect 528146 277538 528382 277774
rect 528466 277538 528702 277774
rect 528146 277218 528382 277454
rect 528466 277218 528702 277454
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 545546 705562 545782 705798
rect 545866 705562 546102 705798
rect 545546 705242 545782 705478
rect 545866 705242 546102 705478
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 537867 438938 538103 439174
rect 537867 438618 538103 438854
rect 549266 706522 549502 706758
rect 549586 706522 549822 706758
rect 549266 706202 549502 706438
rect 549586 706202 549822 706438
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 533647 435218 533883 435454
rect 533647 434898 533883 435134
rect 542088 435218 542324 435454
rect 542088 434898 542324 435134
rect 531866 425258 532102 425494
rect 532186 425258 532422 425494
rect 531866 424938 532102 425174
rect 532186 424938 532422 425174
rect 531866 389258 532102 389494
rect 532186 389258 532422 389494
rect 531866 388938 532102 389174
rect 532186 388938 532422 389174
rect 531866 353258 532102 353494
rect 532186 353258 532422 353494
rect 531866 352938 532102 353174
rect 532186 352938 532422 353174
rect 531866 317258 532102 317494
rect 532186 317258 532422 317494
rect 531866 316938 532102 317174
rect 532186 316938 532422 317174
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 531866 281258 532102 281494
rect 532186 281258 532422 281494
rect 531866 280938 532102 281174
rect 532186 280938 532422 281174
rect 479610 258938 479846 259174
rect 479610 258618 479846 258854
rect 510330 258938 510566 259174
rect 510330 258618 510566 258854
rect 464250 255218 464486 255454
rect 464250 254898 464486 255134
rect 494970 255218 495206 255454
rect 494970 254898 495206 255134
rect 525690 255218 525926 255454
rect 525690 254898 525926 255134
rect 459866 245258 460102 245494
rect 460186 245258 460422 245494
rect 459866 244938 460102 245174
rect 460186 244938 460422 245174
rect 531866 245258 532102 245494
rect 532186 245258 532422 245494
rect 531866 244938 532102 245174
rect 532186 244938 532422 245174
rect 479610 222938 479846 223174
rect 479610 222618 479846 222854
rect 510330 222938 510566 223174
rect 510330 222618 510566 222854
rect 464250 219218 464486 219454
rect 464250 218898 464486 219134
rect 494970 219218 495206 219454
rect 494970 218898 495206 219134
rect 525690 219218 525926 219454
rect 525690 218898 525926 219134
rect 459866 209258 460102 209494
rect 460186 209258 460422 209494
rect 459866 208938 460102 209174
rect 460186 208938 460422 209174
rect 531866 209258 532102 209494
rect 532186 209258 532422 209494
rect 531866 208938 532102 209174
rect 532186 208938 532422 209174
rect 459866 173258 460102 173494
rect 460186 173258 460422 173494
rect 459866 172938 460102 173174
rect 460186 172938 460422 173174
rect 459866 137258 460102 137494
rect 460186 137258 460422 137494
rect 459866 136938 460102 137174
rect 460186 136938 460422 137174
rect 459866 101258 460102 101494
rect 460186 101258 460422 101494
rect 459866 100938 460102 101174
rect 460186 100938 460422 101174
rect 405610 78938 405846 79174
rect 405610 78618 405846 78854
rect 436330 78938 436566 79174
rect 436330 78618 436566 78854
rect 390250 75218 390486 75454
rect 390250 74898 390486 75134
rect 420970 75218 421206 75454
rect 420970 74898 421206 75134
rect 451690 75218 451926 75454
rect 451690 74898 451926 75134
rect 384146 61538 384382 61774
rect 384466 61538 384702 61774
rect 384146 61218 384382 61454
rect 384466 61218 384702 61454
rect 380426 21818 380662 22054
rect 380746 21818 380982 22054
rect 380426 21498 380662 21734
rect 380746 21498 380982 21734
rect 380426 -5382 380662 -5146
rect 380746 -5382 380982 -5146
rect 380426 -5702 380662 -5466
rect 380746 -5702 380982 -5466
rect 459866 65258 460102 65494
rect 460186 65258 460422 65494
rect 459866 64938 460102 65174
rect 460186 64938 460422 65174
rect 405610 42938 405846 43174
rect 405610 42618 405846 42854
rect 436330 42938 436566 43174
rect 436330 42618 436566 42854
rect 390250 39218 390486 39454
rect 390250 38898 390486 39134
rect 420970 39218 421206 39454
rect 420970 38898 421206 39134
rect 451690 39218 451926 39454
rect 451690 38898 451926 39134
rect 384146 25538 384382 25774
rect 384466 25538 384702 25774
rect 384146 25218 384382 25454
rect 384466 25218 384702 25454
rect 384146 -6342 384382 -6106
rect 384466 -6342 384702 -6106
rect 384146 -6662 384382 -6426
rect 384466 -6662 384702 -6426
rect 387866 29258 388102 29494
rect 388186 29258 388422 29494
rect 387866 28938 388102 29174
rect 388186 28938 388422 29174
rect 387866 -7302 388102 -7066
rect 388186 -7302 388422 -7066
rect 387866 -7622 388102 -7386
rect 388186 -7622 388422 -7386
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -1542 401782 -1306
rect 401866 -1542 402102 -1306
rect 401546 -1862 401782 -1626
rect 401866 -1862 402102 -1626
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -2502 405502 -2266
rect 405586 -2502 405822 -2266
rect 405266 -2822 405502 -2586
rect 405586 -2822 405822 -2586
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 408986 -3462 409222 -3226
rect 409306 -3462 409542 -3226
rect 408986 -3782 409222 -3546
rect 409306 -3782 409542 -3546
rect 412706 18098 412942 18334
rect 413026 18098 413262 18334
rect 412706 17778 412942 18014
rect 413026 17778 413262 18014
rect 412706 -4422 412942 -4186
rect 413026 -4422 413262 -4186
rect 412706 -4742 412942 -4506
rect 413026 -4742 413262 -4506
rect 416426 21818 416662 22054
rect 416746 21818 416982 22054
rect 416426 21498 416662 21734
rect 416746 21498 416982 21734
rect 416426 -5382 416662 -5146
rect 416746 -5382 416982 -5146
rect 416426 -5702 416662 -5466
rect 416746 -5702 416982 -5466
rect 420146 25538 420382 25774
rect 420466 25538 420702 25774
rect 420146 25218 420382 25454
rect 420466 25218 420702 25454
rect 420146 -6342 420382 -6106
rect 420466 -6342 420702 -6106
rect 420146 -6662 420382 -6426
rect 420466 -6662 420702 -6426
rect 423866 29258 424102 29494
rect 424186 29258 424422 29494
rect 423866 28938 424102 29174
rect 424186 28938 424422 29174
rect 423866 -7302 424102 -7066
rect 424186 -7302 424422 -7066
rect 423866 -7622 424102 -7386
rect 424186 -7622 424422 -7386
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -1542 437782 -1306
rect 437866 -1542 438102 -1306
rect 437546 -1862 437782 -1626
rect 437866 -1862 438102 -1626
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -2502 441502 -2266
rect 441586 -2502 441822 -2266
rect 441266 -2822 441502 -2586
rect 441586 -2822 441822 -2586
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 444986 -3462 445222 -3226
rect 445306 -3462 445542 -3226
rect 444986 -3782 445222 -3546
rect 445306 -3782 445542 -3546
rect 448706 18098 448942 18334
rect 449026 18098 449262 18334
rect 448706 17778 448942 18014
rect 449026 17778 449262 18014
rect 448706 -4422 448942 -4186
rect 449026 -4422 449262 -4186
rect 448706 -4742 448942 -4506
rect 449026 -4742 449262 -4506
rect 452426 21818 452662 22054
rect 452746 21818 452982 22054
rect 452426 21498 452662 21734
rect 452746 21498 452982 21734
rect 452426 -5382 452662 -5146
rect 452746 -5382 452982 -5146
rect 452426 -5702 452662 -5466
rect 452746 -5702 452982 -5466
rect 456146 25538 456382 25774
rect 456466 25538 456702 25774
rect 456146 25218 456382 25454
rect 456466 25218 456702 25454
rect 456146 -6342 456382 -6106
rect 456466 -6342 456702 -6106
rect 456146 -6662 456382 -6426
rect 456466 -6662 456702 -6426
rect 459866 29258 460102 29494
rect 460186 29258 460422 29494
rect 459866 28938 460102 29174
rect 460186 28938 460422 29174
rect 459866 -7302 460102 -7066
rect 460186 -7302 460422 -7066
rect 459866 -7622 460102 -7386
rect 460186 -7622 460422 -7386
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -1542 473782 -1306
rect 473866 -1542 474102 -1306
rect 473546 -1862 473782 -1626
rect 473866 -1862 474102 -1626
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -2502 477502 -2266
rect 477586 -2502 477822 -2266
rect 477266 -2822 477502 -2586
rect 477586 -2822 477822 -2586
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 484706 198098 484942 198334
rect 485026 198098 485262 198334
rect 484706 197778 484942 198014
rect 485026 197778 485262 198014
rect 484706 162098 484942 162334
rect 485026 162098 485262 162334
rect 484706 161778 484942 162014
rect 485026 161778 485262 162014
rect 484706 126098 484942 126334
rect 485026 126098 485262 126334
rect 484706 125778 484942 126014
rect 485026 125778 485262 126014
rect 484250 111218 484486 111454
rect 484250 110898 484486 111134
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 480986 -3462 481222 -3226
rect 481306 -3462 481542 -3226
rect 480986 -3782 481222 -3546
rect 481306 -3782 481542 -3546
rect 484706 90098 484942 90334
rect 485026 90098 485262 90334
rect 484706 89778 484942 90014
rect 485026 89778 485262 90014
rect 484706 54098 484942 54334
rect 485026 54098 485262 54334
rect 484706 53778 484942 54014
rect 485026 53778 485262 54014
rect 484706 18098 484942 18334
rect 485026 18098 485262 18334
rect 484706 17778 484942 18014
rect 485026 17778 485262 18014
rect 484706 -4422 484942 -4186
rect 485026 -4422 485262 -4186
rect 484706 -4742 484942 -4506
rect 485026 -4742 485262 -4506
rect 488426 165818 488662 166054
rect 488746 165818 488982 166054
rect 488426 165498 488662 165734
rect 488746 165498 488982 165734
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 520706 198098 520942 198334
rect 521026 198098 521262 198334
rect 520706 197778 520942 198014
rect 521026 197778 521262 198014
rect 520706 162098 520942 162334
rect 521026 162098 521262 162334
rect 520706 161778 520942 162014
rect 521026 161778 521262 162014
rect 524426 165818 524662 166054
rect 524746 165818 524982 166054
rect 524426 165498 524662 165734
rect 524746 165498 524982 165734
rect 531866 173258 532102 173494
rect 532186 173258 532422 173494
rect 531866 172938 532102 173174
rect 532186 172938 532422 173174
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 488426 129818 488662 130054
rect 488746 129818 488982 130054
rect 488426 129498 488662 129734
rect 488746 129498 488982 129734
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 499610 114938 499846 115174
rect 499610 114618 499846 114854
rect 530330 114938 530566 115174
rect 530330 114618 530566 114854
rect 514970 111218 515206 111454
rect 514970 110898 515206 111134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 488426 93818 488662 94054
rect 488746 93818 488982 94054
rect 488426 93498 488662 93734
rect 488746 93498 488982 93734
rect 488426 57818 488662 58054
rect 488746 57818 488982 58054
rect 488426 57498 488662 57734
rect 488746 57498 488982 57734
rect 488426 21818 488662 22054
rect 488746 21818 488982 22054
rect 488426 21498 488662 21734
rect 488746 21498 488982 21734
rect 488426 -5382 488662 -5146
rect 488746 -5382 488982 -5146
rect 488426 -5702 488662 -5466
rect 488746 -5702 488982 -5466
rect 492146 61538 492382 61774
rect 492466 61538 492702 61774
rect 492146 61218 492382 61454
rect 492466 61218 492702 61454
rect 492146 25538 492382 25774
rect 492466 25538 492702 25774
rect 492146 25218 492382 25454
rect 492466 25218 492702 25454
rect 492146 -6342 492382 -6106
rect 492466 -6342 492702 -6106
rect 492146 -6662 492382 -6426
rect 492466 -6662 492702 -6426
rect 495866 65258 496102 65494
rect 496186 65258 496422 65494
rect 495866 64938 496102 65174
rect 496186 64938 496422 65174
rect 495866 29258 496102 29494
rect 496186 29258 496422 29494
rect 495866 28938 496102 29174
rect 496186 28938 496422 29174
rect 495866 -7302 496102 -7066
rect 496186 -7302 496422 -7066
rect 495866 -7622 496102 -7386
rect 496186 -7622 496422 -7386
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -1542 509782 -1306
rect 509866 -1542 510102 -1306
rect 509546 -1862 509782 -1626
rect 509866 -1862 510102 -1626
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -2502 513502 -2266
rect 513586 -2502 513822 -2266
rect 513266 -2822 513502 -2586
rect 513586 -2822 513822 -2586
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 516986 -3462 517222 -3226
rect 517306 -3462 517542 -3226
rect 516986 -3782 517222 -3546
rect 517306 -3782 517542 -3546
rect 520706 54098 520942 54334
rect 521026 54098 521262 54334
rect 520706 53778 520942 54014
rect 521026 53778 521262 54014
rect 520706 18098 520942 18334
rect 521026 18098 521262 18334
rect 520706 17778 520942 18014
rect 521026 17778 521262 18014
rect 520706 -4422 520942 -4186
rect 521026 -4422 521262 -4186
rect 520706 -4742 520942 -4506
rect 521026 -4742 521262 -4506
rect 524426 57818 524662 58054
rect 524746 57818 524982 58054
rect 524426 57498 524662 57734
rect 524746 57498 524982 57734
rect 524426 21818 524662 22054
rect 524746 21818 524982 22054
rect 524426 21498 524662 21734
rect 524746 21498 524982 21734
rect 524426 -5382 524662 -5146
rect 524746 -5382 524982 -5146
rect 524426 -5702 524662 -5466
rect 524746 -5702 524982 -5466
rect 528146 61538 528382 61774
rect 528466 61538 528702 61774
rect 528146 61218 528382 61454
rect 528466 61218 528702 61454
rect 528146 25538 528382 25774
rect 528466 25538 528702 25774
rect 528146 25218 528382 25454
rect 528466 25218 528702 25454
rect 528146 -6342 528382 -6106
rect 528466 -6342 528702 -6106
rect 528146 -6662 528382 -6426
rect 528466 -6662 528702 -6426
rect 531866 65258 532102 65494
rect 532186 65258 532422 65494
rect 531866 64938 532102 65174
rect 532186 64938 532422 65174
rect 531866 29258 532102 29494
rect 532186 29258 532422 29494
rect 531866 28938 532102 29174
rect 532186 28938 532422 29174
rect 531866 -7302 532102 -7066
rect 532186 -7302 532422 -7066
rect 531866 -7622 532102 -7386
rect 532186 -7622 532422 -7386
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 546308 438938 546544 439174
rect 546308 438618 546544 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 552986 707482 553222 707718
rect 553306 707482 553542 707718
rect 552986 707162 553222 707398
rect 553306 707162 553542 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 550529 435218 550765 435454
rect 550529 434898 550765 435134
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 556706 708442 556942 708678
rect 557026 708442 557262 708678
rect 556706 708122 556942 708358
rect 557026 708122 557262 708358
rect 560426 709402 560662 709638
rect 560746 709402 560982 709638
rect 560426 709082 560662 709318
rect 560746 709082 560982 709318
rect 556706 666098 556942 666334
rect 557026 666098 557262 666334
rect 556706 665778 556942 666014
rect 557026 665778 557262 666014
rect 556706 630098 556942 630334
rect 557026 630098 557262 630334
rect 556706 629778 556942 630014
rect 557026 629778 557262 630014
rect 556706 594098 556942 594334
rect 557026 594098 557262 594334
rect 556706 593778 556942 594014
rect 557026 593778 557262 594014
rect 556706 558098 556942 558334
rect 557026 558098 557262 558334
rect 556706 557778 556942 558014
rect 557026 557778 557262 558014
rect 556706 522098 556942 522334
rect 557026 522098 557262 522334
rect 556706 521778 556942 522014
rect 557026 521778 557262 522014
rect 556706 486098 556942 486334
rect 557026 486098 557262 486334
rect 556706 485778 556942 486014
rect 557026 485778 557262 486014
rect 556706 450098 556942 450334
rect 557026 450098 557262 450334
rect 556706 449778 556942 450014
rect 557026 449778 557262 450014
rect 554749 438938 554985 439174
rect 554749 438618 554985 438854
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 556706 414098 556942 414334
rect 557026 414098 557262 414334
rect 556706 413778 556942 414014
rect 557026 413778 557262 414014
rect 556706 378007 556942 378243
rect 557026 378007 557262 378243
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 554918 366938 555154 367174
rect 554918 366618 555154 366854
rect 558851 366938 559087 367174
rect 558851 366618 559087 366854
rect 552952 363218 553188 363454
rect 552952 362898 553188 363134
rect 556885 363218 557121 363454
rect 556885 362898 557121 363134
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 556706 342098 556942 342334
rect 557026 342098 557262 342334
rect 556706 341778 556942 342014
rect 557026 341778 557262 342014
rect 560426 669818 560662 670054
rect 560746 669818 560982 670054
rect 560426 669498 560662 669734
rect 560746 669498 560982 669734
rect 560426 633818 560662 634054
rect 560746 633818 560982 634054
rect 560426 633498 560662 633734
rect 560746 633498 560982 633734
rect 560426 597818 560662 598054
rect 560746 597818 560982 598054
rect 560426 597498 560662 597734
rect 560746 597498 560982 597734
rect 560426 561818 560662 562054
rect 560746 561818 560982 562054
rect 560426 561498 560662 561734
rect 560746 561498 560982 561734
rect 560426 525818 560662 526054
rect 560746 525818 560982 526054
rect 560426 525498 560662 525734
rect 560746 525498 560982 525734
rect 560426 489818 560662 490054
rect 560746 489818 560982 490054
rect 560426 489498 560662 489734
rect 560746 489498 560982 489734
rect 560426 453818 560662 454054
rect 560746 453818 560982 454054
rect 560426 453498 560662 453734
rect 560746 453498 560982 453734
rect 560426 417818 560662 418054
rect 560746 417818 560982 418054
rect 560426 417498 560662 417734
rect 560746 417498 560982 417734
rect 560426 381818 560662 382054
rect 560746 381818 560982 382054
rect 560426 381498 560662 381734
rect 560746 381498 560982 381734
rect 564146 710362 564382 710598
rect 564466 710362 564702 710598
rect 564146 710042 564382 710278
rect 564466 710042 564702 710278
rect 564146 673538 564382 673774
rect 564466 673538 564702 673774
rect 564146 673218 564382 673454
rect 564466 673218 564702 673454
rect 564146 637538 564382 637774
rect 564466 637538 564702 637774
rect 564146 637218 564382 637454
rect 564466 637218 564702 637454
rect 564146 601538 564382 601774
rect 564466 601538 564702 601774
rect 564146 601218 564382 601454
rect 564466 601218 564702 601454
rect 564146 565538 564382 565774
rect 564466 565538 564702 565774
rect 564146 565218 564382 565454
rect 564466 565218 564702 565454
rect 564146 529538 564382 529774
rect 564466 529538 564702 529774
rect 564146 529218 564382 529454
rect 564466 529218 564702 529454
rect 564146 493538 564382 493774
rect 564466 493538 564702 493774
rect 564146 493218 564382 493454
rect 564466 493218 564702 493454
rect 564146 457538 564382 457774
rect 564466 457538 564702 457774
rect 564146 457218 564382 457454
rect 564466 457218 564702 457454
rect 564146 421538 564382 421774
rect 564466 421538 564702 421774
rect 564146 421218 564382 421454
rect 564466 421218 564702 421454
rect 564146 385538 564382 385774
rect 564466 385538 564702 385774
rect 564146 385218 564382 385454
rect 564466 385218 564702 385454
rect 567866 711322 568102 711558
rect 568186 711322 568422 711558
rect 567866 711002 568102 711238
rect 568186 711002 568422 711238
rect 567866 677258 568102 677494
rect 568186 677258 568422 677494
rect 567866 676938 568102 677174
rect 568186 676938 568422 677174
rect 567866 641258 568102 641494
rect 568186 641258 568422 641494
rect 567866 640938 568102 641174
rect 568186 640938 568422 641174
rect 567866 605258 568102 605494
rect 568186 605258 568422 605494
rect 567866 604938 568102 605174
rect 568186 604938 568422 605174
rect 567866 569258 568102 569494
rect 568186 569258 568422 569494
rect 567866 568938 568102 569174
rect 568186 568938 568422 569174
rect 567866 533258 568102 533494
rect 568186 533258 568422 533494
rect 567866 532938 568102 533174
rect 568186 532938 568422 533174
rect 567866 497258 568102 497494
rect 568186 497258 568422 497494
rect 567866 496938 568102 497174
rect 568186 496938 568422 497174
rect 567866 461258 568102 461494
rect 568186 461258 568422 461494
rect 567866 460938 568102 461174
rect 568186 460938 568422 461174
rect 567866 425258 568102 425494
rect 568186 425258 568422 425494
rect 567866 424938 568102 425174
rect 568186 424938 568422 425174
rect 567866 389258 568102 389494
rect 568186 389258 568422 389494
rect 567866 388938 568102 389174
rect 568186 388938 568422 389174
rect 562784 366938 563020 367174
rect 562784 366618 563020 366854
rect 566717 366938 566953 367174
rect 566717 366618 566953 366854
rect 560818 363218 561054 363454
rect 560818 362898 561054 363134
rect 564751 363218 564987 363454
rect 564751 362898 564987 363134
rect 560426 345818 560662 346054
rect 560746 345818 560982 346054
rect 560426 345498 560662 345734
rect 560746 345498 560982 345734
rect 556706 306098 556942 306334
rect 557026 306098 557262 306334
rect 556706 305778 556942 306014
rect 557026 305778 557262 306014
rect 556706 270098 556942 270334
rect 557026 270098 557262 270334
rect 556706 269778 556942 270014
rect 557026 269778 557262 270014
rect 556706 234098 556942 234334
rect 557026 234098 557262 234334
rect 556706 233778 556942 234014
rect 557026 233778 557262 234014
rect 556706 198098 556942 198334
rect 557026 198098 557262 198334
rect 556706 197778 556942 198014
rect 557026 197778 557262 198014
rect 556706 162098 556942 162334
rect 557026 162098 557262 162334
rect 556706 161778 556942 162014
rect 557026 161778 557262 162014
rect 556706 126098 556942 126334
rect 557026 126098 557262 126334
rect 556706 125778 556942 126014
rect 557026 125778 557262 126014
rect 556706 90098 556942 90334
rect 557026 90098 557262 90334
rect 556706 89778 556942 90014
rect 557026 89778 557262 90014
rect 556706 54098 556942 54334
rect 557026 54098 557262 54334
rect 556706 53778 556942 54014
rect 557026 53778 557262 54014
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 545930 42938 546166 43174
rect 545930 42618 546166 42854
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 543458 39218 543694 39454
rect 543458 38898 543694 39134
rect 548403 39218 548639 39454
rect 548403 38898 548639 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -1542 545782 -1306
rect 545866 -1542 546102 -1306
rect 545546 -1862 545782 -1626
rect 545866 -1862 546102 -1626
rect 550875 42938 551111 43174
rect 550875 42618 551111 42854
rect 555820 42938 556056 43174
rect 555820 42618 556056 42854
rect 553348 39218 553584 39454
rect 553348 38898 553584 39134
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -2502 549502 -2266
rect 549586 -2502 549822 -2266
rect 549266 -2822 549502 -2586
rect 549586 -2822 549822 -2586
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 552986 -3462 553222 -3226
rect 553306 -3462 553542 -3226
rect 552986 -3782 553222 -3546
rect 553306 -3782 553542 -3546
rect 560426 309818 560662 310054
rect 560746 309818 560982 310054
rect 560426 309498 560662 309734
rect 560746 309498 560982 309734
rect 560426 273818 560662 274054
rect 560746 273818 560982 274054
rect 560426 273498 560662 273734
rect 560746 273498 560982 273734
rect 560426 237818 560662 238054
rect 560746 237818 560982 238054
rect 560426 237498 560662 237734
rect 560746 237498 560982 237734
rect 560426 201818 560662 202054
rect 560746 201818 560982 202054
rect 560426 201498 560662 201734
rect 560746 201498 560982 201734
rect 560426 165818 560662 166054
rect 560746 165818 560982 166054
rect 560426 165498 560662 165734
rect 560746 165498 560982 165734
rect 560426 129818 560662 130054
rect 560746 129818 560982 130054
rect 560426 129498 560662 129734
rect 560746 129498 560982 129734
rect 560426 93818 560662 94054
rect 560746 93818 560982 94054
rect 560426 93498 560662 93734
rect 560746 93498 560982 93734
rect 560426 57818 560662 58054
rect 560746 57818 560982 58054
rect 560426 57498 560662 57734
rect 560746 57498 560982 57734
rect 564146 349538 564382 349774
rect 564466 349538 564702 349774
rect 564146 349218 564382 349454
rect 564466 349218 564702 349454
rect 564146 313538 564382 313774
rect 564466 313538 564702 313774
rect 564146 313218 564382 313454
rect 564466 313218 564702 313454
rect 564146 277538 564382 277774
rect 564466 277538 564702 277774
rect 564146 277218 564382 277454
rect 564466 277218 564702 277454
rect 564146 241538 564382 241774
rect 564466 241538 564702 241774
rect 564146 241218 564382 241454
rect 564466 241218 564702 241454
rect 564146 205538 564382 205774
rect 564466 205538 564702 205774
rect 564146 205218 564382 205454
rect 564466 205218 564702 205454
rect 564146 169538 564382 169774
rect 564466 169538 564702 169774
rect 564146 169218 564382 169454
rect 564466 169218 564702 169454
rect 564146 133538 564382 133774
rect 564466 133538 564702 133774
rect 564146 133218 564382 133454
rect 564466 133218 564702 133454
rect 564146 97538 564382 97774
rect 564466 97538 564702 97774
rect 564146 97218 564382 97454
rect 564466 97218 564702 97454
rect 564146 61538 564382 61774
rect 564466 61538 564702 61774
rect 564146 61218 564382 61454
rect 564466 61218 564702 61454
rect 560765 42938 561001 43174
rect 560765 42618 561001 42854
rect 558293 39218 558529 39454
rect 558293 38898 558529 39134
rect 556706 18098 556942 18334
rect 557026 18098 557262 18334
rect 556706 17778 556942 18014
rect 557026 17778 557262 18014
rect 556706 -4422 556942 -4186
rect 557026 -4422 557262 -4186
rect 556706 -4742 556942 -4506
rect 557026 -4742 557262 -4506
rect 560426 21818 560662 22054
rect 560746 21818 560982 22054
rect 560426 21498 560662 21734
rect 560746 21498 560982 21734
rect 560426 -5382 560662 -5146
rect 560746 -5382 560982 -5146
rect 560426 -5702 560662 -5466
rect 560746 -5702 560982 -5466
rect 564146 25538 564382 25774
rect 564466 25538 564702 25774
rect 564146 25218 564382 25454
rect 564466 25218 564702 25454
rect 564146 -6342 564382 -6106
rect 564466 -6342 564702 -6106
rect 564146 -6662 564382 -6426
rect 564466 -6662 564702 -6426
rect 567866 353258 568102 353494
rect 568186 353258 568422 353494
rect 567866 352938 568102 353174
rect 568186 352938 568422 353174
rect 567866 317258 568102 317494
rect 568186 317258 568422 317494
rect 567866 316938 568102 317174
rect 568186 316938 568422 317174
rect 567866 281258 568102 281494
rect 568186 281258 568422 281494
rect 567866 280938 568102 281174
rect 568186 280938 568422 281174
rect 567866 245258 568102 245494
rect 568186 245258 568422 245494
rect 567866 244938 568102 245174
rect 568186 244938 568422 245174
rect 567866 209258 568102 209494
rect 568186 209258 568422 209494
rect 567866 208938 568102 209174
rect 568186 208938 568422 209174
rect 567866 173258 568102 173494
rect 568186 173258 568422 173494
rect 567866 172938 568102 173174
rect 568186 172938 568422 173174
rect 567866 137258 568102 137494
rect 568186 137258 568422 137494
rect 567866 136938 568102 137174
rect 568186 136938 568422 137174
rect 567866 101258 568102 101494
rect 568186 101258 568422 101494
rect 567866 100938 568102 101174
rect 568186 100938 568422 101174
rect 567866 65258 568102 65494
rect 568186 65258 568422 65494
rect 567866 64938 568102 65174
rect 568186 64938 568422 65174
rect 567866 29258 568102 29494
rect 568186 29258 568422 29494
rect 567866 28938 568102 29174
rect 568186 28938 568422 29174
rect 567866 -7302 568102 -7066
rect 568186 -7302 568422 -7066
rect 567866 -7622 568102 -7386
rect 568186 -7622 568422 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 581546 705562 581782 705798
rect 581866 705562 582102 705798
rect 581546 705242 581782 705478
rect 581866 705242 582102 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 690938 586538 691174
rect 586622 690938 586858 691174
rect 586302 690618 586538 690854
rect 586622 690618 586858 690854
rect 586302 654938 586538 655174
rect 586622 654938 586858 655174
rect 586302 654618 586538 654854
rect 586622 654618 586858 654854
rect 586302 618938 586538 619174
rect 586622 618938 586858 619174
rect 586302 618618 586538 618854
rect 586622 618618 586858 618854
rect 586302 582938 586538 583174
rect 586622 582938 586858 583174
rect 586302 582618 586538 582854
rect 586622 582618 586858 582854
rect 586302 546938 586538 547174
rect 586622 546938 586858 547174
rect 586302 546618 586538 546854
rect 586622 546618 586858 546854
rect 586302 510938 586538 511174
rect 586622 510938 586858 511174
rect 586302 510618 586538 510854
rect 586622 510618 586858 510854
rect 586302 474938 586538 475174
rect 586622 474938 586858 475174
rect 586302 474618 586538 474854
rect 586622 474618 586858 474854
rect 586302 438938 586538 439174
rect 586622 438938 586858 439174
rect 586302 438618 586538 438854
rect 586622 438618 586858 438854
rect 586302 402938 586538 403174
rect 586622 402938 586858 403174
rect 586302 402618 586538 402854
rect 586622 402618 586858 402854
rect 586302 366938 586538 367174
rect 586622 366938 586858 367174
rect 586302 366618 586538 366854
rect 586622 366618 586858 366854
rect 586302 330938 586538 331174
rect 586622 330938 586858 331174
rect 586302 330618 586538 330854
rect 586622 330618 586858 330854
rect 586302 294938 586538 295174
rect 586622 294938 586858 295174
rect 586302 294618 586538 294854
rect 586622 294618 586858 294854
rect 586302 258938 586538 259174
rect 586622 258938 586858 259174
rect 586302 258618 586538 258854
rect 586622 258618 586858 258854
rect 586302 222938 586538 223174
rect 586622 222938 586858 223174
rect 586302 222618 586538 222854
rect 586622 222618 586858 222854
rect 586302 186938 586538 187174
rect 586622 186938 586858 187174
rect 586302 186618 586538 186854
rect 586622 186618 586858 186854
rect 586302 150938 586538 151174
rect 586622 150938 586858 151174
rect 586302 150618 586538 150854
rect 586622 150618 586858 150854
rect 586302 114938 586538 115174
rect 586622 114938 586858 115174
rect 586302 114618 586538 114854
rect 586622 114618 586858 114854
rect 586302 78938 586538 79174
rect 586622 78938 586858 79174
rect 586302 78618 586538 78854
rect 586622 78618 586858 78854
rect 586302 42938 586538 43174
rect 586622 42938 586858 43174
rect 586302 42618 586538 42854
rect 586622 42618 586858 42854
rect 586302 6938 586538 7174
rect 586622 6938 586858 7174
rect 586302 6618 586538 6854
rect 586622 6618 586858 6854
rect 581546 -1542 581782 -1306
rect 581866 -1542 582102 -1306
rect 581546 -1862 581782 -1626
rect 581866 -1862 582102 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 694658 587498 694894
rect 587582 694658 587818 694894
rect 587262 694338 587498 694574
rect 587582 694338 587818 694574
rect 587262 658658 587498 658894
rect 587582 658658 587818 658894
rect 587262 658338 587498 658574
rect 587582 658338 587818 658574
rect 587262 622658 587498 622894
rect 587582 622658 587818 622894
rect 587262 622338 587498 622574
rect 587582 622338 587818 622574
rect 587262 586658 587498 586894
rect 587582 586658 587818 586894
rect 587262 586338 587498 586574
rect 587582 586338 587818 586574
rect 587262 550658 587498 550894
rect 587582 550658 587818 550894
rect 587262 550338 587498 550574
rect 587582 550338 587818 550574
rect 587262 514658 587498 514894
rect 587582 514658 587818 514894
rect 587262 514338 587498 514574
rect 587582 514338 587818 514574
rect 587262 478658 587498 478894
rect 587582 478658 587818 478894
rect 587262 478338 587498 478574
rect 587582 478338 587818 478574
rect 587262 442658 587498 442894
rect 587582 442658 587818 442894
rect 587262 442338 587498 442574
rect 587582 442338 587818 442574
rect 587262 406658 587498 406894
rect 587582 406658 587818 406894
rect 587262 406338 587498 406574
rect 587582 406338 587818 406574
rect 587262 370658 587498 370894
rect 587582 370658 587818 370894
rect 587262 370338 587498 370574
rect 587582 370338 587818 370574
rect 587262 334658 587498 334894
rect 587582 334658 587818 334894
rect 587262 334338 587498 334574
rect 587582 334338 587818 334574
rect 587262 298658 587498 298894
rect 587582 298658 587818 298894
rect 587262 298338 587498 298574
rect 587582 298338 587818 298574
rect 587262 262658 587498 262894
rect 587582 262658 587818 262894
rect 587262 262338 587498 262574
rect 587582 262338 587818 262574
rect 587262 226658 587498 226894
rect 587582 226658 587818 226894
rect 587262 226338 587498 226574
rect 587582 226338 587818 226574
rect 587262 190658 587498 190894
rect 587582 190658 587818 190894
rect 587262 190338 587498 190574
rect 587582 190338 587818 190574
rect 587262 154658 587498 154894
rect 587582 154658 587818 154894
rect 587262 154338 587498 154574
rect 587582 154338 587818 154574
rect 587262 118658 587498 118894
rect 587582 118658 587818 118894
rect 587262 118338 587498 118574
rect 587582 118338 587818 118574
rect 587262 82658 587498 82894
rect 587582 82658 587818 82894
rect 587262 82338 587498 82574
rect 587582 82338 587818 82574
rect 587262 46658 587498 46894
rect 587582 46658 587818 46894
rect 587262 46338 587498 46574
rect 587582 46338 587818 46574
rect 587262 10658 587498 10894
rect 587582 10658 587818 10894
rect 587262 10338 587498 10574
rect 587582 10338 587818 10574
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 698378 588458 698614
rect 588542 698378 588778 698614
rect 588222 698058 588458 698294
rect 588542 698058 588778 698294
rect 588222 662378 588458 662614
rect 588542 662378 588778 662614
rect 588222 662058 588458 662294
rect 588542 662058 588778 662294
rect 588222 626378 588458 626614
rect 588542 626378 588778 626614
rect 588222 626058 588458 626294
rect 588542 626058 588778 626294
rect 588222 590378 588458 590614
rect 588542 590378 588778 590614
rect 588222 590058 588458 590294
rect 588542 590058 588778 590294
rect 588222 554378 588458 554614
rect 588542 554378 588778 554614
rect 588222 554058 588458 554294
rect 588542 554058 588778 554294
rect 588222 518378 588458 518614
rect 588542 518378 588778 518614
rect 588222 518058 588458 518294
rect 588542 518058 588778 518294
rect 588222 482378 588458 482614
rect 588542 482378 588778 482614
rect 588222 482058 588458 482294
rect 588542 482058 588778 482294
rect 588222 446378 588458 446614
rect 588542 446378 588778 446614
rect 588222 446058 588458 446294
rect 588542 446058 588778 446294
rect 588222 410378 588458 410614
rect 588542 410378 588778 410614
rect 588222 410058 588458 410294
rect 588542 410058 588778 410294
rect 588222 374378 588458 374614
rect 588542 374378 588778 374614
rect 588222 374058 588458 374294
rect 588542 374058 588778 374294
rect 588222 338378 588458 338614
rect 588542 338378 588778 338614
rect 588222 338058 588458 338294
rect 588542 338058 588778 338294
rect 588222 302378 588458 302614
rect 588542 302378 588778 302614
rect 588222 302058 588458 302294
rect 588542 302058 588778 302294
rect 588222 266378 588458 266614
rect 588542 266378 588778 266614
rect 588222 266058 588458 266294
rect 588542 266058 588778 266294
rect 588222 230378 588458 230614
rect 588542 230378 588778 230614
rect 588222 230058 588458 230294
rect 588542 230058 588778 230294
rect 588222 194378 588458 194614
rect 588542 194378 588778 194614
rect 588222 194058 588458 194294
rect 588542 194058 588778 194294
rect 588222 158378 588458 158614
rect 588542 158378 588778 158614
rect 588222 158058 588458 158294
rect 588542 158058 588778 158294
rect 588222 122378 588458 122614
rect 588542 122378 588778 122614
rect 588222 122058 588458 122294
rect 588542 122058 588778 122294
rect 588222 86378 588458 86614
rect 588542 86378 588778 86614
rect 588222 86058 588458 86294
rect 588542 86058 588778 86294
rect 588222 50378 588458 50614
rect 588542 50378 588778 50614
rect 588222 50058 588458 50294
rect 588542 50058 588778 50294
rect 588222 14378 588458 14614
rect 588542 14378 588778 14614
rect 588222 14058 588458 14294
rect 588542 14058 588778 14294
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 666098 589418 666334
rect 589502 666098 589738 666334
rect 589182 665778 589418 666014
rect 589502 665778 589738 666014
rect 589182 630098 589418 630334
rect 589502 630098 589738 630334
rect 589182 629778 589418 630014
rect 589502 629778 589738 630014
rect 589182 594098 589418 594334
rect 589502 594098 589738 594334
rect 589182 593778 589418 594014
rect 589502 593778 589738 594014
rect 589182 558098 589418 558334
rect 589502 558098 589738 558334
rect 589182 557778 589418 558014
rect 589502 557778 589738 558014
rect 589182 522098 589418 522334
rect 589502 522098 589738 522334
rect 589182 521778 589418 522014
rect 589502 521778 589738 522014
rect 589182 486098 589418 486334
rect 589502 486098 589738 486334
rect 589182 485778 589418 486014
rect 589502 485778 589738 486014
rect 589182 450098 589418 450334
rect 589502 450098 589738 450334
rect 589182 449778 589418 450014
rect 589502 449778 589738 450014
rect 589182 414098 589418 414334
rect 589502 414098 589738 414334
rect 589182 413778 589418 414014
rect 589502 413778 589738 414014
rect 589182 378098 589418 378334
rect 589502 378098 589738 378334
rect 589182 377778 589418 378014
rect 589502 377778 589738 378014
rect 589182 342098 589418 342334
rect 589502 342098 589738 342334
rect 589182 341778 589418 342014
rect 589502 341778 589738 342014
rect 589182 306098 589418 306334
rect 589502 306098 589738 306334
rect 589182 305778 589418 306014
rect 589502 305778 589738 306014
rect 589182 270098 589418 270334
rect 589502 270098 589738 270334
rect 589182 269778 589418 270014
rect 589502 269778 589738 270014
rect 589182 234098 589418 234334
rect 589502 234098 589738 234334
rect 589182 233778 589418 234014
rect 589502 233778 589738 234014
rect 589182 198098 589418 198334
rect 589502 198098 589738 198334
rect 589182 197778 589418 198014
rect 589502 197778 589738 198014
rect 589182 162098 589418 162334
rect 589502 162098 589738 162334
rect 589182 161778 589418 162014
rect 589502 161778 589738 162014
rect 589182 126098 589418 126334
rect 589502 126098 589738 126334
rect 589182 125778 589418 126014
rect 589502 125778 589738 126014
rect 589182 90098 589418 90334
rect 589502 90098 589738 90334
rect 589182 89778 589418 90014
rect 589502 89778 589738 90014
rect 589182 54098 589418 54334
rect 589502 54098 589738 54334
rect 589182 53778 589418 54014
rect 589502 53778 589738 54014
rect 589182 18098 589418 18334
rect 589502 18098 589738 18334
rect 589182 17778 589418 18014
rect 589502 17778 589738 18014
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 669818 590378 670054
rect 590462 669818 590698 670054
rect 590142 669498 590378 669734
rect 590462 669498 590698 669734
rect 590142 633818 590378 634054
rect 590462 633818 590698 634054
rect 590142 633498 590378 633734
rect 590462 633498 590698 633734
rect 590142 597818 590378 598054
rect 590462 597818 590698 598054
rect 590142 597498 590378 597734
rect 590462 597498 590698 597734
rect 590142 561818 590378 562054
rect 590462 561818 590698 562054
rect 590142 561498 590378 561734
rect 590462 561498 590698 561734
rect 590142 525818 590378 526054
rect 590462 525818 590698 526054
rect 590142 525498 590378 525734
rect 590462 525498 590698 525734
rect 590142 489818 590378 490054
rect 590462 489818 590698 490054
rect 590142 489498 590378 489734
rect 590462 489498 590698 489734
rect 590142 453818 590378 454054
rect 590462 453818 590698 454054
rect 590142 453498 590378 453734
rect 590462 453498 590698 453734
rect 590142 417818 590378 418054
rect 590462 417818 590698 418054
rect 590142 417498 590378 417734
rect 590462 417498 590698 417734
rect 590142 381818 590378 382054
rect 590462 381818 590698 382054
rect 590142 381498 590378 381734
rect 590462 381498 590698 381734
rect 590142 345818 590378 346054
rect 590462 345818 590698 346054
rect 590142 345498 590378 345734
rect 590462 345498 590698 345734
rect 590142 309818 590378 310054
rect 590462 309818 590698 310054
rect 590142 309498 590378 309734
rect 590462 309498 590698 309734
rect 590142 273818 590378 274054
rect 590462 273818 590698 274054
rect 590142 273498 590378 273734
rect 590462 273498 590698 273734
rect 590142 237818 590378 238054
rect 590462 237818 590698 238054
rect 590142 237498 590378 237734
rect 590462 237498 590698 237734
rect 590142 201818 590378 202054
rect 590462 201818 590698 202054
rect 590142 201498 590378 201734
rect 590462 201498 590698 201734
rect 590142 165818 590378 166054
rect 590462 165818 590698 166054
rect 590142 165498 590378 165734
rect 590462 165498 590698 165734
rect 590142 129818 590378 130054
rect 590462 129818 590698 130054
rect 590142 129498 590378 129734
rect 590462 129498 590698 129734
rect 590142 93818 590378 94054
rect 590462 93818 590698 94054
rect 590142 93498 590378 93734
rect 590462 93498 590698 93734
rect 590142 57818 590378 58054
rect 590462 57818 590698 58054
rect 590142 57498 590378 57734
rect 590462 57498 590698 57734
rect 590142 21818 590378 22054
rect 590462 21818 590698 22054
rect 590142 21498 590378 21734
rect 590462 21498 590698 21734
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 673538 591338 673774
rect 591422 673538 591658 673774
rect 591102 673218 591338 673454
rect 591422 673218 591658 673454
rect 591102 637538 591338 637774
rect 591422 637538 591658 637774
rect 591102 637218 591338 637454
rect 591422 637218 591658 637454
rect 591102 601538 591338 601774
rect 591422 601538 591658 601774
rect 591102 601218 591338 601454
rect 591422 601218 591658 601454
rect 591102 565538 591338 565774
rect 591422 565538 591658 565774
rect 591102 565218 591338 565454
rect 591422 565218 591658 565454
rect 591102 529538 591338 529774
rect 591422 529538 591658 529774
rect 591102 529218 591338 529454
rect 591422 529218 591658 529454
rect 591102 493538 591338 493774
rect 591422 493538 591658 493774
rect 591102 493218 591338 493454
rect 591422 493218 591658 493454
rect 591102 457538 591338 457774
rect 591422 457538 591658 457774
rect 591102 457218 591338 457454
rect 591422 457218 591658 457454
rect 591102 421538 591338 421774
rect 591422 421538 591658 421774
rect 591102 421218 591338 421454
rect 591422 421218 591658 421454
rect 591102 385538 591338 385774
rect 591422 385538 591658 385774
rect 591102 385218 591338 385454
rect 591422 385218 591658 385454
rect 591102 349538 591338 349774
rect 591422 349538 591658 349774
rect 591102 349218 591338 349454
rect 591422 349218 591658 349454
rect 591102 313538 591338 313774
rect 591422 313538 591658 313774
rect 591102 313218 591338 313454
rect 591422 313218 591658 313454
rect 591102 277538 591338 277774
rect 591422 277538 591658 277774
rect 591102 277218 591338 277454
rect 591422 277218 591658 277454
rect 591102 241538 591338 241774
rect 591422 241538 591658 241774
rect 591102 241218 591338 241454
rect 591422 241218 591658 241454
rect 591102 205538 591338 205774
rect 591422 205538 591658 205774
rect 591102 205218 591338 205454
rect 591422 205218 591658 205454
rect 591102 169538 591338 169774
rect 591422 169538 591658 169774
rect 591102 169218 591338 169454
rect 591422 169218 591658 169454
rect 591102 133538 591338 133774
rect 591422 133538 591658 133774
rect 591102 133218 591338 133454
rect 591422 133218 591658 133454
rect 591102 97538 591338 97774
rect 591422 97538 591658 97774
rect 591102 97218 591338 97454
rect 591422 97218 591658 97454
rect 591102 61538 591338 61774
rect 591422 61538 591658 61774
rect 591102 61218 591338 61454
rect 591422 61218 591658 61454
rect 591102 25538 591338 25774
rect 591422 25538 591658 25774
rect 591102 25218 591338 25454
rect 591422 25218 591658 25454
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 677258 592298 677494
rect 592382 677258 592618 677494
rect 592062 676938 592298 677174
rect 592382 676938 592618 677174
rect 592062 641258 592298 641494
rect 592382 641258 592618 641494
rect 592062 640938 592298 641174
rect 592382 640938 592618 641174
rect 592062 605258 592298 605494
rect 592382 605258 592618 605494
rect 592062 604938 592298 605174
rect 592382 604938 592618 605174
rect 592062 569258 592298 569494
rect 592382 569258 592618 569494
rect 592062 568938 592298 569174
rect 592382 568938 592618 569174
rect 592062 533258 592298 533494
rect 592382 533258 592618 533494
rect 592062 532938 592298 533174
rect 592382 532938 592618 533174
rect 592062 497258 592298 497494
rect 592382 497258 592618 497494
rect 592062 496938 592298 497174
rect 592382 496938 592618 497174
rect 592062 461258 592298 461494
rect 592382 461258 592618 461494
rect 592062 460938 592298 461174
rect 592382 460938 592618 461174
rect 592062 425258 592298 425494
rect 592382 425258 592618 425494
rect 592062 424938 592298 425174
rect 592382 424938 592618 425174
rect 592062 389258 592298 389494
rect 592382 389258 592618 389494
rect 592062 388938 592298 389174
rect 592382 388938 592618 389174
rect 592062 353258 592298 353494
rect 592382 353258 592618 353494
rect 592062 352938 592298 353174
rect 592382 352938 592618 353174
rect 592062 317258 592298 317494
rect 592382 317258 592618 317494
rect 592062 316938 592298 317174
rect 592382 316938 592618 317174
rect 592062 281258 592298 281494
rect 592382 281258 592618 281494
rect 592062 280938 592298 281174
rect 592382 280938 592618 281174
rect 592062 245258 592298 245494
rect 592382 245258 592618 245494
rect 592062 244938 592298 245174
rect 592382 244938 592618 245174
rect 592062 209258 592298 209494
rect 592382 209258 592618 209494
rect 592062 208938 592298 209174
rect 592382 208938 592618 209174
rect 592062 173258 592298 173494
rect 592382 173258 592618 173494
rect 592062 172938 592298 173174
rect 592382 172938 592618 173174
rect 592062 137258 592298 137494
rect 592382 137258 592618 137494
rect 592062 136938 592298 137174
rect 592382 136938 592618 137174
rect 592062 101258 592298 101494
rect 592382 101258 592618 101494
rect 592062 100938 592298 101174
rect 592382 100938 592618 101174
rect 592062 65258 592298 65494
rect 592382 65258 592618 65494
rect 592062 64938 592298 65174
rect 592382 64938 592618 65174
rect 592062 29258 592298 29494
rect 592382 29258 592618 29494
rect 592062 28938 592298 29174
rect 592382 28938 592618 29174
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 348146 710598
rect 348382 710362 348466 710598
rect 348702 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 348146 710278
rect 348382 710042 348466 710278
rect 348702 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 344426 709638
rect 344662 709402 344746 709638
rect 344982 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 344426 709318
rect 344662 709082 344746 709318
rect 344982 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 520706 708678
rect 520942 708442 521026 708678
rect 521262 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 520706 708358
rect 520942 708122 521026 708358
rect 521262 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 592650 698294
rect -8726 698026 592650 698058
rect -8726 694894 592650 694926
rect -8726 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 592650 694894
rect -8726 694574 592650 694658
rect -8726 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 592650 694574
rect -8726 694306 592650 694338
rect -8726 691174 592650 691206
rect -8726 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 592650 691174
rect -8726 690854 592650 690938
rect -8726 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 592650 690854
rect -8726 690586 592650 690618
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 677494 592650 677526
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect -8726 677174 592650 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect -8726 676906 592650 676938
rect -8726 673774 592650 673806
rect -8726 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 348146 673774
rect 348382 673538 348466 673774
rect 348702 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 592650 673774
rect -8726 673454 592650 673538
rect -8726 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 348146 673454
rect 348382 673218 348466 673454
rect 348702 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 592650 673454
rect -8726 673186 592650 673218
rect -8726 670054 592650 670086
rect -8726 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 344426 670054
rect 344662 669818 344746 670054
rect 344982 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 592650 670054
rect -8726 669734 592650 669818
rect -8726 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 344426 669734
rect 344662 669498 344746 669734
rect 344982 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 592650 669734
rect -8726 669466 592650 669498
rect -8726 666334 592650 666366
rect -8726 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 520706 666334
rect 520942 666098 521026 666334
rect 521262 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 592650 666334
rect -8726 666014 592650 666098
rect -8726 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 520706 666014
rect 520942 665778 521026 666014
rect 521262 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 592650 666014
rect -8726 665746 592650 665778
rect -8726 662614 592650 662646
rect -8726 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 592650 662294
rect -8726 662026 592650 662058
rect -8726 658894 592650 658926
rect -8726 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 592650 658894
rect -8726 658574 592650 658658
rect -8726 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 592650 658574
rect -8726 658306 592650 658338
rect -8726 655174 592650 655206
rect -8726 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 39610 655174
rect 39846 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 70330 655174
rect 70566 654938 101050 655174
rect 101286 654938 131770 655174
rect 132006 654938 162490 655174
rect 162726 654938 193210 655174
rect 193446 654938 223930 655174
rect 224166 654938 254650 655174
rect 254886 654938 285370 655174
rect 285606 654938 316090 655174
rect 316326 654938 346810 655174
rect 347046 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 479610 655174
rect 479846 654938 510330 655174
rect 510566 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 592650 655174
rect -8726 654854 592650 654938
rect -8726 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 39610 654854
rect 39846 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 70330 654854
rect 70566 654618 101050 654854
rect 101286 654618 131770 654854
rect 132006 654618 162490 654854
rect 162726 654618 193210 654854
rect 193446 654618 223930 654854
rect 224166 654618 254650 654854
rect 254886 654618 285370 654854
rect 285606 654618 316090 654854
rect 316326 654618 346810 654854
rect 347046 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 479610 654854
rect 479846 654618 510330 654854
rect 510566 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 592650 654854
rect -8726 654586 592650 654618
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 24250 651454
rect 24486 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 54970 651454
rect 55206 651218 85690 651454
rect 85926 651218 116410 651454
rect 116646 651218 147130 651454
rect 147366 651218 177850 651454
rect 178086 651218 208570 651454
rect 208806 651218 239290 651454
rect 239526 651218 270010 651454
rect 270246 651218 300730 651454
rect 300966 651218 331450 651454
rect 331686 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 464250 651454
rect 464486 651218 494970 651454
rect 495206 651218 525690 651454
rect 525926 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 24250 651134
rect 24486 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 54970 651134
rect 55206 650898 85690 651134
rect 85926 650898 116410 651134
rect 116646 650898 147130 651134
rect 147366 650898 177850 651134
rect 178086 650898 208570 651134
rect 208806 650898 239290 651134
rect 239526 650898 270010 651134
rect 270246 650898 300730 651134
rect 300966 650898 331450 651134
rect 331686 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 464250 651134
rect 464486 650898 494970 651134
rect 495206 650898 525690 651134
rect 525926 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 641494 592650 641526
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 351866 641494
rect 352102 641258 352186 641494
rect 352422 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 423866 641494
rect 424102 641258 424186 641494
rect 424422 641258 531866 641494
rect 532102 641258 532186 641494
rect 532422 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect -8726 641174 592650 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 351866 641174
rect 352102 640938 352186 641174
rect 352422 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 423866 641174
rect 424102 640938 424186 641174
rect 424422 640938 531866 641174
rect 532102 640938 532186 641174
rect 532422 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect -8726 640906 592650 640938
rect -8726 637774 592650 637806
rect -8726 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 348146 637774
rect 348382 637538 348466 637774
rect 348702 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 420146 637774
rect 420382 637538 420466 637774
rect 420702 637538 456146 637774
rect 456382 637538 456466 637774
rect 456702 637538 528146 637774
rect 528382 637538 528466 637774
rect 528702 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 592650 637774
rect -8726 637454 592650 637538
rect -8726 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 348146 637454
rect 348382 637218 348466 637454
rect 348702 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 420146 637454
rect 420382 637218 420466 637454
rect 420702 637218 456146 637454
rect 456382 637218 456466 637454
rect 456702 637218 528146 637454
rect 528382 637218 528466 637454
rect 528702 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 592650 637454
rect -8726 637186 592650 637218
rect -8726 634054 592650 634086
rect -8726 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 344426 634054
rect 344662 633818 344746 634054
rect 344982 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 416426 634054
rect 416662 633818 416746 634054
rect 416982 633818 452426 634054
rect 452662 633818 452746 634054
rect 452982 633818 524426 634054
rect 524662 633818 524746 634054
rect 524982 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 592650 634054
rect -8726 633734 592650 633818
rect -8726 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 344426 633734
rect 344662 633498 344746 633734
rect 344982 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 416426 633734
rect 416662 633498 416746 633734
rect 416982 633498 452426 633734
rect 452662 633498 452746 633734
rect 452982 633498 524426 633734
rect 524662 633498 524746 633734
rect 524982 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 592650 633734
rect -8726 633466 592650 633498
rect -8726 630334 592650 630366
rect -8726 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 412706 630334
rect 412942 630098 413026 630334
rect 413262 630098 448706 630334
rect 448942 630098 449026 630334
rect 449262 630098 520706 630334
rect 520942 630098 521026 630334
rect 521262 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 592650 630334
rect -8726 630014 592650 630098
rect -8726 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 412706 630014
rect 412942 629778 413026 630014
rect 413262 629778 448706 630014
rect 448942 629778 449026 630014
rect 449262 629778 520706 630014
rect 520942 629778 521026 630014
rect 521262 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 592650 630014
rect -8726 629746 592650 629778
rect -8726 626614 592650 626646
rect -8726 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 592650 626294
rect -8726 626026 592650 626058
rect -8726 622894 592650 622926
rect -8726 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 592650 622894
rect -8726 622574 592650 622658
rect -8726 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 592650 622574
rect -8726 622306 592650 622338
rect -8726 619174 592650 619206
rect -8726 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 39610 619174
rect 39846 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 70330 619174
rect 70566 618938 101050 619174
rect 101286 618938 131770 619174
rect 132006 618938 162490 619174
rect 162726 618938 193210 619174
rect 193446 618938 223930 619174
rect 224166 618938 254650 619174
rect 254886 618938 285370 619174
rect 285606 618938 316090 619174
rect 316326 618938 346810 619174
rect 347046 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 479610 619174
rect 479846 618938 510330 619174
rect 510566 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 592650 619174
rect -8726 618854 592650 618938
rect -8726 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 39610 618854
rect 39846 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 70330 618854
rect 70566 618618 101050 618854
rect 101286 618618 131770 618854
rect 132006 618618 162490 618854
rect 162726 618618 193210 618854
rect 193446 618618 223930 618854
rect 224166 618618 254650 618854
rect 254886 618618 285370 618854
rect 285606 618618 316090 618854
rect 316326 618618 346810 618854
rect 347046 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 479610 618854
rect 479846 618618 510330 618854
rect 510566 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 592650 618854
rect -8726 618586 592650 618618
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 24250 615454
rect 24486 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 54970 615454
rect 55206 615218 85690 615454
rect 85926 615218 116410 615454
rect 116646 615218 147130 615454
rect 147366 615218 177850 615454
rect 178086 615218 208570 615454
rect 208806 615218 239290 615454
rect 239526 615218 270010 615454
rect 270246 615218 300730 615454
rect 300966 615218 331450 615454
rect 331686 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 464250 615454
rect 464486 615218 494970 615454
rect 495206 615218 525690 615454
rect 525926 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 24250 615134
rect 24486 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 54970 615134
rect 55206 614898 85690 615134
rect 85926 614898 116410 615134
rect 116646 614898 147130 615134
rect 147366 614898 177850 615134
rect 178086 614898 208570 615134
rect 208806 614898 239290 615134
rect 239526 614898 270010 615134
rect 270246 614898 300730 615134
rect 300966 614898 331450 615134
rect 331686 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 464250 615134
rect 464486 614898 494970 615134
rect 495206 614898 525690 615134
rect 525926 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 605494 592650 605526
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 351866 605494
rect 352102 605258 352186 605494
rect 352422 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 423866 605494
rect 424102 605258 424186 605494
rect 424422 605258 531866 605494
rect 532102 605258 532186 605494
rect 532422 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect -8726 605174 592650 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 351866 605174
rect 352102 604938 352186 605174
rect 352422 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 423866 605174
rect 424102 604938 424186 605174
rect 424422 604938 531866 605174
rect 532102 604938 532186 605174
rect 532422 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect -8726 604906 592650 604938
rect -8726 601774 592650 601806
rect -8726 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 348146 601774
rect 348382 601538 348466 601774
rect 348702 601538 384146 601774
rect 384382 601538 384466 601774
rect 384702 601538 420146 601774
rect 420382 601538 420466 601774
rect 420702 601538 456146 601774
rect 456382 601538 456466 601774
rect 456702 601538 528146 601774
rect 528382 601538 528466 601774
rect 528702 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 592650 601774
rect -8726 601454 592650 601538
rect -8726 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 348146 601454
rect 348382 601218 348466 601454
rect 348702 601218 384146 601454
rect 384382 601218 384466 601454
rect 384702 601218 420146 601454
rect 420382 601218 420466 601454
rect 420702 601218 456146 601454
rect 456382 601218 456466 601454
rect 456702 601218 528146 601454
rect 528382 601218 528466 601454
rect 528702 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 592650 601454
rect -8726 601186 592650 601218
rect -8726 598054 592650 598086
rect -8726 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 344426 598054
rect 344662 597818 344746 598054
rect 344982 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 416426 598054
rect 416662 597818 416746 598054
rect 416982 597818 452426 598054
rect 452662 597818 452746 598054
rect 452982 597818 488426 598054
rect 488662 597818 488746 598054
rect 488982 597818 524426 598054
rect 524662 597818 524746 598054
rect 524982 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 592650 598054
rect -8726 597734 592650 597818
rect -8726 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 344426 597734
rect 344662 597498 344746 597734
rect 344982 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 416426 597734
rect 416662 597498 416746 597734
rect 416982 597498 452426 597734
rect 452662 597498 452746 597734
rect 452982 597498 488426 597734
rect 488662 597498 488746 597734
rect 488982 597498 524426 597734
rect 524662 597498 524746 597734
rect 524982 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 592650 597734
rect -8726 597466 592650 597498
rect -8726 594334 592650 594366
rect -8726 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 412706 594334
rect 412942 594098 413026 594334
rect 413262 594098 448706 594334
rect 448942 594098 449026 594334
rect 449262 594098 484706 594334
rect 484942 594098 485026 594334
rect 485262 594098 520706 594334
rect 520942 594098 521026 594334
rect 521262 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 592650 594334
rect -8726 594014 592650 594098
rect -8726 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 412706 594014
rect 412942 593778 413026 594014
rect 413262 593778 448706 594014
rect 448942 593778 449026 594014
rect 449262 593778 484706 594014
rect 484942 593778 485026 594014
rect 485262 593778 520706 594014
rect 520942 593778 521026 594014
rect 521262 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 592650 594014
rect -8726 593746 592650 593778
rect -8726 590614 592650 590646
rect -8726 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 592650 590294
rect -8726 590026 592650 590058
rect -8726 586894 592650 586926
rect -8726 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 592650 586894
rect -8726 586574 592650 586658
rect -8726 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 592650 586574
rect -8726 586306 592650 586338
rect -8726 583174 592650 583206
rect -8726 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 39610 583174
rect 39846 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 70330 583174
rect 70566 582938 101050 583174
rect 101286 582938 131770 583174
rect 132006 582938 162490 583174
rect 162726 582938 193210 583174
rect 193446 582938 223930 583174
rect 224166 582938 254650 583174
rect 254886 582938 285370 583174
rect 285606 582938 316090 583174
rect 316326 582938 346810 583174
rect 347046 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 592650 583174
rect -8726 582854 592650 582938
rect -8726 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 39610 582854
rect 39846 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 70330 582854
rect 70566 582618 101050 582854
rect 101286 582618 131770 582854
rect 132006 582618 162490 582854
rect 162726 582618 193210 582854
rect 193446 582618 223930 582854
rect 224166 582618 254650 582854
rect 254886 582618 285370 582854
rect 285606 582618 316090 582854
rect 316326 582618 346810 582854
rect 347046 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 592650 582854
rect -8726 582586 592650 582618
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 24250 579454
rect 24486 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 54970 579454
rect 55206 579218 85690 579454
rect 85926 579218 116410 579454
rect 116646 579218 147130 579454
rect 147366 579218 177850 579454
rect 178086 579218 208570 579454
rect 208806 579218 239290 579454
rect 239526 579218 270010 579454
rect 270246 579218 300730 579454
rect 300966 579218 331450 579454
rect 331686 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 24250 579134
rect 24486 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 54970 579134
rect 55206 578898 85690 579134
rect 85926 578898 116410 579134
rect 116646 578898 147130 579134
rect 147366 578898 177850 579134
rect 178086 578898 208570 579134
rect 208806 578898 239290 579134
rect 239526 578898 270010 579134
rect 270246 578898 300730 579134
rect 300966 578898 331450 579134
rect 331686 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 569494 592650 569526
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 351866 569494
rect 352102 569258 352186 569494
rect 352422 569258 387866 569494
rect 388102 569258 388186 569494
rect 388422 569258 423866 569494
rect 424102 569258 424186 569494
rect 424422 569258 459866 569494
rect 460102 569258 460186 569494
rect 460422 569258 495866 569494
rect 496102 569258 496186 569494
rect 496422 569258 531866 569494
rect 532102 569258 532186 569494
rect 532422 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect -8726 569174 592650 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 351866 569174
rect 352102 568938 352186 569174
rect 352422 568938 387866 569174
rect 388102 568938 388186 569174
rect 388422 568938 423866 569174
rect 424102 568938 424186 569174
rect 424422 568938 459866 569174
rect 460102 568938 460186 569174
rect 460422 568938 495866 569174
rect 496102 568938 496186 569174
rect 496422 568938 531866 569174
rect 532102 568938 532186 569174
rect 532422 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect -8726 568906 592650 568938
rect -8726 565774 592650 565806
rect -8726 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 348146 565774
rect 348382 565538 348466 565774
rect 348702 565538 384146 565774
rect 384382 565538 384466 565774
rect 384702 565538 420146 565774
rect 420382 565538 420466 565774
rect 420702 565538 456146 565774
rect 456382 565538 456466 565774
rect 456702 565538 492146 565774
rect 492382 565538 492466 565774
rect 492702 565538 528146 565774
rect 528382 565538 528466 565774
rect 528702 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 592650 565774
rect -8726 565454 592650 565538
rect -8726 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 348146 565454
rect 348382 565218 348466 565454
rect 348702 565218 384146 565454
rect 384382 565218 384466 565454
rect 384702 565218 420146 565454
rect 420382 565218 420466 565454
rect 420702 565218 456146 565454
rect 456382 565218 456466 565454
rect 456702 565218 492146 565454
rect 492382 565218 492466 565454
rect 492702 565218 528146 565454
rect 528382 565218 528466 565454
rect 528702 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 592650 565454
rect -8726 565186 592650 565218
rect -8726 562054 592650 562086
rect -8726 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 344426 562054
rect 344662 561818 344746 562054
rect 344982 561818 380426 562054
rect 380662 561818 380746 562054
rect 380982 561818 416426 562054
rect 416662 561818 416746 562054
rect 416982 561818 452426 562054
rect 452662 561818 452746 562054
rect 452982 561818 488426 562054
rect 488662 561818 488746 562054
rect 488982 561818 524426 562054
rect 524662 561818 524746 562054
rect 524982 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 592650 562054
rect -8726 561734 592650 561818
rect -8726 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 344426 561734
rect 344662 561498 344746 561734
rect 344982 561498 380426 561734
rect 380662 561498 380746 561734
rect 380982 561498 416426 561734
rect 416662 561498 416746 561734
rect 416982 561498 452426 561734
rect 452662 561498 452746 561734
rect 452982 561498 488426 561734
rect 488662 561498 488746 561734
rect 488982 561498 524426 561734
rect 524662 561498 524746 561734
rect 524982 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 592650 561734
rect -8726 561466 592650 561498
rect -8726 558334 592650 558366
rect -8726 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 376706 558334
rect 376942 558098 377026 558334
rect 377262 558098 412706 558334
rect 412942 558098 413026 558334
rect 413262 558098 448706 558334
rect 448942 558098 449026 558334
rect 449262 558098 484706 558334
rect 484942 558098 485026 558334
rect 485262 558098 520706 558334
rect 520942 558098 521026 558334
rect 521262 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 592650 558334
rect -8726 558014 592650 558098
rect -8726 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 376706 558014
rect 376942 557778 377026 558014
rect 377262 557778 412706 558014
rect 412942 557778 413026 558014
rect 413262 557778 448706 558014
rect 448942 557778 449026 558014
rect 449262 557778 484706 558014
rect 484942 557778 485026 558014
rect 485262 557778 520706 558014
rect 520942 557778 521026 558014
rect 521262 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 592650 558014
rect -8726 557746 592650 557778
rect -8726 554614 592650 554646
rect -8726 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 592650 554294
rect -8726 554026 592650 554058
rect -8726 550894 592650 550926
rect -8726 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 592650 550894
rect -8726 550574 592650 550658
rect -8726 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 592650 550574
rect -8726 550306 592650 550338
rect -8726 547174 592650 547206
rect -8726 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 39610 547174
rect 39846 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 70330 547174
rect 70566 546938 101050 547174
rect 101286 546938 131770 547174
rect 132006 546938 162490 547174
rect 162726 546938 193210 547174
rect 193446 546938 223930 547174
rect 224166 546938 254650 547174
rect 254886 546938 285370 547174
rect 285606 546938 316090 547174
rect 316326 546938 346810 547174
rect 347046 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 592650 547174
rect -8726 546854 592650 546938
rect -8726 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 39610 546854
rect 39846 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 70330 546854
rect 70566 546618 101050 546854
rect 101286 546618 131770 546854
rect 132006 546618 162490 546854
rect 162726 546618 193210 546854
rect 193446 546618 223930 546854
rect 224166 546618 254650 546854
rect 254886 546618 285370 546854
rect 285606 546618 316090 546854
rect 316326 546618 346810 546854
rect 347046 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 592650 546854
rect -8726 546586 592650 546618
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 24250 543454
rect 24486 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 54970 543454
rect 55206 543218 85690 543454
rect 85926 543218 116410 543454
rect 116646 543218 147130 543454
rect 147366 543218 177850 543454
rect 178086 543218 208570 543454
rect 208806 543218 239290 543454
rect 239526 543218 270010 543454
rect 270246 543218 300730 543454
rect 300966 543218 331450 543454
rect 331686 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 24250 543134
rect 24486 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 54970 543134
rect 55206 542898 85690 543134
rect 85926 542898 116410 543134
rect 116646 542898 147130 543134
rect 147366 542898 177850 543134
rect 178086 542898 208570 543134
rect 208806 542898 239290 543134
rect 239526 542898 270010 543134
rect 270246 542898 300730 543134
rect 300966 542898 331450 543134
rect 331686 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 533494 592650 533526
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 351866 533494
rect 352102 533258 352186 533494
rect 352422 533258 387866 533494
rect 388102 533258 388186 533494
rect 388422 533258 423866 533494
rect 424102 533258 424186 533494
rect 424422 533258 459866 533494
rect 460102 533258 460186 533494
rect 460422 533258 495866 533494
rect 496102 533258 496186 533494
rect 496422 533258 531866 533494
rect 532102 533258 532186 533494
rect 532422 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect -8726 533174 592650 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 351866 533174
rect 352102 532938 352186 533174
rect 352422 532938 387866 533174
rect 388102 532938 388186 533174
rect 388422 532938 423866 533174
rect 424102 532938 424186 533174
rect 424422 532938 459866 533174
rect 460102 532938 460186 533174
rect 460422 532938 495866 533174
rect 496102 532938 496186 533174
rect 496422 532938 531866 533174
rect 532102 532938 532186 533174
rect 532422 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect -8726 532906 592650 532938
rect -8726 529774 592650 529806
rect -8726 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 348146 529774
rect 348382 529538 348466 529774
rect 348702 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 420146 529774
rect 420382 529538 420466 529774
rect 420702 529538 456146 529774
rect 456382 529538 456466 529774
rect 456702 529538 492146 529774
rect 492382 529538 492466 529774
rect 492702 529538 528146 529774
rect 528382 529538 528466 529774
rect 528702 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 592650 529774
rect -8726 529454 592650 529538
rect -8726 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 348146 529454
rect 348382 529218 348466 529454
rect 348702 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 420146 529454
rect 420382 529218 420466 529454
rect 420702 529218 456146 529454
rect 456382 529218 456466 529454
rect 456702 529218 492146 529454
rect 492382 529218 492466 529454
rect 492702 529218 528146 529454
rect 528382 529218 528466 529454
rect 528702 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 592650 529454
rect -8726 529186 592650 529218
rect -8726 526054 592650 526086
rect -8726 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 344426 526054
rect 344662 525818 344746 526054
rect 344982 525818 380426 526054
rect 380662 525818 380746 526054
rect 380982 525818 416426 526054
rect 416662 525818 416746 526054
rect 416982 525818 452426 526054
rect 452662 525818 452746 526054
rect 452982 525818 488426 526054
rect 488662 525818 488746 526054
rect 488982 525818 524426 526054
rect 524662 525818 524746 526054
rect 524982 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 592650 526054
rect -8726 525734 592650 525818
rect -8726 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 344426 525734
rect 344662 525498 344746 525734
rect 344982 525498 380426 525734
rect 380662 525498 380746 525734
rect 380982 525498 416426 525734
rect 416662 525498 416746 525734
rect 416982 525498 452426 525734
rect 452662 525498 452746 525734
rect 452982 525498 488426 525734
rect 488662 525498 488746 525734
rect 488982 525498 524426 525734
rect 524662 525498 524746 525734
rect 524982 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 592650 525734
rect -8726 525466 592650 525498
rect -8726 522334 592650 522366
rect -8726 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 376706 522334
rect 376942 522098 377026 522334
rect 377262 522098 412706 522334
rect 412942 522098 413026 522334
rect 413262 522098 448706 522334
rect 448942 522098 449026 522334
rect 449262 522098 484706 522334
rect 484942 522098 485026 522334
rect 485262 522098 520706 522334
rect 520942 522098 521026 522334
rect 521262 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 592650 522334
rect -8726 522014 592650 522098
rect -8726 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 376706 522014
rect 376942 521778 377026 522014
rect 377262 521778 412706 522014
rect 412942 521778 413026 522014
rect 413262 521778 448706 522014
rect 448942 521778 449026 522014
rect 449262 521778 484706 522014
rect 484942 521778 485026 522014
rect 485262 521778 520706 522014
rect 520942 521778 521026 522014
rect 521262 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 592650 522014
rect -8726 521746 592650 521778
rect -8726 518614 592650 518646
rect -8726 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 592650 518294
rect -8726 518026 592650 518058
rect -8726 514894 592650 514926
rect -8726 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 592650 514894
rect -8726 514574 592650 514658
rect -8726 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 592650 514574
rect -8726 514306 592650 514338
rect -8726 511174 592650 511206
rect -8726 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 39610 511174
rect 39846 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 70330 511174
rect 70566 510938 101050 511174
rect 101286 510938 131770 511174
rect 132006 510938 162490 511174
rect 162726 510938 193210 511174
rect 193446 510938 223930 511174
rect 224166 510938 254650 511174
rect 254886 510938 285370 511174
rect 285606 510938 316090 511174
rect 316326 510938 346810 511174
rect 347046 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 453424 511174
rect 453660 510938 455862 511174
rect 456098 510938 458300 511174
rect 458536 510938 460738 511174
rect 460974 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 483424 511174
rect 483660 510938 485862 511174
rect 486098 510938 488300 511174
rect 488536 510938 490738 511174
rect 490974 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 592650 511174
rect -8726 510854 592650 510938
rect -8726 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 39610 510854
rect 39846 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 70330 510854
rect 70566 510618 101050 510854
rect 101286 510618 131770 510854
rect 132006 510618 162490 510854
rect 162726 510618 193210 510854
rect 193446 510618 223930 510854
rect 224166 510618 254650 510854
rect 254886 510618 285370 510854
rect 285606 510618 316090 510854
rect 316326 510618 346810 510854
rect 347046 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 453424 510854
rect 453660 510618 455862 510854
rect 456098 510618 458300 510854
rect 458536 510618 460738 510854
rect 460974 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 483424 510854
rect 483660 510618 485862 510854
rect 486098 510618 488300 510854
rect 488536 510618 490738 510854
rect 490974 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 592650 510854
rect -8726 510586 592650 510618
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 24250 507454
rect 24486 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 54970 507454
rect 55206 507218 85690 507454
rect 85926 507218 116410 507454
rect 116646 507218 147130 507454
rect 147366 507218 177850 507454
rect 178086 507218 208570 507454
rect 208806 507218 239290 507454
rect 239526 507218 270010 507454
rect 270246 507218 300730 507454
rect 300966 507218 331450 507454
rect 331686 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 452205 507454
rect 452441 507218 454643 507454
rect 454879 507218 457081 507454
rect 457317 507218 459519 507454
rect 459755 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 482205 507454
rect 482441 507218 484643 507454
rect 484879 507218 487081 507454
rect 487317 507218 489519 507454
rect 489755 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 24250 507134
rect 24486 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 54970 507134
rect 55206 506898 85690 507134
rect 85926 506898 116410 507134
rect 116646 506898 147130 507134
rect 147366 506898 177850 507134
rect 178086 506898 208570 507134
rect 208806 506898 239290 507134
rect 239526 506898 270010 507134
rect 270246 506898 300730 507134
rect 300966 506898 331450 507134
rect 331686 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 452205 507134
rect 452441 506898 454643 507134
rect 454879 506898 457081 507134
rect 457317 506898 459519 507134
rect 459755 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 482205 507134
rect 482441 506898 484643 507134
rect 484879 506898 487081 507134
rect 487317 506898 489519 507134
rect 489755 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 497494 592650 497526
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 351866 497494
rect 352102 497258 352186 497494
rect 352422 497258 387866 497494
rect 388102 497258 388186 497494
rect 388422 497258 423866 497494
rect 424102 497258 424186 497494
rect 424422 497258 459866 497494
rect 460102 497258 460186 497494
rect 460422 497258 495866 497494
rect 496102 497258 496186 497494
rect 496422 497258 531866 497494
rect 532102 497258 532186 497494
rect 532422 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect -8726 497174 592650 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 351866 497174
rect 352102 496938 352186 497174
rect 352422 496938 387866 497174
rect 388102 496938 388186 497174
rect 388422 496938 423866 497174
rect 424102 496938 424186 497174
rect 424422 496938 459866 497174
rect 460102 496938 460186 497174
rect 460422 496938 495866 497174
rect 496102 496938 496186 497174
rect 496422 496938 531866 497174
rect 532102 496938 532186 497174
rect 532422 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect -8726 496906 592650 496938
rect -8726 493774 592650 493806
rect -8726 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 348146 493774
rect 348382 493538 348466 493774
rect 348702 493538 384146 493774
rect 384382 493538 384466 493774
rect 384702 493538 420146 493774
rect 420382 493538 420466 493774
rect 420702 493538 456146 493774
rect 456382 493538 456466 493774
rect 456702 493538 492146 493774
rect 492382 493538 492466 493774
rect 492702 493538 528146 493774
rect 528382 493538 528466 493774
rect 528702 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 592650 493774
rect -8726 493454 592650 493538
rect -8726 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 348146 493454
rect 348382 493218 348466 493454
rect 348702 493218 384146 493454
rect 384382 493218 384466 493454
rect 384702 493218 420146 493454
rect 420382 493218 420466 493454
rect 420702 493218 456146 493454
rect 456382 493218 456466 493454
rect 456702 493218 492146 493454
rect 492382 493218 492466 493454
rect 492702 493218 528146 493454
rect 528382 493218 528466 493454
rect 528702 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 592650 493454
rect -8726 493186 592650 493218
rect -8726 490054 592650 490086
rect -8726 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 344426 490054
rect 344662 489818 344746 490054
rect 344982 489818 380426 490054
rect 380662 489818 380746 490054
rect 380982 489818 416426 490054
rect 416662 489818 416746 490054
rect 416982 489818 452426 490054
rect 452662 489818 452746 490054
rect 452982 489818 488426 490054
rect 488662 489818 488746 490054
rect 488982 489818 524426 490054
rect 524662 489818 524746 490054
rect 524982 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 592650 490054
rect -8726 489734 592650 489818
rect -8726 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 344426 489734
rect 344662 489498 344746 489734
rect 344982 489498 380426 489734
rect 380662 489498 380746 489734
rect 380982 489498 416426 489734
rect 416662 489498 416746 489734
rect 416982 489498 452426 489734
rect 452662 489498 452746 489734
rect 452982 489498 488426 489734
rect 488662 489498 488746 489734
rect 488982 489498 524426 489734
rect 524662 489498 524746 489734
rect 524982 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 592650 489734
rect -8726 489466 592650 489498
rect -8726 486334 592650 486366
rect -8726 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 376706 486334
rect 376942 486098 377026 486334
rect 377262 486098 412706 486334
rect 412942 486098 413026 486334
rect 413262 486098 448706 486334
rect 448942 486098 449026 486334
rect 449262 486098 484706 486334
rect 484942 486098 485026 486334
rect 485262 486098 520706 486334
rect 520942 486098 521026 486334
rect 521262 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 592650 486334
rect -8726 486014 592650 486098
rect -8726 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 376706 486014
rect 376942 485778 377026 486014
rect 377262 485778 412706 486014
rect 412942 485778 413026 486014
rect 413262 485778 448706 486014
rect 448942 485778 449026 486014
rect 449262 485778 484706 486014
rect 484942 485778 485026 486014
rect 485262 485778 520706 486014
rect 520942 485778 521026 486014
rect 521262 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 592650 486014
rect -8726 485746 592650 485778
rect -8726 482614 592650 482646
rect -8726 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 592650 482294
rect -8726 482026 592650 482058
rect -8726 478894 592650 478926
rect -8726 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 592650 478894
rect -8726 478574 592650 478658
rect -8726 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 592650 478574
rect -8726 478306 592650 478338
rect -8726 475174 592650 475206
rect -8726 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 39610 475174
rect 39846 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 70330 475174
rect 70566 474938 101050 475174
rect 101286 474938 131770 475174
rect 132006 474938 162490 475174
rect 162726 474938 193210 475174
rect 193446 474938 223930 475174
rect 224166 474938 254650 475174
rect 254886 474938 285370 475174
rect 285606 474938 316090 475174
rect 316326 474938 346810 475174
rect 347046 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 592650 475174
rect -8726 474854 592650 474938
rect -8726 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 39610 474854
rect 39846 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 70330 474854
rect 70566 474618 101050 474854
rect 101286 474618 131770 474854
rect 132006 474618 162490 474854
rect 162726 474618 193210 474854
rect 193446 474618 223930 474854
rect 224166 474618 254650 474854
rect 254886 474618 285370 474854
rect 285606 474618 316090 474854
rect 316326 474618 346810 474854
rect 347046 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 592650 474854
rect -8726 474586 592650 474618
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 24250 471454
rect 24486 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 54970 471454
rect 55206 471218 85690 471454
rect 85926 471218 116410 471454
rect 116646 471218 147130 471454
rect 147366 471218 177850 471454
rect 178086 471218 208570 471454
rect 208806 471218 239290 471454
rect 239526 471218 270010 471454
rect 270246 471218 300730 471454
rect 300966 471218 331450 471454
rect 331686 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 24250 471134
rect 24486 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 54970 471134
rect 55206 470898 85690 471134
rect 85926 470898 116410 471134
rect 116646 470898 147130 471134
rect 147366 470898 177850 471134
rect 178086 470898 208570 471134
rect 208806 470898 239290 471134
rect 239526 470898 270010 471134
rect 270246 470898 300730 471134
rect 300966 470898 331450 471134
rect 331686 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 461494 592650 461526
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 351866 461494
rect 352102 461258 352186 461494
rect 352422 461258 387866 461494
rect 388102 461258 388186 461494
rect 388422 461258 423866 461494
rect 424102 461258 424186 461494
rect 424422 461258 459866 461494
rect 460102 461258 460186 461494
rect 460422 461258 495866 461494
rect 496102 461258 496186 461494
rect 496422 461258 531866 461494
rect 532102 461258 532186 461494
rect 532422 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect -8726 461174 592650 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 351866 461174
rect 352102 460938 352186 461174
rect 352422 460938 387866 461174
rect 388102 460938 388186 461174
rect 388422 460938 423866 461174
rect 424102 460938 424186 461174
rect 424422 460938 459866 461174
rect 460102 460938 460186 461174
rect 460422 460938 495866 461174
rect 496102 460938 496186 461174
rect 496422 460938 531866 461174
rect 532102 460938 532186 461174
rect 532422 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect -8726 460906 592650 460938
rect -8726 457774 592650 457806
rect -8726 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 348146 457774
rect 348382 457538 348466 457774
rect 348702 457538 384146 457774
rect 384382 457538 384466 457774
rect 384702 457538 420146 457774
rect 420382 457538 420466 457774
rect 420702 457538 456146 457774
rect 456382 457538 456466 457774
rect 456702 457538 492146 457774
rect 492382 457538 492466 457774
rect 492702 457538 528146 457774
rect 528382 457538 528466 457774
rect 528702 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 592650 457774
rect -8726 457454 592650 457538
rect -8726 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 348146 457454
rect 348382 457218 348466 457454
rect 348702 457218 384146 457454
rect 384382 457218 384466 457454
rect 384702 457218 420146 457454
rect 420382 457218 420466 457454
rect 420702 457218 456146 457454
rect 456382 457218 456466 457454
rect 456702 457218 492146 457454
rect 492382 457218 492466 457454
rect 492702 457218 528146 457454
rect 528382 457218 528466 457454
rect 528702 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 592650 457454
rect -8726 457186 592650 457218
rect -8726 454054 592650 454086
rect -8726 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 344426 454054
rect 344662 453818 344746 454054
rect 344982 453818 380426 454054
rect 380662 453818 380746 454054
rect 380982 453818 416426 454054
rect 416662 453818 416746 454054
rect 416982 453818 452426 454054
rect 452662 453818 452746 454054
rect 452982 454007 524426 454054
rect 452982 453818 488426 454007
rect -8726 453771 488426 453818
rect 488662 453771 488746 454007
rect 488982 453818 524426 454007
rect 524662 453818 524746 454054
rect 524982 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 592650 454054
rect 488982 453771 592650 453818
rect -8726 453734 592650 453771
rect -8726 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 344426 453734
rect 344662 453498 344746 453734
rect 344982 453498 380426 453734
rect 380662 453498 380746 453734
rect 380982 453498 416426 453734
rect 416662 453498 416746 453734
rect 416982 453498 452426 453734
rect 452662 453498 452746 453734
rect 452982 453498 524426 453734
rect 524662 453498 524746 453734
rect 524982 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 592650 453734
rect -8726 453466 592650 453498
rect -8726 450334 592650 450366
rect -8726 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 376706 450334
rect 376942 450098 377026 450334
rect 377262 450098 412706 450334
rect 412942 450098 413026 450334
rect 413262 450098 448706 450334
rect 448942 450098 449026 450334
rect 449262 450098 484706 450334
rect 484942 450098 485026 450334
rect 485262 450098 520706 450334
rect 520942 450098 521026 450334
rect 521262 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 592650 450334
rect -8726 450014 592650 450098
rect -8726 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 376706 450014
rect 376942 449778 377026 450014
rect 377262 449778 412706 450014
rect 412942 449778 413026 450014
rect 413262 449778 448706 450014
rect 448942 449778 449026 450014
rect 449262 449778 484706 450014
rect 484942 449778 485026 450014
rect 485262 449778 520706 450014
rect 520942 449778 521026 450014
rect 521262 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 592650 450014
rect -8726 449746 592650 449778
rect -8726 446614 592650 446646
rect -8726 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 592650 446294
rect -8726 446026 592650 446058
rect -8726 442894 592650 442926
rect -8726 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 592650 442894
rect -8726 442574 592650 442658
rect -8726 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 592650 442574
rect -8726 442306 592650 442338
rect -8726 439174 592650 439206
rect -8726 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 39610 439174
rect 39846 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 70330 439174
rect 70566 438938 101050 439174
rect 101286 438938 131770 439174
rect 132006 438938 162490 439174
rect 162726 438938 193210 439174
rect 193446 438938 223930 439174
rect 224166 438938 254650 439174
rect 254886 438938 285370 439174
rect 285606 438938 316090 439174
rect 316326 438938 346810 439174
rect 347046 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 426666 439174
rect 426902 438938 432347 439174
rect 432583 438938 438028 439174
rect 438264 438938 443709 439174
rect 443945 438938 475930 439174
rect 476166 438938 480875 439174
rect 481111 438938 485820 439174
rect 486056 438938 490765 439174
rect 491001 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 529426 439174
rect 529662 438938 537867 439174
rect 538103 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546308 439174
rect 546544 438938 554749 439174
rect 554985 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 592650 439174
rect -8726 438854 592650 438938
rect -8726 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 39610 438854
rect 39846 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 70330 438854
rect 70566 438618 101050 438854
rect 101286 438618 131770 438854
rect 132006 438618 162490 438854
rect 162726 438618 193210 438854
rect 193446 438618 223930 438854
rect 224166 438618 254650 438854
rect 254886 438618 285370 438854
rect 285606 438618 316090 438854
rect 316326 438618 346810 438854
rect 347046 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 426666 438854
rect 426902 438618 432347 438854
rect 432583 438618 438028 438854
rect 438264 438618 443709 438854
rect 443945 438618 475930 438854
rect 476166 438618 480875 438854
rect 481111 438618 485820 438854
rect 486056 438618 490765 438854
rect 491001 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 529426 438854
rect 529662 438618 537867 438854
rect 538103 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546308 438854
rect 546544 438618 554749 438854
rect 554985 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 592650 438854
rect -8726 438586 592650 438618
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 24250 435454
rect 24486 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 54970 435454
rect 55206 435218 85690 435454
rect 85926 435218 116410 435454
rect 116646 435218 147130 435454
rect 147366 435218 177850 435454
rect 178086 435218 208570 435454
rect 208806 435218 239290 435454
rect 239526 435218 270010 435454
rect 270246 435218 300730 435454
rect 300966 435218 331450 435454
rect 331686 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 423826 435454
rect 424062 435218 429507 435454
rect 429743 435218 435188 435454
rect 435424 435218 440869 435454
rect 441105 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 473458 435454
rect 473694 435218 478403 435454
rect 478639 435218 483348 435454
rect 483584 435218 488293 435454
rect 488529 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 525206 435454
rect 525442 435218 533647 435454
rect 533883 435218 542088 435454
rect 542324 435218 550529 435454
rect 550765 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 24250 435134
rect 24486 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 54970 435134
rect 55206 434898 85690 435134
rect 85926 434898 116410 435134
rect 116646 434898 147130 435134
rect 147366 434898 177850 435134
rect 178086 434898 208570 435134
rect 208806 434898 239290 435134
rect 239526 434898 270010 435134
rect 270246 434898 300730 435134
rect 300966 434898 331450 435134
rect 331686 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 423826 435134
rect 424062 434898 429507 435134
rect 429743 434898 435188 435134
rect 435424 434898 440869 435134
rect 441105 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 473458 435134
rect 473694 434898 478403 435134
rect 478639 434898 483348 435134
rect 483584 434898 488293 435134
rect 488529 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 525206 435134
rect 525442 434898 533647 435134
rect 533883 434898 542088 435134
rect 542324 434898 550529 435134
rect 550765 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 425494 592650 425526
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 351866 425494
rect 352102 425258 352186 425494
rect 352422 425258 387866 425494
rect 388102 425258 388186 425494
rect 388422 425258 459866 425494
rect 460102 425258 460186 425494
rect 460422 425258 495866 425494
rect 496102 425258 496186 425494
rect 496422 425258 531866 425494
rect 532102 425258 532186 425494
rect 532422 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect -8726 425174 592650 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 351866 425174
rect 352102 424938 352186 425174
rect 352422 424938 387866 425174
rect 388102 424938 388186 425174
rect 388422 424938 459866 425174
rect 460102 424938 460186 425174
rect 460422 424938 495866 425174
rect 496102 424938 496186 425174
rect 496422 424938 531866 425174
rect 532102 424938 532186 425174
rect 532422 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect -8726 424906 592650 424938
rect -8726 421774 592650 421806
rect -8726 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 348146 421774
rect 348382 421538 348466 421774
rect 348702 421538 384146 421774
rect 384382 421538 384466 421774
rect 384702 421538 420146 421774
rect 420382 421538 420466 421774
rect 420702 421538 456146 421774
rect 456382 421538 456466 421774
rect 456702 421538 492146 421774
rect 492382 421538 492466 421774
rect 492702 421538 528146 421774
rect 528382 421538 528466 421774
rect 528702 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 592650 421774
rect -8726 421454 592650 421538
rect -8726 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 348146 421454
rect 348382 421218 348466 421454
rect 348702 421218 384146 421454
rect 384382 421218 384466 421454
rect 384702 421218 420146 421454
rect 420382 421218 420466 421454
rect 420702 421218 456146 421454
rect 456382 421218 456466 421454
rect 456702 421218 492146 421454
rect 492382 421218 492466 421454
rect 492702 421218 528146 421454
rect 528382 421218 528466 421454
rect 528702 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 592650 421454
rect -8726 421186 592650 421218
rect -8726 418054 592650 418086
rect -8726 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 344426 418054
rect 344662 417818 344746 418054
rect 344982 417818 380426 418054
rect 380662 417818 380746 418054
rect 380982 417818 416426 418054
rect 416662 417818 416746 418054
rect 416982 417818 452426 418054
rect 452662 417818 452746 418054
rect 452982 417818 524426 418054
rect 524662 417818 524746 418054
rect 524982 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 592650 418054
rect -8726 417734 592650 417818
rect -8726 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 344426 417734
rect 344662 417498 344746 417734
rect 344982 417498 380426 417734
rect 380662 417498 380746 417734
rect 380982 417498 416426 417734
rect 416662 417498 416746 417734
rect 416982 417498 452426 417734
rect 452662 417498 452746 417734
rect 452982 417498 524426 417734
rect 524662 417498 524746 417734
rect 524982 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 592650 417734
rect -8726 417466 592650 417498
rect -8726 414334 592650 414366
rect -8726 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 376706 414334
rect 376942 414098 377026 414334
rect 377262 414098 412706 414334
rect 412942 414098 413026 414334
rect 413262 414098 448706 414334
rect 448942 414098 449026 414334
rect 449262 414098 484706 414334
rect 484942 414098 485026 414334
rect 485262 414098 520706 414334
rect 520942 414098 521026 414334
rect 521262 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 592650 414334
rect -8726 414014 592650 414098
rect -8726 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 376706 414014
rect 376942 413778 377026 414014
rect 377262 413778 412706 414014
rect 412942 413778 413026 414014
rect 413262 413778 448706 414014
rect 448942 413778 449026 414014
rect 449262 413778 484706 414014
rect 484942 413778 485026 414014
rect 485262 413778 520706 414014
rect 520942 413778 521026 414014
rect 521262 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 592650 414014
rect -8726 413746 592650 413778
rect -8726 410614 592650 410646
rect -8726 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 592650 410294
rect -8726 410026 592650 410058
rect -8726 406894 592650 406926
rect -8726 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 592650 406894
rect -8726 406574 592650 406658
rect -8726 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 592650 406574
rect -8726 406306 592650 406338
rect -8726 403174 592650 403206
rect -8726 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 39610 403174
rect 39846 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 70330 403174
rect 70566 402938 101050 403174
rect 101286 402938 131770 403174
rect 132006 402938 162490 403174
rect 162726 402938 193210 403174
rect 193446 402938 223930 403174
rect 224166 402938 254650 403174
rect 254886 402938 285370 403174
rect 285606 402938 316090 403174
rect 316326 402938 346810 403174
rect 347046 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 592650 403174
rect -8726 402854 592650 402938
rect -8726 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 39610 402854
rect 39846 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 70330 402854
rect 70566 402618 101050 402854
rect 101286 402618 131770 402854
rect 132006 402618 162490 402854
rect 162726 402618 193210 402854
rect 193446 402618 223930 402854
rect 224166 402618 254650 402854
rect 254886 402618 285370 402854
rect 285606 402618 316090 402854
rect 316326 402618 346810 402854
rect 347046 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 592650 402854
rect -8726 402586 592650 402618
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 24250 399454
rect 24486 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 54970 399454
rect 55206 399218 85690 399454
rect 85926 399218 116410 399454
rect 116646 399218 147130 399454
rect 147366 399218 177850 399454
rect 178086 399218 208570 399454
rect 208806 399218 239290 399454
rect 239526 399218 270010 399454
rect 270246 399218 300730 399454
rect 300966 399218 331450 399454
rect 331686 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 24250 399134
rect 24486 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 54970 399134
rect 55206 398898 85690 399134
rect 85926 398898 116410 399134
rect 116646 398898 147130 399134
rect 147366 398898 177850 399134
rect 178086 398898 208570 399134
rect 208806 398898 239290 399134
rect 239526 398898 270010 399134
rect 270246 398898 300730 399134
rect 300966 398898 331450 399134
rect 331686 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 389494 592650 389526
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 351866 389494
rect 352102 389258 352186 389494
rect 352422 389258 387866 389494
rect 388102 389258 388186 389494
rect 388422 389258 423866 389494
rect 424102 389258 424186 389494
rect 424422 389258 459866 389494
rect 460102 389258 460186 389494
rect 460422 389258 495866 389494
rect 496102 389258 496186 389494
rect 496422 389258 531866 389494
rect 532102 389258 532186 389494
rect 532422 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect -8726 389174 592650 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 351866 389174
rect 352102 388938 352186 389174
rect 352422 388938 387866 389174
rect 388102 388938 388186 389174
rect 388422 388938 423866 389174
rect 424102 388938 424186 389174
rect 424422 388938 459866 389174
rect 460102 388938 460186 389174
rect 460422 388938 495866 389174
rect 496102 388938 496186 389174
rect 496422 388938 531866 389174
rect 532102 388938 532186 389174
rect 532422 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect -8726 388906 592650 388938
rect -8726 385774 592650 385806
rect -8726 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 348146 385774
rect 348382 385538 348466 385774
rect 348702 385538 384146 385774
rect 384382 385538 384466 385774
rect 384702 385538 420146 385774
rect 420382 385538 420466 385774
rect 420702 385538 456146 385774
rect 456382 385538 456466 385774
rect 456702 385538 528146 385774
rect 528382 385538 528466 385774
rect 528702 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 592650 385774
rect -8726 385454 592650 385538
rect -8726 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 348146 385454
rect 348382 385218 348466 385454
rect 348702 385218 384146 385454
rect 384382 385218 384466 385454
rect 384702 385218 420146 385454
rect 420382 385218 420466 385454
rect 420702 385218 456146 385454
rect 456382 385218 456466 385454
rect 456702 385218 528146 385454
rect 528382 385218 528466 385454
rect 528702 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 592650 385454
rect -8726 385186 592650 385218
rect -8726 382054 592650 382086
rect -8726 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 344426 382054
rect 344662 381818 344746 382054
rect 344982 381818 380426 382054
rect 380662 381818 380746 382054
rect 380982 381818 416426 382054
rect 416662 381818 416746 382054
rect 416982 381818 452426 382054
rect 452662 381818 452746 382054
rect 452982 381818 524426 382054
rect 524662 381818 524746 382054
rect 524982 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 592650 382054
rect -8726 381734 592650 381818
rect -8726 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 344426 381734
rect 344662 381498 344746 381734
rect 344982 381498 380426 381734
rect 380662 381498 380746 381734
rect 380982 381498 416426 381734
rect 416662 381498 416746 381734
rect 416982 381498 452426 381734
rect 452662 381498 452746 381734
rect 452982 381498 524426 381734
rect 524662 381498 524746 381734
rect 524982 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 592650 381734
rect -8726 381466 592650 381498
rect -8726 378334 592650 378366
rect -8726 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 376706 378334
rect 376942 378098 377026 378334
rect 377262 378098 412706 378334
rect 412942 378098 413026 378334
rect 413262 378098 448706 378334
rect 448942 378098 449026 378334
rect 449262 378098 520706 378334
rect 520942 378098 521026 378334
rect 521262 378243 589182 378334
rect 521262 378098 556706 378243
rect -8726 378014 556706 378098
rect -8726 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 376706 378014
rect 376942 377778 377026 378014
rect 377262 377778 412706 378014
rect 412942 377778 413026 378014
rect 413262 377778 448706 378014
rect 448942 377778 449026 378014
rect 449262 377778 520706 378014
rect 520942 377778 521026 378014
rect 521262 378007 556706 378014
rect 556942 378007 557026 378243
rect 557262 378098 589182 378243
rect 589418 378098 589502 378334
rect 589738 378098 592650 378334
rect 557262 378014 592650 378098
rect 557262 378007 589182 378014
rect 521262 377778 589182 378007
rect 589418 377778 589502 378014
rect 589738 377778 592650 378014
rect -8726 377746 592650 377778
rect -8726 374614 592650 374646
rect -8726 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 592650 374294
rect -8726 374026 592650 374058
rect -8726 370894 592650 370926
rect -8726 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 592650 370894
rect -8726 370574 592650 370658
rect -8726 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 592650 370574
rect -8726 370306 592650 370338
rect -8726 367174 592650 367206
rect -8726 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 39610 367174
rect 39846 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 70330 367174
rect 70566 366938 101050 367174
rect 101286 366938 131770 367174
rect 132006 366938 162490 367174
rect 162726 366938 193210 367174
rect 193446 366938 223930 367174
rect 224166 366938 254650 367174
rect 254886 366938 285370 367174
rect 285606 366938 316090 367174
rect 316326 366938 346810 367174
rect 347046 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 469610 367174
rect 469846 366938 500330 367174
rect 500566 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 554918 367174
rect 555154 366938 558851 367174
rect 559087 366938 562784 367174
rect 563020 366938 566717 367174
rect 566953 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 592650 367174
rect -8726 366854 592650 366938
rect -8726 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 39610 366854
rect 39846 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 70330 366854
rect 70566 366618 101050 366854
rect 101286 366618 131770 366854
rect 132006 366618 162490 366854
rect 162726 366618 193210 366854
rect 193446 366618 223930 366854
rect 224166 366618 254650 366854
rect 254886 366618 285370 366854
rect 285606 366618 316090 366854
rect 316326 366618 346810 366854
rect 347046 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 469610 366854
rect 469846 366618 500330 366854
rect 500566 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 554918 366854
rect 555154 366618 558851 366854
rect 559087 366618 562784 366854
rect 563020 366618 566717 366854
rect 566953 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 592650 366854
rect -8726 366586 592650 366618
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 24250 363454
rect 24486 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 54970 363454
rect 55206 363218 85690 363454
rect 85926 363218 116410 363454
rect 116646 363218 147130 363454
rect 147366 363218 177850 363454
rect 178086 363218 208570 363454
rect 208806 363218 239290 363454
rect 239526 363218 270010 363454
rect 270246 363218 300730 363454
rect 300966 363218 331450 363454
rect 331686 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 454250 363454
rect 454486 363218 484970 363454
rect 485206 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 552952 363454
rect 553188 363218 556885 363454
rect 557121 363218 560818 363454
rect 561054 363218 564751 363454
rect 564987 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 24250 363134
rect 24486 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 54970 363134
rect 55206 362898 85690 363134
rect 85926 362898 116410 363134
rect 116646 362898 147130 363134
rect 147366 362898 177850 363134
rect 178086 362898 208570 363134
rect 208806 362898 239290 363134
rect 239526 362898 270010 363134
rect 270246 362898 300730 363134
rect 300966 362898 331450 363134
rect 331686 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 454250 363134
rect 454486 362898 484970 363134
rect 485206 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 552952 363134
rect 553188 362898 556885 363134
rect 557121 362898 560818 363134
rect 561054 362898 564751 363134
rect 564987 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 353494 592650 353526
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 351866 353494
rect 352102 353258 352186 353494
rect 352422 353258 387866 353494
rect 388102 353258 388186 353494
rect 388422 353258 423866 353494
rect 424102 353258 424186 353494
rect 424422 353258 459866 353494
rect 460102 353258 460186 353494
rect 460422 353258 531866 353494
rect 532102 353258 532186 353494
rect 532422 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect -8726 353174 592650 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 351866 353174
rect 352102 352938 352186 353174
rect 352422 352938 387866 353174
rect 388102 352938 388186 353174
rect 388422 352938 423866 353174
rect 424102 352938 424186 353174
rect 424422 352938 459866 353174
rect 460102 352938 460186 353174
rect 460422 352938 531866 353174
rect 532102 352938 532186 353174
rect 532422 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect -8726 352906 592650 352938
rect -8726 349774 592650 349806
rect -8726 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 348146 349774
rect 348382 349538 348466 349774
rect 348702 349538 384146 349774
rect 384382 349538 384466 349774
rect 384702 349538 420146 349774
rect 420382 349538 420466 349774
rect 420702 349538 456146 349774
rect 456382 349538 456466 349774
rect 456702 349538 528146 349774
rect 528382 349538 528466 349774
rect 528702 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 592650 349774
rect -8726 349454 592650 349538
rect -8726 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 348146 349454
rect 348382 349218 348466 349454
rect 348702 349218 384146 349454
rect 384382 349218 384466 349454
rect 384702 349218 420146 349454
rect 420382 349218 420466 349454
rect 420702 349218 456146 349454
rect 456382 349218 456466 349454
rect 456702 349218 528146 349454
rect 528382 349218 528466 349454
rect 528702 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 592650 349454
rect -8726 349186 592650 349218
rect -8726 346054 592650 346086
rect -8726 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 344426 346054
rect 344662 345818 344746 346054
rect 344982 345818 380426 346054
rect 380662 345818 380746 346054
rect 380982 345818 416426 346054
rect 416662 345818 416746 346054
rect 416982 345818 452426 346054
rect 452662 345818 452746 346054
rect 452982 345818 524426 346054
rect 524662 345818 524746 346054
rect 524982 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 592650 346054
rect -8726 345734 592650 345818
rect -8726 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 344426 345734
rect 344662 345498 344746 345734
rect 344982 345498 380426 345734
rect 380662 345498 380746 345734
rect 380982 345498 416426 345734
rect 416662 345498 416746 345734
rect 416982 345498 452426 345734
rect 452662 345498 452746 345734
rect 452982 345498 524426 345734
rect 524662 345498 524746 345734
rect 524982 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 592650 345734
rect -8726 345466 592650 345498
rect -8726 342334 592650 342366
rect -8726 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 376706 342334
rect 376942 342098 377026 342334
rect 377262 342098 412706 342334
rect 412942 342098 413026 342334
rect 413262 342098 448706 342334
rect 448942 342098 449026 342334
rect 449262 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 592650 342334
rect -8726 342014 592650 342098
rect -8726 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 376706 342014
rect 376942 341778 377026 342014
rect 377262 341778 412706 342014
rect 412942 341778 413026 342014
rect 413262 341778 448706 342014
rect 448942 341778 449026 342014
rect 449262 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 592650 342014
rect -8726 341746 592650 341778
rect -8726 338614 592650 338646
rect -8726 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 592650 338294
rect -8726 338026 592650 338058
rect -8726 334894 592650 334926
rect -8726 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 592650 334894
rect -8726 334574 592650 334658
rect -8726 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 592650 334574
rect -8726 334306 592650 334338
rect -8726 331174 592650 331206
rect -8726 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 39610 331174
rect 39846 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 70330 331174
rect 70566 330938 101050 331174
rect 101286 330938 131770 331174
rect 132006 330938 162490 331174
rect 162726 330938 193210 331174
rect 193446 330938 223930 331174
rect 224166 330938 254650 331174
rect 254886 330938 285370 331174
rect 285606 330938 316090 331174
rect 316326 330938 346810 331174
rect 347046 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 407932 331174
rect 408168 330938 414878 331174
rect 415114 330938 421824 331174
rect 422060 330938 428770 331174
rect 429006 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 469610 331174
rect 469846 330938 500330 331174
rect 500566 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 592650 331174
rect -8726 330854 592650 330938
rect -8726 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 39610 330854
rect 39846 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 70330 330854
rect 70566 330618 101050 330854
rect 101286 330618 131770 330854
rect 132006 330618 162490 330854
rect 162726 330618 193210 330854
rect 193446 330618 223930 330854
rect 224166 330618 254650 330854
rect 254886 330618 285370 330854
rect 285606 330618 316090 330854
rect 316326 330618 346810 330854
rect 347046 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 407932 330854
rect 408168 330618 414878 330854
rect 415114 330618 421824 330854
rect 422060 330618 428770 330854
rect 429006 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 469610 330854
rect 469846 330618 500330 330854
rect 500566 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 592650 330854
rect -8726 330586 592650 330618
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 24250 327454
rect 24486 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 54970 327454
rect 55206 327218 85690 327454
rect 85926 327218 116410 327454
rect 116646 327218 147130 327454
rect 147366 327218 177850 327454
rect 178086 327218 208570 327454
rect 208806 327218 239290 327454
rect 239526 327218 270010 327454
rect 270246 327218 300730 327454
rect 300966 327218 331450 327454
rect 331686 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 404459 327454
rect 404695 327218 411405 327454
rect 411641 327218 418351 327454
rect 418587 327218 425297 327454
rect 425533 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 454250 327454
rect 454486 327218 484970 327454
rect 485206 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 24250 327134
rect 24486 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 54970 327134
rect 55206 326898 85690 327134
rect 85926 326898 116410 327134
rect 116646 326898 147130 327134
rect 147366 326898 177850 327134
rect 178086 326898 208570 327134
rect 208806 326898 239290 327134
rect 239526 326898 270010 327134
rect 270246 326898 300730 327134
rect 300966 326898 331450 327134
rect 331686 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 404459 327134
rect 404695 326898 411405 327134
rect 411641 326898 418351 327134
rect 418587 326898 425297 327134
rect 425533 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 454250 327134
rect 454486 326898 484970 327134
rect 485206 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 317494 592650 317526
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 351866 317494
rect 352102 317258 352186 317494
rect 352422 317258 387866 317494
rect 388102 317258 388186 317494
rect 388422 317258 423866 317494
rect 424102 317258 424186 317494
rect 424422 317258 459866 317494
rect 460102 317258 460186 317494
rect 460422 317258 495866 317494
rect 496102 317258 496186 317494
rect 496422 317258 531866 317494
rect 532102 317258 532186 317494
rect 532422 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect -8726 317174 592650 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 351866 317174
rect 352102 316938 352186 317174
rect 352422 316938 387866 317174
rect 388102 316938 388186 317174
rect 388422 316938 423866 317174
rect 424102 316938 424186 317174
rect 424422 316938 459866 317174
rect 460102 316938 460186 317174
rect 460422 316938 495866 317174
rect 496102 316938 496186 317174
rect 496422 316938 531866 317174
rect 532102 316938 532186 317174
rect 532422 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect -8726 316906 592650 316938
rect -8726 313774 592650 313806
rect -8726 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 348146 313774
rect 348382 313538 348466 313774
rect 348702 313538 384146 313774
rect 384382 313538 384466 313774
rect 384702 313538 420146 313774
rect 420382 313538 420466 313774
rect 420702 313538 456146 313774
rect 456382 313538 456466 313774
rect 456702 313538 492146 313774
rect 492382 313538 492466 313774
rect 492702 313538 528146 313774
rect 528382 313538 528466 313774
rect 528702 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 592650 313774
rect -8726 313454 592650 313538
rect -8726 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 348146 313454
rect 348382 313218 348466 313454
rect 348702 313218 384146 313454
rect 384382 313218 384466 313454
rect 384702 313218 420146 313454
rect 420382 313218 420466 313454
rect 420702 313218 456146 313454
rect 456382 313218 456466 313454
rect 456702 313218 492146 313454
rect 492382 313218 492466 313454
rect 492702 313218 528146 313454
rect 528382 313218 528466 313454
rect 528702 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 592650 313454
rect -8726 313186 592650 313218
rect -8726 310054 592650 310086
rect -8726 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 344426 310054
rect 344662 309818 344746 310054
rect 344982 309818 380426 310054
rect 380662 309818 380746 310054
rect 380982 309818 416426 310054
rect 416662 309818 416746 310054
rect 416982 309818 452426 310054
rect 452662 309818 452746 310054
rect 452982 309818 488426 310054
rect 488662 309818 488746 310054
rect 488982 309818 524426 310054
rect 524662 309818 524746 310054
rect 524982 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 592650 310054
rect -8726 309734 592650 309818
rect -8726 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 344426 309734
rect 344662 309498 344746 309734
rect 344982 309498 380426 309734
rect 380662 309498 380746 309734
rect 380982 309498 416426 309734
rect 416662 309498 416746 309734
rect 416982 309498 452426 309734
rect 452662 309498 452746 309734
rect 452982 309498 488426 309734
rect 488662 309498 488746 309734
rect 488982 309498 524426 309734
rect 524662 309498 524746 309734
rect 524982 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 592650 309734
rect -8726 309466 592650 309498
rect -8726 306334 592650 306366
rect -8726 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 376706 306334
rect 376942 306098 377026 306334
rect 377262 306098 412706 306334
rect 412942 306098 413026 306334
rect 413262 306098 448706 306334
rect 448942 306098 449026 306334
rect 449262 306098 484706 306334
rect 484942 306098 485026 306334
rect 485262 306098 520706 306334
rect 520942 306098 521026 306334
rect 521262 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 592650 306334
rect -8726 306014 592650 306098
rect -8726 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 376706 306014
rect 376942 305778 377026 306014
rect 377262 305778 412706 306014
rect 412942 305778 413026 306014
rect 413262 305778 448706 306014
rect 448942 305778 449026 306014
rect 449262 305778 484706 306014
rect 484942 305778 485026 306014
rect 485262 305778 520706 306014
rect 520942 305778 521026 306014
rect 521262 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 592650 306014
rect -8726 305746 592650 305778
rect -8726 302614 592650 302646
rect -8726 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 592650 302294
rect -8726 302026 592650 302058
rect -8726 298894 592650 298926
rect -8726 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 592650 298894
rect -8726 298574 592650 298658
rect -8726 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 592650 298574
rect -8726 298306 592650 298338
rect -8726 295174 592650 295206
rect -8726 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 39610 295174
rect 39846 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 70330 295174
rect 70566 294938 101050 295174
rect 101286 294938 131770 295174
rect 132006 294938 162490 295174
rect 162726 294938 193210 295174
rect 193446 294938 223930 295174
rect 224166 294938 254650 295174
rect 254886 294938 285370 295174
rect 285606 294938 316090 295174
rect 316326 294938 346810 295174
rect 347046 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 592650 295174
rect -8726 294854 592650 294938
rect -8726 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 39610 294854
rect 39846 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 70330 294854
rect 70566 294618 101050 294854
rect 101286 294618 131770 294854
rect 132006 294618 162490 294854
rect 162726 294618 193210 294854
rect 193446 294618 223930 294854
rect 224166 294618 254650 294854
rect 254886 294618 285370 294854
rect 285606 294618 316090 294854
rect 316326 294618 346810 294854
rect 347046 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 592650 294854
rect -8726 294586 592650 294618
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 24250 291454
rect 24486 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 54970 291454
rect 55206 291218 85690 291454
rect 85926 291218 116410 291454
rect 116646 291218 147130 291454
rect 147366 291218 177850 291454
rect 178086 291218 208570 291454
rect 208806 291218 239290 291454
rect 239526 291218 270010 291454
rect 270246 291218 300730 291454
rect 300966 291218 331450 291454
rect 331686 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 24250 291134
rect 24486 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 54970 291134
rect 55206 290898 85690 291134
rect 85926 290898 116410 291134
rect 116646 290898 147130 291134
rect 147366 290898 177850 291134
rect 178086 290898 208570 291134
rect 208806 290898 239290 291134
rect 239526 290898 270010 291134
rect 270246 290898 300730 291134
rect 300966 290898 331450 291134
rect 331686 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 281494 592650 281526
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 351866 281494
rect 352102 281258 352186 281494
rect 352422 281258 387866 281494
rect 388102 281258 388186 281494
rect 388422 281258 423866 281494
rect 424102 281258 424186 281494
rect 424422 281258 459866 281494
rect 460102 281258 460186 281494
rect 460422 281258 495866 281494
rect 496102 281258 496186 281494
rect 496422 281258 531866 281494
rect 532102 281258 532186 281494
rect 532422 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect -8726 281174 592650 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 351866 281174
rect 352102 280938 352186 281174
rect 352422 280938 387866 281174
rect 388102 280938 388186 281174
rect 388422 280938 423866 281174
rect 424102 280938 424186 281174
rect 424422 280938 459866 281174
rect 460102 280938 460186 281174
rect 460422 280938 495866 281174
rect 496102 280938 496186 281174
rect 496422 280938 531866 281174
rect 532102 280938 532186 281174
rect 532422 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect -8726 280906 592650 280938
rect -8726 277774 592650 277806
rect -8726 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 348146 277774
rect 348382 277538 348466 277774
rect 348702 277538 384146 277774
rect 384382 277538 384466 277774
rect 384702 277538 420146 277774
rect 420382 277538 420466 277774
rect 420702 277538 456146 277774
rect 456382 277538 456466 277774
rect 456702 277538 492146 277774
rect 492382 277538 492466 277774
rect 492702 277538 528146 277774
rect 528382 277538 528466 277774
rect 528702 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 592650 277774
rect -8726 277454 592650 277538
rect -8726 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 348146 277454
rect 348382 277218 348466 277454
rect 348702 277218 384146 277454
rect 384382 277218 384466 277454
rect 384702 277218 420146 277454
rect 420382 277218 420466 277454
rect 420702 277218 456146 277454
rect 456382 277218 456466 277454
rect 456702 277218 492146 277454
rect 492382 277218 492466 277454
rect 492702 277218 528146 277454
rect 528382 277218 528466 277454
rect 528702 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 592650 277454
rect -8726 277186 592650 277218
rect -8726 274054 592650 274086
rect -8726 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 344426 274054
rect 344662 273818 344746 274054
rect 344982 273818 380426 274054
rect 380662 273818 380746 274054
rect 380982 273818 416426 274054
rect 416662 273818 416746 274054
rect 416982 273818 452426 274054
rect 452662 273818 452746 274054
rect 452982 273818 488426 274054
rect 488662 273818 488746 274054
rect 488982 273818 524426 274054
rect 524662 273818 524746 274054
rect 524982 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 592650 274054
rect -8726 273734 592650 273818
rect -8726 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 344426 273734
rect 344662 273498 344746 273734
rect 344982 273498 380426 273734
rect 380662 273498 380746 273734
rect 380982 273498 416426 273734
rect 416662 273498 416746 273734
rect 416982 273498 452426 273734
rect 452662 273498 452746 273734
rect 452982 273498 488426 273734
rect 488662 273498 488746 273734
rect 488982 273498 524426 273734
rect 524662 273498 524746 273734
rect 524982 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 592650 273734
rect -8726 273466 592650 273498
rect -8726 270334 592650 270366
rect -8726 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 376706 270334
rect 376942 270098 377026 270334
rect 377262 270098 412706 270334
rect 412942 270098 413026 270334
rect 413262 270098 448706 270334
rect 448942 270098 449026 270334
rect 449262 270098 484706 270334
rect 484942 270098 485026 270334
rect 485262 270098 520706 270334
rect 520942 270098 521026 270334
rect 521262 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 592650 270334
rect -8726 270014 592650 270098
rect -8726 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 376706 270014
rect 376942 269778 377026 270014
rect 377262 269778 412706 270014
rect 412942 269778 413026 270014
rect 413262 269778 448706 270014
rect 448942 269778 449026 270014
rect 449262 269778 484706 270014
rect 484942 269778 485026 270014
rect 485262 269778 520706 270014
rect 520942 269778 521026 270014
rect 521262 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 592650 270014
rect -8726 269746 592650 269778
rect -8726 266614 592650 266646
rect -8726 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 592650 266294
rect -8726 266026 592650 266058
rect -8726 262894 592650 262926
rect -8726 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 592650 262894
rect -8726 262574 592650 262658
rect -8726 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 592650 262574
rect -8726 262306 592650 262338
rect -8726 259174 592650 259206
rect -8726 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 39610 259174
rect 39846 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 70330 259174
rect 70566 258938 101050 259174
rect 101286 258938 131770 259174
rect 132006 258938 162490 259174
rect 162726 258938 193210 259174
rect 193446 258938 223930 259174
rect 224166 258938 254650 259174
rect 254886 258938 285370 259174
rect 285606 258938 316090 259174
rect 316326 258938 346810 259174
rect 347046 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 479610 259174
rect 479846 258938 510330 259174
rect 510566 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 592650 259174
rect -8726 258854 592650 258938
rect -8726 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 39610 258854
rect 39846 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 70330 258854
rect 70566 258618 101050 258854
rect 101286 258618 131770 258854
rect 132006 258618 162490 258854
rect 162726 258618 193210 258854
rect 193446 258618 223930 258854
rect 224166 258618 254650 258854
rect 254886 258618 285370 258854
rect 285606 258618 316090 258854
rect 316326 258618 346810 258854
rect 347046 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 479610 258854
rect 479846 258618 510330 258854
rect 510566 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 592650 258854
rect -8726 258586 592650 258618
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 24250 255454
rect 24486 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 54970 255454
rect 55206 255218 85690 255454
rect 85926 255218 116410 255454
rect 116646 255218 147130 255454
rect 147366 255218 177850 255454
rect 178086 255218 208570 255454
rect 208806 255218 239290 255454
rect 239526 255218 270010 255454
rect 270246 255218 300730 255454
rect 300966 255218 331450 255454
rect 331686 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 464250 255454
rect 464486 255218 494970 255454
rect 495206 255218 525690 255454
rect 525926 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 24250 255134
rect 24486 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 54970 255134
rect 55206 254898 85690 255134
rect 85926 254898 116410 255134
rect 116646 254898 147130 255134
rect 147366 254898 177850 255134
rect 178086 254898 208570 255134
rect 208806 254898 239290 255134
rect 239526 254898 270010 255134
rect 270246 254898 300730 255134
rect 300966 254898 331450 255134
rect 331686 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 464250 255134
rect 464486 254898 494970 255134
rect 495206 254898 525690 255134
rect 525926 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 245494 592650 245526
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 351866 245494
rect 352102 245258 352186 245494
rect 352422 245258 387866 245494
rect 388102 245258 388186 245494
rect 388422 245258 423866 245494
rect 424102 245258 424186 245494
rect 424422 245258 459866 245494
rect 460102 245258 460186 245494
rect 460422 245258 531866 245494
rect 532102 245258 532186 245494
rect 532422 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect -8726 245174 592650 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 351866 245174
rect 352102 244938 352186 245174
rect 352422 244938 387866 245174
rect 388102 244938 388186 245174
rect 388422 244938 423866 245174
rect 424102 244938 424186 245174
rect 424422 244938 459866 245174
rect 460102 244938 460186 245174
rect 460422 244938 531866 245174
rect 532102 244938 532186 245174
rect 532422 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect -8726 244906 592650 244938
rect -8726 241774 592650 241806
rect -8726 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 348146 241774
rect 348382 241538 348466 241774
rect 348702 241538 384146 241774
rect 384382 241538 384466 241774
rect 384702 241538 420146 241774
rect 420382 241538 420466 241774
rect 420702 241538 456146 241774
rect 456382 241538 456466 241774
rect 456702 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 592650 241774
rect -8726 241454 592650 241538
rect -8726 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 348146 241454
rect 348382 241218 348466 241454
rect 348702 241218 384146 241454
rect 384382 241218 384466 241454
rect 384702 241218 420146 241454
rect 420382 241218 420466 241454
rect 420702 241218 456146 241454
rect 456382 241218 456466 241454
rect 456702 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 592650 241454
rect -8726 241186 592650 241218
rect -8726 238054 592650 238086
rect -8726 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 344426 238054
rect 344662 237818 344746 238054
rect 344982 237818 380426 238054
rect 380662 237818 380746 238054
rect 380982 237818 416426 238054
rect 416662 237818 416746 238054
rect 416982 237818 452426 238054
rect 452662 237818 452746 238054
rect 452982 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 592650 238054
rect -8726 237734 592650 237818
rect -8726 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 344426 237734
rect 344662 237498 344746 237734
rect 344982 237498 380426 237734
rect 380662 237498 380746 237734
rect 380982 237498 416426 237734
rect 416662 237498 416746 237734
rect 416982 237498 452426 237734
rect 452662 237498 452746 237734
rect 452982 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 592650 237734
rect -8726 237466 592650 237498
rect -8726 234334 592650 234366
rect -8726 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 376706 234334
rect 376942 234098 377026 234334
rect 377262 234098 412706 234334
rect 412942 234098 413026 234334
rect 413262 234098 448706 234334
rect 448942 234098 449026 234334
rect 449262 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 592650 234334
rect -8726 234014 592650 234098
rect -8726 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 376706 234014
rect 376942 233778 377026 234014
rect 377262 233778 412706 234014
rect 412942 233778 413026 234014
rect 413262 233778 448706 234014
rect 448942 233778 449026 234014
rect 449262 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 592650 234014
rect -8726 233746 592650 233778
rect -8726 230614 592650 230646
rect -8726 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 592650 230294
rect -8726 230026 592650 230058
rect -8726 226894 592650 226926
rect -8726 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 592650 226894
rect -8726 226574 592650 226658
rect -8726 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 592650 226574
rect -8726 226306 592650 226338
rect -8726 223174 592650 223206
rect -8726 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 39610 223174
rect 39846 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 70330 223174
rect 70566 222938 101050 223174
rect 101286 222938 131770 223174
rect 132006 222938 162490 223174
rect 162726 222938 193210 223174
rect 193446 222938 223930 223174
rect 224166 222938 254650 223174
rect 254886 222938 285370 223174
rect 285606 222938 316090 223174
rect 316326 222938 346810 223174
rect 347046 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 479610 223174
rect 479846 222938 510330 223174
rect 510566 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 592650 223174
rect -8726 222854 592650 222938
rect -8726 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 39610 222854
rect 39846 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 70330 222854
rect 70566 222618 101050 222854
rect 101286 222618 131770 222854
rect 132006 222618 162490 222854
rect 162726 222618 193210 222854
rect 193446 222618 223930 222854
rect 224166 222618 254650 222854
rect 254886 222618 285370 222854
rect 285606 222618 316090 222854
rect 316326 222618 346810 222854
rect 347046 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 479610 222854
rect 479846 222618 510330 222854
rect 510566 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 592650 222854
rect -8726 222586 592650 222618
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 24250 219454
rect 24486 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 54970 219454
rect 55206 219218 85690 219454
rect 85926 219218 116410 219454
rect 116646 219218 147130 219454
rect 147366 219218 177850 219454
rect 178086 219218 208570 219454
rect 208806 219218 239290 219454
rect 239526 219218 270010 219454
rect 270246 219218 300730 219454
rect 300966 219218 331450 219454
rect 331686 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 464250 219454
rect 464486 219218 494970 219454
rect 495206 219218 525690 219454
rect 525926 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 24250 219134
rect 24486 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 54970 219134
rect 55206 218898 85690 219134
rect 85926 218898 116410 219134
rect 116646 218898 147130 219134
rect 147366 218898 177850 219134
rect 178086 218898 208570 219134
rect 208806 218898 239290 219134
rect 239526 218898 270010 219134
rect 270246 218898 300730 219134
rect 300966 218898 331450 219134
rect 331686 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 464250 219134
rect 464486 218898 494970 219134
rect 495206 218898 525690 219134
rect 525926 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 209494 592650 209526
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 351866 209494
rect 352102 209258 352186 209494
rect 352422 209258 387866 209494
rect 388102 209258 388186 209494
rect 388422 209258 423866 209494
rect 424102 209258 424186 209494
rect 424422 209258 459866 209494
rect 460102 209258 460186 209494
rect 460422 209258 531866 209494
rect 532102 209258 532186 209494
rect 532422 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect -8726 209174 592650 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 351866 209174
rect 352102 208938 352186 209174
rect 352422 208938 387866 209174
rect 388102 208938 388186 209174
rect 388422 208938 423866 209174
rect 424102 208938 424186 209174
rect 424422 208938 459866 209174
rect 460102 208938 460186 209174
rect 460422 208938 531866 209174
rect 532102 208938 532186 209174
rect 532422 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect -8726 208906 592650 208938
rect -8726 205774 592650 205806
rect -8726 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 348146 205774
rect 348382 205538 348466 205774
rect 348702 205538 384146 205774
rect 384382 205538 384466 205774
rect 384702 205538 420146 205774
rect 420382 205538 420466 205774
rect 420702 205538 456146 205774
rect 456382 205538 456466 205774
rect 456702 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 592650 205774
rect -8726 205454 592650 205538
rect -8726 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 348146 205454
rect 348382 205218 348466 205454
rect 348702 205218 384146 205454
rect 384382 205218 384466 205454
rect 384702 205218 420146 205454
rect 420382 205218 420466 205454
rect 420702 205218 456146 205454
rect 456382 205218 456466 205454
rect 456702 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 592650 205454
rect -8726 205186 592650 205218
rect -8726 202054 592650 202086
rect -8726 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 344426 202054
rect 344662 201818 344746 202054
rect 344982 201818 380426 202054
rect 380662 201818 380746 202054
rect 380982 201818 416426 202054
rect 416662 201818 416746 202054
rect 416982 201818 452426 202054
rect 452662 201818 452746 202054
rect 452982 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 592650 202054
rect -8726 201734 592650 201818
rect -8726 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 344426 201734
rect 344662 201498 344746 201734
rect 344982 201498 380426 201734
rect 380662 201498 380746 201734
rect 380982 201498 416426 201734
rect 416662 201498 416746 201734
rect 416982 201498 452426 201734
rect 452662 201498 452746 201734
rect 452982 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 592650 201734
rect -8726 201466 592650 201498
rect -8726 198334 592650 198366
rect -8726 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 376706 198334
rect 376942 198098 377026 198334
rect 377262 198098 412706 198334
rect 412942 198098 413026 198334
rect 413262 198098 448706 198334
rect 448942 198098 449026 198334
rect 449262 198098 484706 198334
rect 484942 198098 485026 198334
rect 485262 198098 520706 198334
rect 520942 198098 521026 198334
rect 521262 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 592650 198334
rect -8726 198014 592650 198098
rect -8726 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 376706 198014
rect 376942 197778 377026 198014
rect 377262 197778 412706 198014
rect 412942 197778 413026 198014
rect 413262 197778 448706 198014
rect 448942 197778 449026 198014
rect 449262 197778 484706 198014
rect 484942 197778 485026 198014
rect 485262 197778 520706 198014
rect 520942 197778 521026 198014
rect 521262 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 592650 198014
rect -8726 197746 592650 197778
rect -8726 194614 592650 194646
rect -8726 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 592650 194294
rect -8726 194026 592650 194058
rect -8726 190894 592650 190926
rect -8726 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 592650 190894
rect -8726 190574 592650 190658
rect -8726 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 592650 190574
rect -8726 190306 592650 190338
rect -8726 187174 592650 187206
rect -8726 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 39610 187174
rect 39846 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 70330 187174
rect 70566 186938 101050 187174
rect 101286 186938 131770 187174
rect 132006 186938 162490 187174
rect 162726 186938 193210 187174
rect 193446 186938 223930 187174
rect 224166 186938 254650 187174
rect 254886 186938 285370 187174
rect 285606 186938 316090 187174
rect 316326 186938 346810 187174
rect 347046 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 592650 187174
rect -8726 186854 592650 186938
rect -8726 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 39610 186854
rect 39846 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 70330 186854
rect 70566 186618 101050 186854
rect 101286 186618 131770 186854
rect 132006 186618 162490 186854
rect 162726 186618 193210 186854
rect 193446 186618 223930 186854
rect 224166 186618 254650 186854
rect 254886 186618 285370 186854
rect 285606 186618 316090 186854
rect 316326 186618 346810 186854
rect 347046 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 592650 186854
rect -8726 186586 592650 186618
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 24250 183454
rect 24486 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 54970 183454
rect 55206 183218 85690 183454
rect 85926 183218 116410 183454
rect 116646 183218 147130 183454
rect 147366 183218 177850 183454
rect 178086 183218 208570 183454
rect 208806 183218 239290 183454
rect 239526 183218 270010 183454
rect 270246 183218 300730 183454
rect 300966 183218 331450 183454
rect 331686 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 24250 183134
rect 24486 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 54970 183134
rect 55206 182898 85690 183134
rect 85926 182898 116410 183134
rect 116646 182898 147130 183134
rect 147366 182898 177850 183134
rect 178086 182898 208570 183134
rect 208806 182898 239290 183134
rect 239526 182898 270010 183134
rect 270246 182898 300730 183134
rect 300966 182898 331450 183134
rect 331686 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 173494 592650 173526
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 27866 173494
rect 28102 173258 28186 173494
rect 28422 173258 351866 173494
rect 352102 173258 352186 173494
rect 352422 173258 387866 173494
rect 388102 173258 388186 173494
rect 388422 173258 423866 173494
rect 424102 173258 424186 173494
rect 424422 173258 459866 173494
rect 460102 173258 460186 173494
rect 460422 173258 531866 173494
rect 532102 173258 532186 173494
rect 532422 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect -8726 173174 592650 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 27866 173174
rect 28102 172938 28186 173174
rect 28422 172938 351866 173174
rect 352102 172938 352186 173174
rect 352422 172938 387866 173174
rect 388102 172938 388186 173174
rect 388422 172938 423866 173174
rect 424102 172938 424186 173174
rect 424422 172938 459866 173174
rect 460102 172938 460186 173174
rect 460422 172938 531866 173174
rect 532102 172938 532186 173174
rect 532422 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect -8726 172906 592650 172938
rect -8726 169774 592650 169806
rect -8726 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 348146 169774
rect 348382 169538 348466 169774
rect 348702 169538 384146 169774
rect 384382 169538 384466 169774
rect 384702 169538 420146 169774
rect 420382 169538 420466 169774
rect 420702 169538 456146 169774
rect 456382 169538 456466 169774
rect 456702 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 592650 169774
rect -8726 169454 592650 169538
rect -8726 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 348146 169454
rect 348382 169218 348466 169454
rect 348702 169218 384146 169454
rect 384382 169218 384466 169454
rect 384702 169218 420146 169454
rect 420382 169218 420466 169454
rect 420702 169218 456146 169454
rect 456382 169218 456466 169454
rect 456702 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 592650 169454
rect -8726 169186 592650 169218
rect -8726 166054 592650 166086
rect -8726 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 344426 166054
rect 344662 165818 344746 166054
rect 344982 165818 380426 166054
rect 380662 165818 380746 166054
rect 380982 165818 416426 166054
rect 416662 165818 416746 166054
rect 416982 165818 452426 166054
rect 452662 165818 452746 166054
rect 452982 165818 488426 166054
rect 488662 165818 488746 166054
rect 488982 165818 524426 166054
rect 524662 165818 524746 166054
rect 524982 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 592650 166054
rect -8726 165734 592650 165818
rect -8726 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 344426 165734
rect 344662 165498 344746 165734
rect 344982 165498 380426 165734
rect 380662 165498 380746 165734
rect 380982 165498 416426 165734
rect 416662 165498 416746 165734
rect 416982 165498 452426 165734
rect 452662 165498 452746 165734
rect 452982 165498 488426 165734
rect 488662 165498 488746 165734
rect 488982 165498 524426 165734
rect 524662 165498 524746 165734
rect 524982 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 592650 165734
rect -8726 165466 592650 165498
rect -8726 162334 592650 162366
rect -8726 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 376706 162334
rect 376942 162098 377026 162334
rect 377262 162098 412706 162334
rect 412942 162098 413026 162334
rect 413262 162098 448706 162334
rect 448942 162098 449026 162334
rect 449262 162098 484706 162334
rect 484942 162098 485026 162334
rect 485262 162098 520706 162334
rect 520942 162098 521026 162334
rect 521262 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 592650 162334
rect -8726 162014 592650 162098
rect -8726 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 376706 162014
rect 376942 161778 377026 162014
rect 377262 161778 412706 162014
rect 412942 161778 413026 162014
rect 413262 161778 448706 162014
rect 448942 161778 449026 162014
rect 449262 161778 484706 162014
rect 484942 161778 485026 162014
rect 485262 161778 520706 162014
rect 520942 161778 521026 162014
rect 521262 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 592650 162014
rect -8726 161746 592650 161778
rect -8726 158614 592650 158646
rect -8726 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 592650 158294
rect -8726 158026 592650 158058
rect -8726 154894 592650 154926
rect -8726 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 592650 154894
rect -8726 154574 592650 154658
rect -8726 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 592650 154574
rect -8726 154306 592650 154338
rect -8726 151174 592650 151206
rect -8726 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 39610 151174
rect 39846 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 70330 151174
rect 70566 150938 101050 151174
rect 101286 150938 131770 151174
rect 132006 150938 162490 151174
rect 162726 150938 193210 151174
rect 193446 150938 223930 151174
rect 224166 150938 254650 151174
rect 254886 150938 285370 151174
rect 285606 150938 316090 151174
rect 316326 150938 346810 151174
rect 347046 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 429610 151174
rect 429846 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 592650 151174
rect -8726 150854 592650 150938
rect -8726 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 39610 150854
rect 39846 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 70330 150854
rect 70566 150618 101050 150854
rect 101286 150618 131770 150854
rect 132006 150618 162490 150854
rect 162726 150618 193210 150854
rect 193446 150618 223930 150854
rect 224166 150618 254650 150854
rect 254886 150618 285370 150854
rect 285606 150618 316090 150854
rect 316326 150618 346810 150854
rect 347046 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 429610 150854
rect 429846 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 592650 150854
rect -8726 150586 592650 150618
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 24250 147454
rect 24486 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 54970 147454
rect 55206 147218 85690 147454
rect 85926 147218 116410 147454
rect 116646 147218 147130 147454
rect 147366 147218 177850 147454
rect 178086 147218 208570 147454
rect 208806 147218 239290 147454
rect 239526 147218 270010 147454
rect 270246 147218 300730 147454
rect 300966 147218 331450 147454
rect 331686 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 414250 147454
rect 414486 147218 444970 147454
rect 445206 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 24250 147134
rect 24486 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 54970 147134
rect 55206 146898 85690 147134
rect 85926 146898 116410 147134
rect 116646 146898 147130 147134
rect 147366 146898 177850 147134
rect 178086 146898 208570 147134
rect 208806 146898 239290 147134
rect 239526 146898 270010 147134
rect 270246 146898 300730 147134
rect 300966 146898 331450 147134
rect 331686 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 414250 147134
rect 414486 146898 444970 147134
rect 445206 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 137494 592650 137526
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 27866 137494
rect 28102 137258 28186 137494
rect 28422 137258 351866 137494
rect 352102 137258 352186 137494
rect 352422 137258 387866 137494
rect 388102 137258 388186 137494
rect 388422 137258 459866 137494
rect 460102 137258 460186 137494
rect 460422 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect -8726 137174 592650 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 27866 137174
rect 28102 136938 28186 137174
rect 28422 136938 351866 137174
rect 352102 136938 352186 137174
rect 352422 136938 387866 137174
rect 388102 136938 388186 137174
rect 388422 136938 459866 137174
rect 460102 136938 460186 137174
rect 460422 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect -8726 136906 592650 136938
rect -8726 133774 592650 133806
rect -8726 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 348146 133774
rect 348382 133538 348466 133774
rect 348702 133538 384146 133774
rect 384382 133538 384466 133774
rect 384702 133538 456146 133774
rect 456382 133538 456466 133774
rect 456702 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 592650 133774
rect -8726 133454 592650 133538
rect -8726 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 348146 133454
rect 348382 133218 348466 133454
rect 348702 133218 384146 133454
rect 384382 133218 384466 133454
rect 384702 133218 456146 133454
rect 456382 133218 456466 133454
rect 456702 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 592650 133454
rect -8726 133186 592650 133218
rect -8726 130054 592650 130086
rect -8726 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 344426 130054
rect 344662 129818 344746 130054
rect 344982 129818 380426 130054
rect 380662 129818 380746 130054
rect 380982 129818 452426 130054
rect 452662 129818 452746 130054
rect 452982 129818 488426 130054
rect 488662 129818 488746 130054
rect 488982 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 592650 130054
rect -8726 129734 592650 129818
rect -8726 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 344426 129734
rect 344662 129498 344746 129734
rect 344982 129498 380426 129734
rect 380662 129498 380746 129734
rect 380982 129498 452426 129734
rect 452662 129498 452746 129734
rect 452982 129498 488426 129734
rect 488662 129498 488746 129734
rect 488982 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 592650 129734
rect -8726 129466 592650 129498
rect -8726 126334 592650 126366
rect -8726 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 376706 126334
rect 376942 126098 377026 126334
rect 377262 126098 484706 126334
rect 484942 126098 485026 126334
rect 485262 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 592650 126334
rect -8726 126014 592650 126098
rect -8726 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 376706 126014
rect 376942 125778 377026 126014
rect 377262 125778 484706 126014
rect 484942 125778 485026 126014
rect 485262 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 592650 126014
rect -8726 125746 592650 125778
rect -8726 122614 592650 122646
rect -8726 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 592650 122294
rect -8726 122026 592650 122058
rect -8726 118894 592650 118926
rect -8726 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 592650 118894
rect -8726 118574 592650 118658
rect -8726 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 592650 118574
rect -8726 118306 592650 118338
rect -8726 115174 592650 115206
rect -8726 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 39610 115174
rect 39846 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 70330 115174
rect 70566 114938 101050 115174
rect 101286 114938 131770 115174
rect 132006 114938 162490 115174
rect 162726 114938 193210 115174
rect 193446 114938 223930 115174
rect 224166 114938 254650 115174
rect 254886 114938 285370 115174
rect 285606 114938 316090 115174
rect 316326 114938 346810 115174
rect 347046 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 499610 115174
rect 499846 114938 530330 115174
rect 530566 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 592650 115174
rect -8726 114854 592650 114938
rect -8726 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 39610 114854
rect 39846 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 70330 114854
rect 70566 114618 101050 114854
rect 101286 114618 131770 114854
rect 132006 114618 162490 114854
rect 162726 114618 193210 114854
rect 193446 114618 223930 114854
rect 224166 114618 254650 114854
rect 254886 114618 285370 114854
rect 285606 114618 316090 114854
rect 316326 114618 346810 114854
rect 347046 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 499610 114854
rect 499846 114618 530330 114854
rect 530566 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 592650 114854
rect -8726 114586 592650 114618
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 24250 111454
rect 24486 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 54970 111454
rect 55206 111218 85690 111454
rect 85926 111218 116410 111454
rect 116646 111218 147130 111454
rect 147366 111218 177850 111454
rect 178086 111218 208570 111454
rect 208806 111218 239290 111454
rect 239526 111218 270010 111454
rect 270246 111218 300730 111454
rect 300966 111218 331450 111454
rect 331686 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 484250 111454
rect 484486 111218 514970 111454
rect 515206 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 24250 111134
rect 24486 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 54970 111134
rect 55206 110898 85690 111134
rect 85926 110898 116410 111134
rect 116646 110898 147130 111134
rect 147366 110898 177850 111134
rect 178086 110898 208570 111134
rect 208806 110898 239290 111134
rect 239526 110898 270010 111134
rect 270246 110898 300730 111134
rect 300966 110898 331450 111134
rect 331686 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 484250 111134
rect 484486 110898 514970 111134
rect 515206 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 101494 592650 101526
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 27866 101494
rect 28102 101258 28186 101494
rect 28422 101258 351866 101494
rect 352102 101258 352186 101494
rect 352422 101258 387866 101494
rect 388102 101258 388186 101494
rect 388422 101258 423866 101494
rect 424102 101258 424186 101494
rect 424422 101258 459866 101494
rect 460102 101258 460186 101494
rect 460422 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect -8726 101174 592650 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 27866 101174
rect 28102 100938 28186 101174
rect 28422 100938 351866 101174
rect 352102 100938 352186 101174
rect 352422 100938 387866 101174
rect 388102 100938 388186 101174
rect 388422 100938 423866 101174
rect 424102 100938 424186 101174
rect 424422 100938 459866 101174
rect 460102 100938 460186 101174
rect 460422 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect -8726 100906 592650 100938
rect -8726 97774 592650 97806
rect -8726 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 348146 97774
rect 348382 97538 348466 97774
rect 348702 97538 384146 97774
rect 384382 97538 384466 97774
rect 384702 97538 420146 97774
rect 420382 97538 420466 97774
rect 420702 97538 456146 97774
rect 456382 97538 456466 97774
rect 456702 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 592650 97774
rect -8726 97454 592650 97538
rect -8726 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 348146 97454
rect 348382 97218 348466 97454
rect 348702 97218 384146 97454
rect 384382 97218 384466 97454
rect 384702 97218 420146 97454
rect 420382 97218 420466 97454
rect 420702 97218 456146 97454
rect 456382 97218 456466 97454
rect 456702 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 592650 97454
rect -8726 97186 592650 97218
rect -8726 94054 592650 94086
rect -8726 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 344426 94054
rect 344662 93818 344746 94054
rect 344982 93818 380426 94054
rect 380662 93818 380746 94054
rect 380982 93818 416426 94054
rect 416662 93818 416746 94054
rect 416982 93818 452426 94054
rect 452662 93818 452746 94054
rect 452982 93818 488426 94054
rect 488662 93818 488746 94054
rect 488982 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 592650 94054
rect -8726 93734 592650 93818
rect -8726 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 344426 93734
rect 344662 93498 344746 93734
rect 344982 93498 380426 93734
rect 380662 93498 380746 93734
rect 380982 93498 416426 93734
rect 416662 93498 416746 93734
rect 416982 93498 452426 93734
rect 452662 93498 452746 93734
rect 452982 93498 488426 93734
rect 488662 93498 488746 93734
rect 488982 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 592650 93734
rect -8726 93466 592650 93498
rect -8726 90334 592650 90366
rect -8726 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 376706 90334
rect 376942 90098 377026 90334
rect 377262 90098 484706 90334
rect 484942 90098 485026 90334
rect 485262 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 592650 90334
rect -8726 90014 592650 90098
rect -8726 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 376706 90014
rect 376942 89778 377026 90014
rect 377262 89778 484706 90014
rect 484942 89778 485026 90014
rect 485262 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 592650 90014
rect -8726 89746 592650 89778
rect -8726 86614 592650 86646
rect -8726 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 592650 86294
rect -8726 86026 592650 86058
rect -8726 82894 592650 82926
rect -8726 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 592650 82894
rect -8726 82574 592650 82658
rect -8726 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 592650 82574
rect -8726 82306 592650 82338
rect -8726 79174 592650 79206
rect -8726 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 39610 79174
rect 39846 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 70330 79174
rect 70566 78938 101050 79174
rect 101286 78938 131770 79174
rect 132006 78938 162490 79174
rect 162726 78938 193210 79174
rect 193446 78938 223930 79174
rect 224166 78938 254650 79174
rect 254886 78938 285370 79174
rect 285606 78938 316090 79174
rect 316326 78938 346810 79174
rect 347046 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 405610 79174
rect 405846 78938 436330 79174
rect 436566 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 592650 79174
rect -8726 78854 592650 78938
rect -8726 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 39610 78854
rect 39846 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 70330 78854
rect 70566 78618 101050 78854
rect 101286 78618 131770 78854
rect 132006 78618 162490 78854
rect 162726 78618 193210 78854
rect 193446 78618 223930 78854
rect 224166 78618 254650 78854
rect 254886 78618 285370 78854
rect 285606 78618 316090 78854
rect 316326 78618 346810 78854
rect 347046 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 405610 78854
rect 405846 78618 436330 78854
rect 436566 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 592650 78854
rect -8726 78586 592650 78618
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 24250 75454
rect 24486 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 54970 75454
rect 55206 75218 85690 75454
rect 85926 75218 116410 75454
rect 116646 75218 147130 75454
rect 147366 75218 177850 75454
rect 178086 75218 208570 75454
rect 208806 75218 239290 75454
rect 239526 75218 270010 75454
rect 270246 75218 300730 75454
rect 300966 75218 331450 75454
rect 331686 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 390250 75454
rect 390486 75218 420970 75454
rect 421206 75218 451690 75454
rect 451926 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 24250 75134
rect 24486 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 54970 75134
rect 55206 74898 85690 75134
rect 85926 74898 116410 75134
rect 116646 74898 147130 75134
rect 147366 74898 177850 75134
rect 178086 74898 208570 75134
rect 208806 74898 239290 75134
rect 239526 74898 270010 75134
rect 270246 74898 300730 75134
rect 300966 74898 331450 75134
rect 331686 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 390250 75134
rect 390486 74898 420970 75134
rect 421206 74898 451690 75134
rect 451926 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 65494 592650 65526
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 27866 65494
rect 28102 65258 28186 65494
rect 28422 65258 351866 65494
rect 352102 65258 352186 65494
rect 352422 65258 459866 65494
rect 460102 65258 460186 65494
rect 460422 65258 495866 65494
rect 496102 65258 496186 65494
rect 496422 65258 531866 65494
rect 532102 65258 532186 65494
rect 532422 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect -8726 65174 592650 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 27866 65174
rect 28102 64938 28186 65174
rect 28422 64938 351866 65174
rect 352102 64938 352186 65174
rect 352422 64938 459866 65174
rect 460102 64938 460186 65174
rect 460422 64938 495866 65174
rect 496102 64938 496186 65174
rect 496422 64938 531866 65174
rect 532102 64938 532186 65174
rect 532422 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect -8726 64906 592650 64938
rect -8726 61774 592650 61806
rect -8726 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 348146 61774
rect 348382 61538 348466 61774
rect 348702 61538 384146 61774
rect 384382 61538 384466 61774
rect 384702 61538 492146 61774
rect 492382 61538 492466 61774
rect 492702 61538 528146 61774
rect 528382 61538 528466 61774
rect 528702 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 592650 61774
rect -8726 61454 592650 61538
rect -8726 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 348146 61454
rect 348382 61218 348466 61454
rect 348702 61218 384146 61454
rect 384382 61218 384466 61454
rect 384702 61218 492146 61454
rect 492382 61218 492466 61454
rect 492702 61218 528146 61454
rect 528382 61218 528466 61454
rect 528702 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 592650 61454
rect -8726 61186 592650 61218
rect -8726 58054 592650 58086
rect -8726 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 344426 58054
rect 344662 57818 344746 58054
rect 344982 57818 380426 58054
rect 380662 57818 380746 58054
rect 380982 57818 488426 58054
rect 488662 57818 488746 58054
rect 488982 57818 524426 58054
rect 524662 57818 524746 58054
rect 524982 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 592650 58054
rect -8726 57734 592650 57818
rect -8726 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 344426 57734
rect 344662 57498 344746 57734
rect 344982 57498 380426 57734
rect 380662 57498 380746 57734
rect 380982 57498 488426 57734
rect 488662 57498 488746 57734
rect 488982 57498 524426 57734
rect 524662 57498 524746 57734
rect 524982 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 592650 57734
rect -8726 57466 592650 57498
rect -8726 54334 592650 54366
rect -8726 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 52706 54334
rect 52942 54098 53026 54334
rect 53262 54098 88706 54334
rect 88942 54098 89026 54334
rect 89262 54098 124706 54334
rect 124942 54098 125026 54334
rect 125262 54098 160706 54334
rect 160942 54098 161026 54334
rect 161262 54098 196706 54334
rect 196942 54098 197026 54334
rect 197262 54098 232706 54334
rect 232942 54098 233026 54334
rect 233262 54098 268706 54334
rect 268942 54098 269026 54334
rect 269262 54098 304706 54334
rect 304942 54098 305026 54334
rect 305262 54098 340706 54334
rect 340942 54098 341026 54334
rect 341262 54098 376706 54334
rect 376942 54098 377026 54334
rect 377262 54098 484706 54334
rect 484942 54098 485026 54334
rect 485262 54098 520706 54334
rect 520942 54098 521026 54334
rect 521262 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 592650 54334
rect -8726 54014 592650 54098
rect -8726 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 52706 54014
rect 52942 53778 53026 54014
rect 53262 53778 88706 54014
rect 88942 53778 89026 54014
rect 89262 53778 124706 54014
rect 124942 53778 125026 54014
rect 125262 53778 160706 54014
rect 160942 53778 161026 54014
rect 161262 53778 196706 54014
rect 196942 53778 197026 54014
rect 197262 53778 232706 54014
rect 232942 53778 233026 54014
rect 233262 53778 268706 54014
rect 268942 53778 269026 54014
rect 269262 53778 304706 54014
rect 304942 53778 305026 54014
rect 305262 53778 340706 54014
rect 340942 53778 341026 54014
rect 341262 53778 376706 54014
rect 376942 53778 377026 54014
rect 377262 53778 484706 54014
rect 484942 53778 485026 54014
rect 485262 53778 520706 54014
rect 520942 53778 521026 54014
rect 521262 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 592650 54014
rect -8726 53746 592650 53778
rect -8726 50614 592650 50646
rect -8726 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 592650 50294
rect -8726 50026 592650 50058
rect -8726 46894 592650 46926
rect -8726 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 592650 46894
rect -8726 46574 592650 46658
rect -8726 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 592650 46574
rect -8726 46306 592650 46338
rect -8726 43174 592650 43206
rect -8726 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 405610 43174
rect 405846 42938 436330 43174
rect 436566 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545930 43174
rect 546166 42938 550875 43174
rect 551111 42938 555820 43174
rect 556056 42938 560765 43174
rect 561001 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 592650 43174
rect -8726 42854 592650 42938
rect -8726 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 405610 42854
rect 405846 42618 436330 42854
rect 436566 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545930 42854
rect 546166 42618 550875 42854
rect 551111 42618 555820 42854
rect 556056 42618 560765 42854
rect 561001 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 592650 42854
rect -8726 42586 592650 42618
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 390250 39454
rect 390486 39218 420970 39454
rect 421206 39218 451690 39454
rect 451926 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 543458 39454
rect 543694 39218 548403 39454
rect 548639 39218 553348 39454
rect 553584 39218 558293 39454
rect 558529 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 390250 39134
rect 390486 38898 420970 39134
rect 421206 38898 451690 39134
rect 451926 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 543458 39134
rect 543694 38898 548403 39134
rect 548639 38898 553348 39134
rect 553584 38898 558293 39134
rect 558529 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 29494 592650 29526
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 63866 29494
rect 64102 29258 64186 29494
rect 64422 29258 99866 29494
rect 100102 29258 100186 29494
rect 100422 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 351866 29494
rect 352102 29258 352186 29494
rect 352422 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect -8726 29174 592650 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 63866 29174
rect 64102 28938 64186 29174
rect 64422 28938 99866 29174
rect 100102 28938 100186 29174
rect 100422 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 351866 29174
rect 352102 28938 352186 29174
rect 352422 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect -8726 28906 592650 28938
rect -8726 25774 592650 25806
rect -8726 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 60146 25774
rect 60382 25538 60466 25774
rect 60702 25538 96146 25774
rect 96382 25538 96466 25774
rect 96702 25538 132146 25774
rect 132382 25538 132466 25774
rect 132702 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 348146 25774
rect 348382 25538 348466 25774
rect 348702 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 420146 25774
rect 420382 25538 420466 25774
rect 420702 25538 456146 25774
rect 456382 25538 456466 25774
rect 456702 25538 492146 25774
rect 492382 25538 492466 25774
rect 492702 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 592650 25774
rect -8726 25454 592650 25538
rect -8726 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 60146 25454
rect 60382 25218 60466 25454
rect 60702 25218 96146 25454
rect 96382 25218 96466 25454
rect 96702 25218 132146 25454
rect 132382 25218 132466 25454
rect 132702 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 348146 25454
rect 348382 25218 348466 25454
rect 348702 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 420146 25454
rect 420382 25218 420466 25454
rect 420702 25218 456146 25454
rect 456382 25218 456466 25454
rect 456702 25218 492146 25454
rect 492382 25218 492466 25454
rect 492702 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 592650 25454
rect -8726 25186 592650 25218
rect -8726 22054 592650 22086
rect -8726 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 92426 22054
rect 92662 21818 92746 22054
rect 92982 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 592650 22054
rect -8726 21734 592650 21818
rect -8726 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 92426 21734
rect 92662 21498 92746 21734
rect 92982 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 592650 21734
rect -8726 21466 592650 21498
rect -8726 18334 592650 18366
rect -8726 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 592650 18334
rect -8726 18014 592650 18098
rect -8726 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 592650 18014
rect -8726 17746 592650 17778
rect -8726 14614 592650 14646
rect -8726 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 592650 14294
rect -8726 14026 592650 14058
rect -8726 10894 592650 10926
rect -8726 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 592650 10894
rect -8726 10574 592650 10658
rect -8726 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 592650 10574
rect -8726 10306 592650 10338
rect -8726 7174 592650 7206
rect -8726 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 592650 7174
rect -8726 6854 592650 6938
rect -8726 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 592650 6854
rect -8726 6586 592650 6618
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 60146 -6106
rect 60382 -6342 60466 -6106
rect 60702 -6342 96146 -6106
rect 96382 -6342 96466 -6106
rect 96702 -6342 132146 -6106
rect 132382 -6342 132466 -6106
rect 132702 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 60146 -6426
rect 60382 -6662 60466 -6426
rect 60702 -6662 96146 -6426
rect 96382 -6662 96466 -6426
rect 96702 -6662 132146 -6426
rect 132382 -6662 132466 -6426
rect 132702 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 63866 -7066
rect 64102 -7302 64186 -7066
rect 64422 -7302 99866 -7066
rect 100102 -7302 100186 -7066
rect 100422 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 63866 -7386
rect 64102 -7622 64186 -7386
rect 64422 -7622 99866 -7386
rect 100102 -7622 100186 -7386
rect 100422 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use posit_unit  posit_unit
timestamp 0
transform 1 0 460000 0 1 200000
box 0 2128 70000 67504
use multiplexer  proj_multiplexer
timestamp 0
transform 1 0 450000 0 1 322000
box 0 0 60000 64000
use tholin_avalonsemi_5401  tholin_avalonsemi_5401
timestamp 0
transform 1 0 520000 0 1 425000
box 1066 0 36000 36000
use tholin_avalonsemi_tbb1143  tholin_avalonsemi_tbb1143
timestamp 0
transform 1 0 400000 0 1 305000
box 1066 2048 30000 30000
use tt2_tholin_diceroll  tt2_tholin_diceroll
timestamp 0
transform 1 0 470000 0 1 432000
box 1066 0 21043 22000
use tt2_tholin_multiplexed_counter  tt2_tholin_multiplexed_counter
timestamp 0
transform 1 0 550000 0 1 360000
box 842 0 17098 18000
use tt2_tholin_multiplier  tt2_tholin_multiplier
timestamp 0
transform 1 0 450000 0 1 500000
box 0 0 11118 16584
use tt2_tholin_namebadge  tt2_tholin_namebadge
timestamp 0
transform 1 0 420000 0 1 420000
box 1066 0 23987 25000
use tune_player  tune_player
timestamp 0
transform 1 0 540000 0 1 30000
box 0 2128 21043 19632
use wrapped_6502  wrapped_6502
timestamp 0
transform 1 0 410000 0 1 120000
box 1066 1504 40000 40000
use wrapped_MC14500  wrapped_MC14500
timestamp 0
transform 1 0 480000 0 1 500000
box 566 0 12000 18000
use wrapped_as1802  wrapped_as1802
timestamp 0
transform 1 0 480000 0 1 80000
box 1066 2128 60000 60000
use wrapped_as2650  wrapped_as2650
timestamp 0
transform 1 0 460000 0 1 600000
box 0 0 68816 67992
use wrapped_as512512512  wrapped_as512512512
timestamp 0
transform 1 0 20000 0 1 45000
box 1066 2128 340000 637616
use wrapped_vgatest  wrapped_vgatest
timestamp 0
transform 1 0 386000 0 1 30000
box 749 2128 75000 75000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 56303 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 680513 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 56303 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 680513 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 56303 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 680513 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 56303 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 680513 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 56303 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 680513 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 56303 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 680513 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 56303 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 680513 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 56303 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 680513 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 31919 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 92137 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 31919 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 161465 434414 420423 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 443377 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 201919 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 385580 470414 600287 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 668801 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 83687 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 139417 506414 201919 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 259417 506414 600287 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 668801 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 425068 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 460836 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 9234 -7654 9854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 -7654 45854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 -7654 81854 56303 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 680513 81854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 -7654 117854 56303 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 680513 117854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 -7654 153854 56303 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 680513 153854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 -7654 189854 56303 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 680513 189854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 -7654 225854 56303 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 680513 225854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 -7654 261854 56303 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 680513 261854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 -7654 297854 56303 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 680513 297854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 -7654 333854 56303 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 680513 333854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 369234 -7654 369854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 -7654 405854 30068 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 104460 405854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 -7654 441854 31919 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 161465 441854 420423 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 443377 441854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 -7654 477854 201919 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 259417 477854 320655 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 385225 477854 600287 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 668801 477854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 -7654 513854 83687 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 139417 513854 201919 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 259417 513854 600287 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 668801 513854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 -7654 549854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 10306 592650 10926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 46306 592650 46926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 82306 592650 82926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 118306 592650 118926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 154306 592650 154926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 190306 592650 190926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 226306 592650 226926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 262306 592650 262926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 298306 592650 298926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 334306 592650 334926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 370306 592650 370926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 406306 592650 406926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 442306 592650 442926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 478306 592650 478926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 514306 592650 514926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 550306 592650 550926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 586306 592650 586926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 622306 592650 622926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 658306 592650 658926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 694306 592650 694926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 16674 -7654 17294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 52674 -7654 53294 56303 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 -7654 89294 56303 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 124674 -7654 125294 56303 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 160674 -7654 161294 56303 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 196674 -7654 197294 56303 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 232674 -7654 233294 56303 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 268674 -7654 269294 56303 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 304674 -7654 305294 56303 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 340674 -7654 341294 56303 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 376674 -7654 377294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 412674 -7654 413294 31919 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 412674 161465 413294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 -7654 449294 31919 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 161465 449294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 -7654 485294 201919 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 259417 485294 320655 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 385580 485294 500068 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 517884 485294 600287 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 -7654 521294 83687 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 139417 521294 201919 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 259417 521294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 556674 -7654 557294 360068 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 556674 377884 557294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 17746 592650 18366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 53746 592650 54366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 89746 592650 90366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 125746 592650 126366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 161746 592650 162366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 197746 592650 198366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 233746 592650 234366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 269746 592650 270366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 305746 592650 306366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 341746 592650 342366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 377746 592650 378366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 413746 592650 414366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 449746 592650 450366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 485746 592650 486366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 521746 592650 522366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 557746 592650 558366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 593746 592650 594366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 629746 592650 630366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 665746 592650 666366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 24114 -7654 24734 45068 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 60114 -7654 60734 56303 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 96114 -7654 96734 56303 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 132114 -7654 132734 56303 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 168114 -7654 168734 56303 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 204114 -7654 204734 56303 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 240114 -7654 240734 56303 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 276114 -7654 276734 56303 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 312114 -7654 312734 56303 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 348114 -7654 348734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 384114 -7654 384734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 -7654 420734 31919 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 92137 420734 120423 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 161465 420734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 -7654 456734 31919 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 92137 456734 500068 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 517884 456734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 -7654 492734 83687 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 259417 492734 320655 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 385225 492734 600287 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 668801 492734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 -7654 528734 83687 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 259417 528734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 564114 -7654 564734 360068 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 564114 377884 564734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 25186 592650 25806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 61186 592650 61806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 97186 592650 97806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 133186 592650 133806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 169186 592650 169806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 205186 592650 205806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 241186 592650 241806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 277186 592650 277806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 313186 592650 313806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 349186 592650 349806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 385186 592650 385806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 421186 592650 421806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 457186 592650 457806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 493186 592650 493806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 529186 592650 529806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 565186 592650 565806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 601186 592650 601806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 637186 592650 637806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 673186 592650 673806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 20394 -7654 21014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 56394 -7654 57014 56303 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 -7654 93014 56303 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 128394 -7654 129014 56303 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 164394 -7654 165014 56303 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 200394 -7654 201014 56303 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 236394 -7654 237014 56303 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272394 -7654 273014 56303 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 308394 -7654 309014 56303 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 344394 -7654 345014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 380394 -7654 381014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 -7654 417014 31919 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 92137 417014 120423 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 161465 417014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 -7654 453014 31919 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 92137 453014 500068 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 517884 453014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 -7654 489014 201919 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 259417 489014 320655 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 453692 489014 500068 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 517884 489014 600287 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 668801 489014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 -7654 525014 83687 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 139417 525014 201919 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 259417 525014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560394 -7654 561014 30068 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560394 51692 561014 360068 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560394 377884 561014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 21466 592650 22086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 57466 592650 58086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 93466 592650 94086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 129466 592650 130086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 165466 592650 166086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 201466 592650 202086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 237466 592650 238086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 273466 592650 274086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 309466 592650 310086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 345466 592650 346086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 381466 592650 382086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 417466 592650 418086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 453466 592650 454086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 489466 592650 490086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 525466 592650 526086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 561466 592650 562086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 597466 592650 598086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 633466 592650 634086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 669466 592650 670086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 27834 -7654 28454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 63834 -7654 64454 56303 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 -7654 100454 56303 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 135834 -7654 136454 56303 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 171834 -7654 172454 56303 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 207834 -7654 208454 56303 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 243834 -7654 244454 56303 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 279834 -7654 280454 56303 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 315834 -7654 316454 45068 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 351834 -7654 352454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 387834 -7654 388454 31919 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 387834 92137 388454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 -7654 424454 31919 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 92137 424454 120423 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 161465 424454 420068 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 444412 424454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 -7654 460454 500068 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 517884 460454 600287 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 668801 460454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 -7654 496454 83687 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 259417 496454 320655 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 385225 496454 600287 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 668801 496454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 -7654 532454 83687 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 139417 532454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 567834 -7654 568454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 28906 592650 29526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 64906 592650 65526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 100906 592650 101526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 136906 592650 137526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 172906 592650 173526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 208906 592650 209526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 244906 592650 245526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 280906 592650 281526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 316906 592650 317526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 352906 592650 353526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 388906 592650 389526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 424906 592650 425526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 460906 592650 461526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 496906 592650 497526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 532906 592650 533526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 568906 592650 569526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 604906 592650 605526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 640906 592650 641526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 676906 592650 677526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 5514 -7654 6134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 -7654 42134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 -7654 78134 56303 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 680513 78134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 -7654 114134 56303 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 680513 114134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 -7654 150134 56303 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 680513 150134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 -7654 186134 56303 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 680513 186134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 -7654 222134 56303 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 680513 222134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 -7654 258134 56303 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 680513 258134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 -7654 294134 56303 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 680513 294134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 -7654 330134 56303 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 680513 330134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 -7654 366134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 -7654 402134 31919 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 92137 402134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 -7654 438134 31919 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 161465 438134 420068 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 444412 438134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 -7654 474134 201919 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 453692 474134 600287 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 668801 474134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 -7654 510134 83687 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 139417 510134 201919 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 259417 510134 600287 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 668801 510134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 -7654 546134 30068 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 51692 546134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 581514 -7654 582134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 6586 592650 7206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 42586 592650 43206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 78586 592650 79206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 114586 592650 115206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 150586 592650 151206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 186586 592650 187206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 222586 592650 223206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 258586 592650 259206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 294586 592650 295206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 330586 592650 331206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 366586 592650 367206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 402586 592650 403206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 438586 592650 439206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 474586 592650 475206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 510586 592650 511206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 546586 592650 547206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 582586 592650 583206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 618586 592650 619206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 654586 592650 655206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 690586 592650 691206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 12954 -7654 13574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 -7654 49574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 -7654 85574 56303 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 680513 85574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 -7654 121574 56303 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 680513 121574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 -7654 157574 56303 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 680513 157574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 -7654 193574 45068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 684676 193574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 -7654 229574 56303 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 680513 229574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 -7654 265574 56303 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 680513 265574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 -7654 301574 45068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 684676 301574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 -7654 337574 56303 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 680513 337574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 372954 -7654 373574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 -7654 409574 31919 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 92137 409574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 -7654 445574 31919 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 161465 445574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 -7654 481574 201919 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 259417 481574 320655 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 453692 481574 600287 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 668801 481574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 -7654 517574 83687 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 139417 517574 201919 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 259417 517574 600287 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 668801 517574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 -7654 553574 30068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 51692 553574 360068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 377884 553574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 14026 592650 14646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 50026 592650 50646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 86026 592650 86646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 122026 592650 122646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 158026 592650 158646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 194026 592650 194646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 230026 592650 230646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 266026 592650 266646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 302026 592650 302646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 338026 592650 338646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 374026 592650 374646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 410026 592650 410646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 446026 592650 446646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 482026 592650 482646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 518026 592650 518646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 554026 592650 554646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 590026 592650 590646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 626026 592650 626646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 662026 592650 662646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 698026 592650 698646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
rlabel via4 451808 75336 451808 75336 0 vccd1
rlabel via4 333704 46776 333704 46776 0 vccd2
rlabel via4 341144 54216 341144 54216 0 vdda1
rlabel via4 456584 97656 456584 97656 0 vdda2
rlabel via4 452864 93936 452864 93936 0 vssa1
rlabel via4 460304 101376 460304 101376 0 vssa2
rlabel via4 436448 79056 436448 79056 0 vssd1
rlabel via4 337424 50496 337424 50496 0 vssd2
rlabel metal2 422655 444380 422655 444380 0 design_clk
rlabel metal2 411578 159868 411578 159868 0 dsi_all\[0\]
rlabel metal1 445004 330582 445004 330582 0 dsi_all\[10\]
rlabel metal2 447258 331415 447258 331415 0 dsi_all\[11\]
rlabel metal3 448876 332180 448876 332180 0 dsi_all\[12\]
rlabel metal2 447258 332741 447258 332741 0 dsi_all\[13\]
rlabel metal2 447350 333115 447350 333115 0 dsi_all\[14\]
rlabel metal2 447258 334101 447258 334101 0 dsi_all\[15\]
rlabel metal1 445510 334050 445510 334050 0 dsi_all\[16\]
rlabel metal1 444820 335478 444820 335478 0 dsi_all\[17\]
rlabel metal2 447258 335835 447258 335835 0 dsi_all\[18\]
rlabel metal2 447166 336889 447166 336889 0 dsi_all\[19\]
rlabel metal3 450156 503423 450156 503423 0 dsi_all\[1\]
rlabel metal2 447258 337195 447258 337195 0 dsi_all\[20\]
rlabel metal2 431250 310522 431250 310522 0 dsi_all\[21\]
rlabel metal2 385986 316030 385986 316030 0 dsi_all\[22\]
rlabel metal1 445510 339558 445510 339558 0 dsi_all\[23\]
rlabel metal2 447166 339915 447166 339915 0 dsi_all\[24\]
rlabel metal2 442934 338504 442934 338504 0 dsi_all\[25\]
rlabel metal2 447166 341309 447166 341309 0 dsi_all\[26\]
rlabel metal3 449612 342380 449612 342380 0 dsi_all\[27\]
rlabel metal3 450156 505395 450156 505395 0 dsi_all\[2\]
rlabel metal2 447258 326553 447258 326553 0 dsi_all\[3\]
rlabel metal2 425040 160011 425040 160011 0 dsi_all\[4\]
rlabel metal2 428184 159868 428184 159868 0 dsi_all\[5\]
rlabel metal2 431496 159868 431496 159868 0 dsi_all\[6\]
rlabel metal3 448692 328780 448692 328780 0 dsi_all\[7\]
rlabel metal2 447258 329613 447258 329613 0 dsi_all\[8\]
rlabel metal3 448692 330140 448692 330140 0 dsi_all\[9\]
rlabel metal2 487002 320120 487002 320120 0 dso_6502\[0\]
rlabel metal2 489762 297340 489762 297340 0 dso_6502\[10\]
rlabel via2 451582 136493 451582 136493 0 dso_6502\[11\]
rlabel via2 452594 137853 452594 137853 0 dso_6502\[12\]
rlabel metal3 449788 139313 449788 139313 0 dso_6502\[13\]
rlabel metal3 449788 140673 449788 140673 0 dso_6502\[14\]
rlabel metal3 449788 142033 449788 142033 0 dso_6502\[15\]
rlabel metal3 449788 143393 449788 143393 0 dso_6502\[16\]
rlabel metal3 449788 144753 449788 144753 0 dso_6502\[17\]
rlabel metal3 449788 146113 449788 146113 0 dso_6502\[18\]
rlabel metal3 449788 147473 449788 147473 0 dso_6502\[19\]
rlabel metal3 449788 123265 449788 123265 0 dso_6502\[1\]
rlabel metal3 449788 148901 449788 148901 0 dso_6502\[20\]
rlabel metal3 449788 150261 449788 150261 0 dso_6502\[21\]
rlabel metal3 449788 151621 449788 151621 0 dso_6502\[22\]
rlabel metal3 449788 152981 449788 152981 0 dso_6502\[23\]
rlabel metal3 449788 154273 449788 154273 0 dso_6502\[24\]
rlabel metal3 449788 155701 449788 155701 0 dso_6502\[25\]
rlabel metal3 449788 157129 449788 157129 0 dso_6502\[26\]
rlabel metal3 449788 124625 449788 124625 0 dso_6502\[2\]
rlabel metal3 449788 125985 449788 125985 0 dso_6502\[3\]
rlabel metal2 488106 298700 488106 298700 0 dso_6502\[4\]
rlabel metal2 488382 315972 488382 315972 0 dso_6502\[5\]
rlabel metal2 488658 315292 488658 315292 0 dso_6502\[6\]
rlabel metal2 488934 307710 488934 307710 0 dso_6502\[7\]
rlabel metal2 489210 320086 489210 320086 0 dso_6502\[8\]
rlabel metal2 489486 299448 489486 299448 0 dso_6502\[9\]
rlabel metal2 503785 385900 503785 385900 0 dso_LCD\[0\]
rlabel metal2 504337 385900 504337 385900 0 dso_LCD\[1\]
rlabel metal2 505310 387862 505310 387862 0 dso_LCD\[2\]
rlabel metal2 506046 388576 506046 388576 0 dso_LCD\[3\]
rlabel metal2 506683 385900 506683 385900 0 dso_LCD\[4\]
rlabel metal2 507327 385900 507327 385900 0 dso_LCD\[5\]
rlabel metal2 508109 385900 508109 385900 0 dso_LCD\[6\]
rlabel metal2 508799 385900 508799 385900 0 dso_LCD\[7\]
rlabel metal3 540492 82348 540492 82348 0 dso_as1802\[0\]
rlabel metal3 540538 102748 540538 102748 0 dso_as1802\[10\]
rlabel metal3 540676 104788 540676 104788 0 dso_as1802\[11\]
rlabel metal3 540722 106828 540722 106828 0 dso_as1802\[12\]
rlabel via2 539925 109140 539925 109140 0 dso_as1802\[13\]
rlabel metal3 540584 110908 540584 110908 0 dso_as1802\[14\]
rlabel metal3 539948 112865 539948 112865 0 dso_as1802\[15\]
rlabel metal3 540768 114988 540768 114988 0 dso_as1802\[16\]
rlabel metal3 539948 117179 539948 117179 0 dso_as1802\[17\]
rlabel metal3 541504 119068 541504 119068 0 dso_as1802\[18\]
rlabel metal3 541228 121108 541228 121108 0 dso_as1802\[19\]
rlabel metal3 541274 84388 541274 84388 0 dso_as1802\[1\]
rlabel metal2 499974 296048 499974 296048 0 dso_as1802\[20\]
rlabel metal2 500250 295300 500250 295300 0 dso_as1802\[21\]
rlabel metal2 500526 296082 500526 296082 0 dso_as1802\[22\]
rlabel metal2 500802 318029 500802 318029 0 dso_as1802\[23\]
rlabel metal2 501078 318828 501078 318828 0 dso_as1802\[24\]
rlabel metal3 540170 133348 540170 133348 0 dso_as1802\[25\]
rlabel metal2 539258 135660 539258 135660 0 dso_as1802\[26\]
rlabel via2 539741 86836 539741 86836 0 dso_as1802\[2\]
rlabel metal3 540630 88468 540630 88468 0 dso_as1802\[3\]
rlabel metal3 541320 90508 541320 90508 0 dso_as1802\[4\]
rlabel metal3 541412 92548 541412 92548 0 dso_as1802\[5\]
rlabel metal3 541596 94588 541596 94588 0 dso_as1802\[6\]
rlabel metal3 541458 96628 541458 96628 0 dso_as1802\[7\]
rlabel via2 539603 99212 539603 99212 0 dso_as1802\[8\]
rlabel via2 539787 100572 539787 100572 0 dso_as1802\[9\]
rlabel metal2 463121 385900 463121 385900 0 dso_as2650\[0\]
rlabel metal3 459824 626280 459824 626280 0 dso_as2650\[10\]
rlabel metal2 471217 385900 471217 385900 0 dso_as2650\[11\]
rlabel metal2 472190 388559 472190 388559 0 dso_as2650\[12\]
rlabel metal2 472926 387471 472926 387471 0 dso_as2650\[13\]
rlabel metal3 459747 635460 459747 635460 0 dso_as2650\[14\]
rlabel metal3 459793 637908 459793 637908 0 dso_as2650\[15\]
rlabel metal3 459517 640356 459517 640356 0 dso_as2650\[16\]
rlabel metal2 468510 493544 468510 493544 0 dso_as2650\[17\]
rlabel metal1 458896 603738 458896 603738 0 dso_as2650\[18\]
rlabel metal2 469982 494258 469982 494258 0 dso_as2650\[19\]
rlabel metal2 463903 385900 463903 385900 0 dso_as2650\[1\]
rlabel metal2 469890 494190 469890 494190 0 dso_as2650\[20\]
rlabel metal2 461610 494394 461610 494394 0 dso_as2650\[21\]
rlabel metal3 459640 655724 459640 655724 0 dso_as2650\[22\]
rlabel metal2 480286 387182 480286 387182 0 dso_as2650\[23\]
rlabel metal2 481022 387250 481022 387250 0 dso_as2650\[24\]
rlabel metal2 481758 387352 481758 387352 0 dso_as2650\[25\]
rlabel metal2 482494 387284 482494 387284 0 dso_as2650\[26\]
rlabel metal2 464593 385900 464593 385900 0 dso_as2650\[2\]
rlabel metal2 465375 385900 465375 385900 0 dso_as2650\[3\]
rlabel metal2 466111 385900 466111 385900 0 dso_as2650\[4\]
rlabel metal2 466755 385900 466755 385900 0 dso_as2650\[5\]
rlabel metal2 467537 385900 467537 385900 0 dso_as2650\[6\]
rlabel metal2 468273 385900 468273 385900 0 dso_as2650\[7\]
rlabel metal2 469246 386978 469246 386978 0 dso_as2650\[8\]
rlabel metal2 469982 386944 469982 386944 0 dso_as2650\[9\]
rlabel metal2 429226 367778 429226 367778 0 dso_as512512512\[0\]
rlabel metal2 447258 372045 447258 372045 0 dso_as512512512\[10\]
rlabel metal2 447166 372419 447166 372419 0 dso_as512512512\[11\]
rlabel metal2 447258 373439 447258 373439 0 dso_as512512512\[12\]
rlabel metal2 447166 373813 447166 373813 0 dso_as512512512\[13\]
rlabel metal2 411930 449854 411930 449854 0 dso_as512512512\[14\]
rlabel metal2 447166 375173 447166 375173 0 dso_as512512512\[15\]
rlabel metal2 447258 376193 447258 376193 0 dso_as512512512\[16\]
rlabel metal2 447166 376499 447166 376499 0 dso_as512512512\[17\]
rlabel metal2 367770 473348 367770 473348 0 dso_as512512512\[18\]
rlabel metal2 370530 478856 370530 478856 0 dso_as512512512\[19\]
rlabel metal1 444820 365602 444820 365602 0 dso_as512512512\[1\]
rlabel metal2 372002 485078 372002 485078 0 dso_as512512512\[20\]
rlabel metal2 447166 379253 447166 379253 0 dso_as512512512\[21\]
rlabel metal2 410550 496774 410550 496774 0 dso_as512512512\[22\]
rlabel metal2 447166 380647 447166 380647 0 dso_as512512512\[23\]
rlabel metal2 407790 508470 407790 508470 0 dso_as512512512\[24\]
rlabel metal2 447166 382007 447166 382007 0 dso_as512512512\[25\]
rlabel metal2 406410 520234 406410 520234 0 dso_as512512512\[26\]
rlabel metal2 447166 383401 447166 383401 0 dso_as512512512\[27\]
rlabel metal2 447166 366605 447166 366605 0 dso_as512512512\[2\]
rlabel metal1 444774 366962 444774 366962 0 dso_as512512512\[3\]
rlabel metal2 447258 367999 447258 367999 0 dso_as512512512\[4\]
rlabel metal2 447166 368305 447166 368305 0 dso_as512512512\[5\]
rlabel metal2 447258 369359 447258 369359 0 dso_as512512512\[6\]
rlabel metal2 447166 369665 447166 369665 0 dso_as512512512\[7\]
rlabel metal2 447258 370719 447258 370719 0 dso_as512512512\[8\]
rlabel metal2 447166 371025 447166 371025 0 dso_as512512512\[9\]
rlabel metal2 483177 385900 483177 385900 0 dso_as5401\[0\]
rlabel metal2 490590 389256 490590 389256 0 dso_as5401\[10\]
rlabel metal2 491326 387607 491326 387607 0 dso_as5401\[11\]
rlabel metal2 491825 385900 491825 385900 0 dso_as5401\[12\]
rlabel metal2 537779 425068 537779 425068 0 dso_as5401\[13\]
rlabel metal2 539067 425068 539067 425068 0 dso_as5401\[14\]
rlabel metal2 540355 425068 540355 425068 0 dso_as5401\[15\]
rlabel metal2 541834 422630 541834 422630 0 dso_as5401\[16\]
rlabel metal2 542931 425068 542931 425068 0 dso_as5401\[17\]
rlabel metal2 544219 425068 544219 425068 0 dso_as5401\[18\]
rlabel metal2 545698 424092 545698 424092 0 dso_as5401\[19\]
rlabel metal2 483775 385900 483775 385900 0 dso_as5401\[1\]
rlabel metal2 546795 425068 546795 425068 0 dso_as5401\[20\]
rlabel metal2 498449 385900 498449 385900 0 dso_as5401\[21\]
rlabel metal2 522330 406130 522330 406130 0 dso_as5401\[22\]
rlabel metal2 499921 385900 499921 385900 0 dso_as5401\[23\]
rlabel metal2 500894 387386 500894 387386 0 dso_as5401\[24\]
rlabel metal2 501393 385900 501393 385900 0 dso_as5401\[25\]
rlabel metal2 502366 387318 502366 387318 0 dso_as5401\[26\]
rlabel metal2 484702 387420 484702 387420 0 dso_as5401\[2\]
rlabel metal2 485438 387284 485438 387284 0 dso_as5401\[3\]
rlabel metal2 485983 385900 485983 385900 0 dso_as5401\[4\]
rlabel metal2 486910 387250 486910 387250 0 dso_as5401\[5\]
rlabel metal2 487409 385900 487409 385900 0 dso_as5401\[6\]
rlabel metal2 488382 387182 488382 387182 0 dso_as5401\[7\]
rlabel metal2 488881 385900 488881 385900 0 dso_as5401\[8\]
rlabel metal2 489854 387216 489854 387216 0 dso_as5401\[9\]
rlabel metal2 522330 368628 522330 368628 0 dso_counter\[0\]
rlabel metal2 547170 371348 547170 371348 0 dso_counter\[10\]
rlabel metal2 567042 359458 567042 359458 0 dso_counter\[11\]
rlabel metal3 511650 379236 511650 379236 0 dso_counter\[1\]
rlabel metal2 544410 369308 544410 369308 0 dso_counter\[2\]
rlabel metal3 511052 380324 511052 380324 0 dso_counter\[3\]
rlabel metal3 511420 380868 511420 380868 0 dso_counter\[4\]
rlabel metal2 558210 359594 558210 359594 0 dso_counter\[5\]
rlabel metal2 547262 367268 547262 367268 0 dso_counter\[6\]
rlabel metal2 561154 359254 561154 359254 0 dso_counter\[7\]
rlabel metal2 562626 359356 562626 359356 0 dso_counter\[8\]
rlabel metal2 519662 370498 519662 370498 0 dso_counter\[9\]
rlabel metal2 456734 387182 456734 387182 0 dso_diceroll\[0\]
rlabel metal2 457233 385900 457233 385900 0 dso_diceroll\[1\]
rlabel metal2 458206 389290 458206 389290 0 dso_diceroll\[2\]
rlabel metal2 458705 385900 458705 385900 0 dso_diceroll\[3\]
rlabel metal2 461702 388858 461702 388858 0 dso_diceroll\[4\]
rlabel metal1 483644 429182 483644 429182 0 dso_diceroll\[5\]
rlabel metal2 461150 389256 461150 389256 0 dso_diceroll\[6\]
rlabel metal2 461649 385900 461649 385900 0 dso_diceroll\[7\]
rlabel via2 450317 352988 450317 352988 0 dso_mc14500\[0\]
rlabel metal3 448922 353260 448922 353260 0 dso_mc14500\[1\]
rlabel metal3 449934 353940 449934 353940 0 dso_mc14500\[2\]
rlabel metal3 449888 354620 449888 354620 0 dso_mc14500\[3\]
rlabel metal2 484902 500140 484902 500140 0 dso_mc14500\[4\]
rlabel metal2 486420 500140 486420 500140 0 dso_mc14500\[5\]
rlabel metal2 487478 500140 487478 500140 0 dso_mc14500\[6\]
rlabel metal2 488812 500140 488812 500140 0 dso_mc14500\[7\]
rlabel metal3 449566 358020 449566 358020 0 dso_mc14500\[8\]
rlabel metal2 450793 385900 450793 385900 0 dso_multiplier\[0\]
rlabel metal2 451437 385900 451437 385900 0 dso_multiplier\[1\]
rlabel metal2 452081 385900 452081 385900 0 dso_multiplier\[2\]
rlabel metal2 452955 385900 452955 385900 0 dso_multiplier\[3\]
rlabel metal2 453790 387522 453790 387522 0 dso_multiplier\[4\]
rlabel metal2 454335 385900 454335 385900 0 dso_multiplier\[5\]
rlabel metal2 455071 385900 455071 385900 0 dso_multiplier\[6\]
rlabel metal2 461058 498552 461058 498552 0 dso_multiplier\[7\]
rlabel metal2 485622 318012 485622 318012 0 dso_posit\[0\]
rlabel metal2 485898 312844 485898 312844 0 dso_posit\[1\]
rlabel metal2 486174 303528 486174 303528 0 dso_posit\[2\]
rlabel metal2 486450 311858 486450 311858 0 dso_posit\[3\]
rlabel metal2 447166 359091 447166 359091 0 dso_tbb1143\[0\]
rlabel metal1 444820 358870 444820 358870 0 dso_tbb1143\[1\]
rlabel metal2 447166 360519 447166 360519 0 dso_tbb1143\[2\]
rlabel metal2 447258 360825 447258 360825 0 dso_tbb1143\[3\]
rlabel metal2 447166 361845 447166 361845 0 dso_tbb1143\[4\]
rlabel metal1 444774 361658 444774 361658 0 dso_tbb1143\[5\]
rlabel metal2 447166 363239 447166 363239 0 dso_tbb1143\[6\]
rlabel metal2 447258 363545 447258 363545 0 dso_tbb1143\[7\]
rlabel metal2 502182 320766 502182 320766 0 dso_tune
rlabel metal2 502458 319440 502458 319440 0 dso_vgatest\[0\]
rlabel metal2 407806 104924 407806 104924 0 dso_vgatest\[1\]
rlabel metal2 503010 319406 503010 319406 0 dso_vgatest\[2\]
rlabel metal2 450846 188496 450846 188496 0 dso_vgatest\[3\]
rlabel metal2 426680 104924 426680 104924 0 dso_vgatest\[4\]
rlabel metal2 450570 211276 450570 211276 0 dso_vgatest\[5\]
rlabel metal2 450662 211344 450662 211344 0 dso_vgatest\[6\]
rlabel metal2 445172 104924 445172 104924 0 dso_vgatest\[7\]
rlabel metal2 450954 104924 450954 104924 0 dso_vgatest\[8\]
rlabel metal2 504942 304412 504942 304412 0 dso_vgatest\[9\]
rlabel metal2 580198 6715 580198 6715 0 io_in[0]
rlabel metal3 581218 458116 581218 458116 0 io_in[10]
rlabel metal3 582138 511292 582138 511292 0 io_in[11]
rlabel metal1 578588 563074 578588 563074 0 io_in[12]
rlabel metal2 580198 617185 580198 617185 0 io_in[13]
rlabel metal3 582000 670684 582000 670684 0 io_in[14]
rlabel metal3 559567 699788 559567 699788 0 io_in[15]
rlabel metal2 444314 510272 444314 510272 0 io_in[16]
rlabel metal2 429870 702178 429870 702178 0 io_in[17]
rlabel metal2 365010 702144 365010 702144 0 io_in[18]
rlabel metal2 449190 510952 449190 510952 0 io_in[19]
rlabel metal3 581218 46308 581218 46308 0 io_in[1]
rlabel metal2 235198 702093 235198 702093 0 io_in[20]
rlabel metal4 444268 510748 444268 510748 0 io_in[21]
rlabel metal2 445234 510714 445234 510714 0 io_in[22]
rlabel metal2 40526 701940 40526 701940 0 io_in[23]
rlabel metal3 1786 684284 1786 684284 0 io_in[24]
rlabel metal2 3772 678436 3772 678436 0 io_in[25]
rlabel metal3 1786 579972 1786 579972 0 io_in[26]
rlabel metal3 2154 527884 2154 527884 0 io_in[27]
rlabel metal2 3542 679116 3542 679116 0 io_in[28]
rlabel metal3 2016 423572 2016 423572 0 io_in[29]
rlabel metal2 580198 86547 580198 86547 0 io_in[2]
rlabel metal1 4600 214778 4600 214778 0 io_in[30]
rlabel metal1 4416 253946 4416 253946 0 io_in[31]
rlabel metal3 1924 267172 1924 267172 0 io_in[32]
rlabel metal3 2108 214948 2108 214948 0 io_in[33]
rlabel metal3 1832 162860 1832 162860 0 io_in[34]
rlabel metal3 1947 110636 1947 110636 0 io_in[35]
rlabel metal3 1740 71604 1740 71604 0 io_in[36]
rlabel metal3 1924 32436 1924 32436 0 io_in[37]
rlabel metal2 580198 126463 580198 126463 0 io_in[3]
rlabel metal2 580198 166413 580198 166413 0 io_in[4]
rlabel metal2 579830 206329 579830 206329 0 io_in[5]
rlabel via2 580198 245565 580198 245565 0 io_in[6]
rlabel metal2 461610 308074 461610 308074 0 io_in[7]
rlabel metal3 581862 351900 581862 351900 0 io_in[8]
rlabel metal3 582230 404940 582230 404940 0 io_in[9]
rlabel metal2 563730 171428 563730 171428 0 io_oeb[0]
rlabel metal2 580198 484517 580198 484517 0 io_oeb[10]
rlabel metal3 582092 537812 582092 537812 0 io_oeb[11]
rlabel metal2 580198 590835 580198 590835 0 io_oeb[12]
rlabel metal2 579646 643569 579646 643569 0 io_oeb[13]
rlabel metal3 581908 697204 581908 697204 0 io_oeb[14]
rlabel metal3 526769 699788 526769 699788 0 io_oeb[15]
rlabel metal2 450662 494530 450662 494530 0 io_oeb[16]
rlabel metal2 449098 328542 449098 328542 0 io_oeb[17]
rlabel metal2 332534 702110 332534 702110 0 io_oeb[18]
rlabel metal2 446890 501500 446890 501500 0 io_oeb[19]
rlabel metal2 544410 192134 544410 192134 0 io_oeb[1]
rlabel metal4 450708 501976 450708 501976 0 io_oeb[20]
rlabel metal2 137862 701957 137862 701957 0 io_oeb[21]
rlabel metal2 446982 326740 446982 326740 0 io_oeb[22]
rlabel metal4 446476 501636 446476 501636 0 io_oeb[23]
rlabel metal3 1740 658172 1740 658172 0 io_oeb[24]
rlabel metal3 1855 606084 1855 606084 0 io_oeb[25]
rlabel metal3 2200 553860 2200 553860 0 io_oeb[26]
rlabel metal3 2062 501772 2062 501772 0 io_oeb[27]
rlabel metal3 1878 449548 1878 449548 0 io_oeb[28]
rlabel metal1 5566 60690 5566 60690 0 io_oeb[29]
rlabel metal2 579830 112965 579830 112965 0 io_oeb[2]
rlabel metal1 4232 292774 4232 292774 0 io_oeb[30]
rlabel metal3 1878 293148 1878 293148 0 io_oeb[31]
rlabel metal3 2062 241060 2062 241060 0 io_oeb[32]
rlabel metal1 4094 45560 4094 45560 0 io_oeb[33]
rlabel metal3 1855 136748 1855 136748 0 io_oeb[34]
rlabel metal3 1740 84660 1740 84660 0 io_oeb[35]
rlabel metal3 1924 45492 1924 45492 0 io_oeb[36]
rlabel metal3 1878 6460 1878 6460 0 io_oeb[37]
rlabel metal2 580198 152915 580198 152915 0 io_oeb[3]
rlabel metal2 580198 192831 580198 192831 0 io_oeb[4]
rlabel metal2 580014 232781 580014 232781 0 io_oeb[5]
rlabel metal2 580198 272697 580198 272697 0 io_oeb[6]
rlabel metal2 509174 321164 509174 321164 0 io_oeb[7]
rlabel metal2 579830 378301 579830 378301 0 io_oeb[8]
rlabel metal2 580198 431103 580198 431103 0 io_oeb[9]
rlabel metal2 580014 20213 580014 20213 0 io_out[0]
rlabel metal2 467406 321582 467406 321582 0 io_out[10]
rlabel via2 580198 524467 580198 524467 0 io_out[11]
rlabel metal3 582046 577660 582046 577660 0 io_out[12]
rlabel metal2 468234 321684 468234 321684 0 io_out[13]
rlabel metal2 468510 320868 468510 320868 0 io_out[14]
rlabel metal2 468786 320936 468786 320936 0 io_out[15]
rlabel metal2 445694 510646 445694 510646 0 io_out[16]
rlabel metal2 469154 319583 469154 319583 0 io_out[17]
rlabel metal2 347806 693879 347806 693879 0 io_out[18]
rlabel metal2 446430 510578 446430 510578 0 io_out[19]
rlabel metal2 580198 60163 580198 60163 0 io_out[1]
rlabel metal2 218454 703596 218454 703596 0 io_out[20]
rlabel metal2 154146 702008 154146 702008 0 io_out[21]
rlabel metal2 88366 693811 88366 693811 0 io_out[22]
rlabel metal2 23828 703596 23828 703596 0 io_out[23]
rlabel metal3 2039 671228 2039 671228 0 io_out[24]
rlabel metal3 1947 619140 1947 619140 0 io_out[25]
rlabel metal3 1832 566916 1832 566916 0 io_out[26]
rlabel metal2 3680 679252 3680 679252 0 io_out[27]
rlabel metal3 1924 462604 1924 462604 0 io_out[28]
rlabel metal3 2154 410516 2154 410516 0 io_out[29]
rlabel metal2 580198 100079 580198 100079 0 io_out[2]
rlabel metal2 405674 154666 405674 154666 0 io_out[30]
rlabel metal3 2016 306204 2016 306204 0 io_out[31]
rlabel metal3 1970 254116 1970 254116 0 io_out[32]
rlabel metal3 2154 201892 2154 201892 0 io_out[33]
rlabel metal3 1786 149804 1786 149804 0 io_out[34]
rlabel metal3 2016 97580 2016 97580 0 io_out[35]
rlabel metal3 1878 58548 1878 58548 0 io_out[36]
rlabel metal3 1878 19380 1878 19380 0 io_out[37]
rlabel via2 580198 139349 580198 139349 0 io_out[3]
rlabel metal2 580198 179265 580198 179265 0 io_out[4]
rlabel metal2 580198 219215 580198 219215 0 io_out[5]
rlabel metal2 466302 296626 466302 296626 0 io_out[6]
rlabel metal2 580198 312647 580198 312647 0 io_out[7]
rlabel metal2 580198 364735 580198 364735 0 io_out[8]
rlabel metal2 467130 321072 467130 321072 0 io_out[9]
rlabel metal3 449788 158353 449788 158353 0 oeb_6502
rlabel via2 539373 137700 539373 137700 0 oeb_as1802
rlabel metal2 462477 385900 462477 385900 0 oeb_as2650
rlabel metal2 447166 384421 447166 384421 0 oeb_as512512512
rlabel metal2 502865 385900 502865 385900 0 oeb_as5401
rlabel via2 450501 358836 450501 358836 0 oeb_mc14500
rlabel metal2 448010 159868 448010 159868 0 rst_6502
rlabel metal2 427478 446036 427478 446036 0 rst_LCD
rlabel metal3 449980 345100 449980 345100 0 rst_as1802
rlabel metal3 450041 346188 450041 346188 0 rst_as2650
rlabel metal2 447166 347429 447166 347429 0 rst_as512512512
rlabel metal3 450087 346868 450087 346868 0 rst_as5401
rlabel via2 450363 348228 450363 348228 0 rst_counter
rlabel via2 450179 348908 450179 348908 0 rst_diceroll
rlabel metal3 448968 349180 448968 349180 0 rst_mc14500
rlabel metal3 449888 349860 449888 349860 0 rst_posit
rlabel via2 447166 350557 447166 350557 0 rst_tbb1143
rlabel metal3 449290 351220 449290 351220 0 rst_tune
rlabel via2 447166 351917 447166 351917 0 rst_vgatest
rlabel metal2 444912 160011 444912 160011 0 wb_clk_i
rlabel metal2 1702 1843 1702 1843 0 wb_rst_i
rlabel metal2 2898 1214 2898 1214 0 wbs_ack_o
rlabel metal2 384698 175389 384698 175389 0 wbs_adr_i[0]
rlabel metal2 47649 340 47649 340 0 wbs_adr_i[10]
rlabel metal2 51237 340 51237 340 0 wbs_adr_i[11]
rlabel metal1 217902 44982 217902 44982 0 wbs_adr_i[12]
rlabel metal2 58236 16560 58236 16560 0 wbs_adr_i[13]
rlabel metal2 61863 340 61863 340 0 wbs_adr_i[14]
rlabel metal2 65313 340 65313 340 0 wbs_adr_i[15]
rlabel metal1 224158 45254 224158 45254 0 wbs_adr_i[16]
rlabel metal1 225400 45322 225400 45322 0 wbs_adr_i[17]
rlabel metal2 76077 340 76077 340 0 wbs_adr_i[18]
rlabel metal2 79481 340 79481 340 0 wbs_adr_i[19]
rlabel metal2 12137 340 12137 340 0 wbs_adr_i[1]
rlabel metal2 83076 16560 83076 16560 0 wbs_adr_i[20]
rlabel metal2 86703 340 86703 340 0 wbs_adr_i[21]
rlabel metal2 90153 340 90153 340 0 wbs_adr_i[22]
rlabel metal2 93978 3627 93978 3627 0 wbs_adr_i[23]
rlabel metal2 97060 16560 97060 16560 0 wbs_adr_i[24]
rlabel metal2 100917 340 100917 340 0 wbs_adr_i[25]
rlabel metal2 373474 171496 373474 171496 0 wbs_adr_i[26]
rlabel metal2 373290 172754 373290 172754 0 wbs_adr_i[27]
rlabel metal2 370898 171530 370898 171530 0 wbs_adr_i[28]
rlabel metal2 114993 340 114993 340 0 wbs_adr_i[29]
rlabel metal2 17066 2183 17066 2183 0 wbs_adr_i[2]
rlabel metal2 118818 3627 118818 3627 0 wbs_adr_i[30]
rlabel metal2 121900 16560 121900 16560 0 wbs_adr_i[31]
rlabel metal2 21298 16560 21298 16560 0 wbs_adr_i[3]
rlabel metal2 368046 169745 368046 169745 0 wbs_adr_i[4]
rlabel metal2 367862 150076 367862 150076 0 wbs_adr_i[5]
rlabel metal2 368138 169796 368138 169796 0 wbs_adr_i[6]
rlabel metal2 37214 1996 37214 1996 0 wbs_adr_i[7]
rlabel metal2 40473 340 40473 340 0 wbs_adr_i[8]
rlabel metal2 44298 3627 44298 3627 0 wbs_adr_i[9]
rlabel metal2 3857 340 3857 340 0 wbs_cyc_i
rlabel metal2 365194 150909 365194 150909 0 wbs_dat_i[0]
rlabel metal2 365102 150824 365102 150824 0 wbs_dat_i[10]
rlabel metal2 52578 2030 52578 2030 0 wbs_dat_i[11]
rlabel metal2 56074 2166 56074 2166 0 wbs_dat_i[12]
rlabel metal2 59517 340 59517 340 0 wbs_dat_i[13]
rlabel metal2 62698 16560 62698 16560 0 wbs_dat_i[14]
rlabel metal1 214268 39814 214268 39814 0 wbs_dat_i[15]
rlabel metal2 70097 340 70097 340 0 wbs_dat_i[16]
rlabel metal2 73593 340 73593 340 0 wbs_dat_i[17]
rlabel metal2 77418 3627 77418 3627 0 wbs_dat_i[18]
rlabel metal2 80500 16560 80500 16560 0 wbs_dat_i[19]
rlabel metal2 370530 154632 370530 154632 0 wbs_dat_i[1]
rlabel metal2 84357 340 84357 340 0 wbs_dat_i[20]
rlabel metal2 366482 165886 366482 165886 0 wbs_dat_i[21]
rlabel metal2 368230 165614 368230 165614 0 wbs_dat_i[22]
rlabel metal2 94937 340 94937 340 0 wbs_dat_i[23]
rlabel metal2 98433 340 98433 340 0 wbs_dat_i[24]
rlabel metal2 102258 3627 102258 3627 0 wbs_dat_i[25]
rlabel metal2 369150 166090 369150 166090 0 wbs_dat_i[26]
rlabel metal2 369242 166192 369242 166192 0 wbs_dat_i[27]
rlabel metal2 369334 166056 369334 166056 0 wbs_dat_i[28]
rlabel metal2 116196 16560 116196 16560 0 wbs_dat_i[29]
rlabel metal2 18117 340 18117 340 0 wbs_dat_i[2]
rlabel metal2 119370 16560 119370 16560 0 wbs_dat_i[30]
rlabel metal2 371910 211480 371910 211480 0 wbs_dat_i[31]
rlabel metal2 22809 340 22809 340 0 wbs_dat_i[3]
rlabel metal2 519662 312358 519662 312358 0 wbs_dat_i[4]
rlabel metal2 519478 313140 519478 313140 0 wbs_dat_i[5]
rlabel metal2 520950 314432 520950 314432 0 wbs_dat_i[6]
rlabel metal2 38410 1894 38410 1894 0 wbs_dat_i[7]
rlabel metal2 41906 1962 41906 1962 0 wbs_dat_i[8]
rlabel metal2 45257 340 45257 340 0 wbs_dat_i[9]
rlabel metal2 507702 306527 507702 306527 0 wbs_dat_o[0]
rlabel metal2 520766 318070 520766 318070 0 wbs_dat_o[10]
rlabel metal2 520674 318784 520674 318784 0 wbs_dat_o[11]
rlabel metal2 57270 2132 57270 2132 0 wbs_dat_o[12]
rlabel metal2 60858 17262 60858 17262 0 wbs_dat_o[13]
rlabel metal2 63940 16560 63940 16560 0 wbs_dat_o[14]
rlabel metal2 67797 340 67797 340 0 wbs_dat_o[15]
rlabel metal1 449788 289782 449788 289782 0 wbs_dat_o[16]
rlabel metal2 74796 16560 74796 16560 0 wbs_dat_o[17]
rlabel metal2 78377 340 78377 340 0 wbs_dat_o[18]
rlabel metal2 82110 2200 82110 2200 0 wbs_dat_o[19]
rlabel metal2 385986 160038 385986 160038 0 wbs_dat_o[1]
rlabel metal2 386262 161670 386262 161670 0 wbs_dat_o[20]
rlabel metal2 89194 2234 89194 2234 0 wbs_dat_o[21]
rlabel metal2 92637 340 92637 340 0 wbs_dat_o[22]
rlabel metal2 96278 1860 96278 1860 0 wbs_dat_o[23]
rlabel metal2 99636 16560 99636 16560 0 wbs_dat_o[24]
rlabel metal2 102810 16560 102810 16560 0 wbs_dat_o[25]
rlabel metal2 106950 1758 106950 1758 0 wbs_dat_o[26]
rlabel metal2 110538 1690 110538 1690 0 wbs_dat_o[27]
rlabel metal2 113620 16560 113620 16560 0 wbs_dat_o[28]
rlabel metal2 117477 340 117477 340 0 wbs_dat_o[29]
rlabel metal2 19412 16560 19412 16560 0 wbs_dat_o[2]
rlabel metal2 120881 340 120881 340 0 wbs_dat_o[30]
rlabel metal2 366390 207978 366390 207978 0 wbs_dat_o[31]
rlabel metal2 24242 1911 24242 1911 0 wbs_dat_o[3]
rlabel metal2 386078 160208 386078 160208 0 wbs_dat_o[4]
rlabel metal2 384974 158814 384974 158814 0 wbs_dat_o[5]
rlabel metal2 35972 16560 35972 16560 0 wbs_dat_o[6]
rlabel metal2 39369 340 39369 340 0 wbs_dat_o[7]
rlabel metal2 43102 2064 43102 2064 0 wbs_dat_o[8]
rlabel metal2 521686 314364 521686 314364 0 wbs_dat_o[9]
rlabel metal2 5290 2115 5290 2115 0 wbs_stb_i
rlabel metal2 6486 1792 6486 1792 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
