// This is the unpowered netlist.
module wrapped_as2650 (clk,
    io_oeb,
    rst,
    io_in,
    io_out);
 input clk;
 output io_oeb;
 input rst;
 input [8:0] io_in;
 output [26:0] io_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire \as2650.addr_buff[0] ;
 wire \as2650.addr_buff[1] ;
 wire \as2650.addr_buff[2] ;
 wire \as2650.addr_buff[3] ;
 wire \as2650.addr_buff[4] ;
 wire \as2650.addr_buff[5] ;
 wire \as2650.addr_buff[6] ;
 wire \as2650.addr_buff[7] ;
 wire \as2650.carry ;
 wire \as2650.cycle[0] ;
 wire \as2650.cycle[1] ;
 wire \as2650.cycle[2] ;
 wire \as2650.cycle[3] ;
 wire \as2650.cycle[4] ;
 wire \as2650.cycle[5] ;
 wire \as2650.cycle[6] ;
 wire \as2650.cycle[7] ;
 wire \as2650.halted ;
 wire \as2650.holding_reg[0] ;
 wire \as2650.holding_reg[1] ;
 wire \as2650.holding_reg[2] ;
 wire \as2650.holding_reg[3] ;
 wire \as2650.holding_reg[4] ;
 wire \as2650.holding_reg[5] ;
 wire \as2650.holding_reg[6] ;
 wire \as2650.holding_reg[7] ;
 wire \as2650.idx_ctrl[0] ;
 wire \as2650.idx_ctrl[1] ;
 wire \as2650.ins_reg[0] ;
 wire \as2650.ins_reg[1] ;
 wire \as2650.ins_reg[2] ;
 wire \as2650.ins_reg[3] ;
 wire \as2650.ins_reg[4] ;
 wire \as2650.ins_reg[5] ;
 wire \as2650.ins_reg[6] ;
 wire \as2650.ins_reg[7] ;
 wire \as2650.overflow ;
 wire \as2650.pc[0] ;
 wire \as2650.pc[10] ;
 wire \as2650.pc[11] ;
 wire \as2650.pc[12] ;
 wire \as2650.pc[13] ;
 wire \as2650.pc[14] ;
 wire \as2650.pc[1] ;
 wire \as2650.pc[2] ;
 wire \as2650.pc[3] ;
 wire \as2650.pc[4] ;
 wire \as2650.pc[5] ;
 wire \as2650.pc[6] ;
 wire \as2650.pc[7] ;
 wire \as2650.pc[8] ;
 wire \as2650.pc[9] ;
 wire \as2650.psl[1] ;
 wire \as2650.psl[3] ;
 wire \as2650.psl[4] ;
 wire \as2650.psl[5] ;
 wire \as2650.psl[6] ;
 wire \as2650.psl[7] ;
 wire \as2650.psu[0] ;
 wire \as2650.psu[1] ;
 wire \as2650.psu[2] ;
 wire \as2650.psu[3] ;
 wire \as2650.psu[4] ;
 wire \as2650.psu[5] ;
 wire \as2650.psu[7] ;
 wire \as2650.r0[0] ;
 wire \as2650.r0[1] ;
 wire \as2650.r0[2] ;
 wire \as2650.r0[3] ;
 wire \as2650.r0[4] ;
 wire \as2650.r0[5] ;
 wire \as2650.r0[6] ;
 wire \as2650.r0[7] ;
 wire \as2650.r123[0][0] ;
 wire \as2650.r123[0][1] ;
 wire \as2650.r123[0][2] ;
 wire \as2650.r123[0][3] ;
 wire \as2650.r123[0][4] ;
 wire \as2650.r123[0][5] ;
 wire \as2650.r123[0][6] ;
 wire \as2650.r123[0][7] ;
 wire \as2650.r123[1][0] ;
 wire \as2650.r123[1][1] ;
 wire \as2650.r123[1][2] ;
 wire \as2650.r123[1][3] ;
 wire \as2650.r123[1][4] ;
 wire \as2650.r123[1][5] ;
 wire \as2650.r123[1][6] ;
 wire \as2650.r123[1][7] ;
 wire \as2650.r123[2][0] ;
 wire \as2650.r123[2][1] ;
 wire \as2650.r123[2][2] ;
 wire \as2650.r123[2][3] ;
 wire \as2650.r123[2][4] ;
 wire \as2650.r123[2][5] ;
 wire \as2650.r123[2][6] ;
 wire \as2650.r123[2][7] ;
 wire \as2650.r123[3][0] ;
 wire \as2650.r123[3][1] ;
 wire \as2650.r123[3][2] ;
 wire \as2650.r123[3][3] ;
 wire \as2650.r123[3][4] ;
 wire \as2650.r123[3][5] ;
 wire \as2650.r123[3][6] ;
 wire \as2650.r123[3][7] ;
 wire \as2650.r123_2[0][0] ;
 wire \as2650.r123_2[0][1] ;
 wire \as2650.r123_2[0][2] ;
 wire \as2650.r123_2[0][3] ;
 wire \as2650.r123_2[0][4] ;
 wire \as2650.r123_2[0][5] ;
 wire \as2650.r123_2[0][6] ;
 wire \as2650.r123_2[0][7] ;
 wire \as2650.r123_2[1][0] ;
 wire \as2650.r123_2[1][1] ;
 wire \as2650.r123_2[1][2] ;
 wire \as2650.r123_2[1][3] ;
 wire \as2650.r123_2[1][4] ;
 wire \as2650.r123_2[1][5] ;
 wire \as2650.r123_2[1][6] ;
 wire \as2650.r123_2[1][7] ;
 wire \as2650.r123_2[2][0] ;
 wire \as2650.r123_2[2][1] ;
 wire \as2650.r123_2[2][2] ;
 wire \as2650.r123_2[2][3] ;
 wire \as2650.r123_2[2][4] ;
 wire \as2650.r123_2[2][5] ;
 wire \as2650.r123_2[2][6] ;
 wire \as2650.r123_2[2][7] ;
 wire \as2650.r123_2[3][0] ;
 wire \as2650.r123_2[3][1] ;
 wire \as2650.r123_2[3][2] ;
 wire \as2650.r123_2[3][3] ;
 wire \as2650.r123_2[3][4] ;
 wire \as2650.r123_2[3][5] ;
 wire \as2650.r123_2[3][6] ;
 wire \as2650.r123_2[3][7] ;
 wire \as2650.stack[0][0] ;
 wire \as2650.stack[0][10] ;
 wire \as2650.stack[0][11] ;
 wire \as2650.stack[0][12] ;
 wire \as2650.stack[0][13] ;
 wire \as2650.stack[0][14] ;
 wire \as2650.stack[0][1] ;
 wire \as2650.stack[0][2] ;
 wire \as2650.stack[0][3] ;
 wire \as2650.stack[0][4] ;
 wire \as2650.stack[0][5] ;
 wire \as2650.stack[0][6] ;
 wire \as2650.stack[0][7] ;
 wire \as2650.stack[0][8] ;
 wire \as2650.stack[0][9] ;
 wire \as2650.stack[1][0] ;
 wire \as2650.stack[1][10] ;
 wire \as2650.stack[1][11] ;
 wire \as2650.stack[1][12] ;
 wire \as2650.stack[1][13] ;
 wire \as2650.stack[1][14] ;
 wire \as2650.stack[1][1] ;
 wire \as2650.stack[1][2] ;
 wire \as2650.stack[1][3] ;
 wire \as2650.stack[1][4] ;
 wire \as2650.stack[1][5] ;
 wire \as2650.stack[1][6] ;
 wire \as2650.stack[1][7] ;
 wire \as2650.stack[1][8] ;
 wire \as2650.stack[1][9] ;
 wire \as2650.stack[2][0] ;
 wire \as2650.stack[2][10] ;
 wire \as2650.stack[2][11] ;
 wire \as2650.stack[2][12] ;
 wire \as2650.stack[2][13] ;
 wire \as2650.stack[2][14] ;
 wire \as2650.stack[2][1] ;
 wire \as2650.stack[2][2] ;
 wire \as2650.stack[2][3] ;
 wire \as2650.stack[2][4] ;
 wire \as2650.stack[2][5] ;
 wire \as2650.stack[2][6] ;
 wire \as2650.stack[2][7] ;
 wire \as2650.stack[2][8] ;
 wire \as2650.stack[2][9] ;
 wire \as2650.stack[3][0] ;
 wire \as2650.stack[3][10] ;
 wire \as2650.stack[3][11] ;
 wire \as2650.stack[3][12] ;
 wire \as2650.stack[3][13] ;
 wire \as2650.stack[3][14] ;
 wire \as2650.stack[3][1] ;
 wire \as2650.stack[3][2] ;
 wire \as2650.stack[3][3] ;
 wire \as2650.stack[3][4] ;
 wire \as2650.stack[3][5] ;
 wire \as2650.stack[3][6] ;
 wire \as2650.stack[3][7] ;
 wire \as2650.stack[3][8] ;
 wire \as2650.stack[3][9] ;
 wire \as2650.stack[4][0] ;
 wire \as2650.stack[4][10] ;
 wire \as2650.stack[4][11] ;
 wire \as2650.stack[4][12] ;
 wire \as2650.stack[4][13] ;
 wire \as2650.stack[4][14] ;
 wire \as2650.stack[4][1] ;
 wire \as2650.stack[4][2] ;
 wire \as2650.stack[4][3] ;
 wire \as2650.stack[4][4] ;
 wire \as2650.stack[4][5] ;
 wire \as2650.stack[4][6] ;
 wire \as2650.stack[4][7] ;
 wire \as2650.stack[4][8] ;
 wire \as2650.stack[4][9] ;
 wire \as2650.stack[5][0] ;
 wire \as2650.stack[5][10] ;
 wire \as2650.stack[5][11] ;
 wire \as2650.stack[5][12] ;
 wire \as2650.stack[5][13] ;
 wire \as2650.stack[5][14] ;
 wire \as2650.stack[5][1] ;
 wire \as2650.stack[5][2] ;
 wire \as2650.stack[5][3] ;
 wire \as2650.stack[5][4] ;
 wire \as2650.stack[5][5] ;
 wire \as2650.stack[5][6] ;
 wire \as2650.stack[5][7] ;
 wire \as2650.stack[5][8] ;
 wire \as2650.stack[5][9] ;
 wire \as2650.stack[6][0] ;
 wire \as2650.stack[6][10] ;
 wire \as2650.stack[6][11] ;
 wire \as2650.stack[6][12] ;
 wire \as2650.stack[6][13] ;
 wire \as2650.stack[6][14] ;
 wire \as2650.stack[6][1] ;
 wire \as2650.stack[6][2] ;
 wire \as2650.stack[6][3] ;
 wire \as2650.stack[6][4] ;
 wire \as2650.stack[6][5] ;
 wire \as2650.stack[6][6] ;
 wire \as2650.stack[6][7] ;
 wire \as2650.stack[6][8] ;
 wire \as2650.stack[6][9] ;
 wire \as2650.stack[7][0] ;
 wire \as2650.stack[7][10] ;
 wire \as2650.stack[7][11] ;
 wire \as2650.stack[7][12] ;
 wire \as2650.stack[7][13] ;
 wire \as2650.stack[7][14] ;
 wire \as2650.stack[7][1] ;
 wire \as2650.stack[7][2] ;
 wire \as2650.stack[7][3] ;
 wire \as2650.stack[7][4] ;
 wire \as2650.stack[7][5] ;
 wire \as2650.stack[7][6] ;
 wire \as2650.stack[7][7] ;
 wire \as2650.stack[7][8] ;
 wire \as2650.stack[7][9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 sky130_fd_sc_hd__inv_2 _2933_ (.A(net30),
    .Y(_2524_));
 sky130_fd_sc_hd__inv_4 _2934_ (.A(net213),
    .Y(_2525_));
 sky130_fd_sc_hd__clkinv_2 _2935_ (.A(\as2650.carry ),
    .Y(_2526_));
 sky130_fd_sc_hd__inv_2 _2936_ (.A(net215),
    .Y(_2527_));
 sky130_fd_sc_hd__inv_2 _2937_ (.A(net217),
    .Y(_2528_));
 sky130_fd_sc_hd__inv_2 _2938_ (.A(net220),
    .Y(_2529_));
 sky130_fd_sc_hd__inv_2 _2939_ (.A(net235),
    .Y(_2530_));
 sky130_fd_sc_hd__inv_2 _2940_ (.A(net266),
    .Y(_2531_));
 sky130_fd_sc_hd__inv_2 _2941_ (.A(net268),
    .Y(_2532_));
 sky130_fd_sc_hd__inv_2 _2942_ (.A(net276),
    .Y(_2533_));
 sky130_fd_sc_hd__clkinv_2 _2943_ (.A(net285),
    .Y(_2534_));
 sky130_fd_sc_hd__inv_6 _2944_ (.A(\as2650.halted ),
    .Y(_2535_));
 sky130_fd_sc_hd__clkinv_4 _2945_ (.A(\as2650.cycle[7] ),
    .Y(_2536_));
 sky130_fd_sc_hd__inv_6 _2946_ (.A(\as2650.cycle[1] ),
    .Y(_2537_));
 sky130_fd_sc_hd__clkinv_2 _2947_ (.A(net25),
    .Y(net11));
 sky130_fd_sc_hd__inv_2 _2948_ (.A(net22),
    .Y(_2538_));
 sky130_fd_sc_hd__inv_2 _2949_ (.A(net21),
    .Y(_2539_));
 sky130_fd_sc_hd__inv_2 _2950_ (.A(net16),
    .Y(_2540_));
 sky130_fd_sc_hd__inv_2 _2951_ (.A(net14),
    .Y(_2541_));
 sky130_fd_sc_hd__inv_2 _2952_ (.A(net37),
    .Y(_2542_));
 sky130_fd_sc_hd__inv_2 _2953_ (.A(net304),
    .Y(_2543_));
 sky130_fd_sc_hd__inv_2 _2954_ (.A(net302),
    .Y(_2544_));
 sky130_fd_sc_hd__inv_2 _2955_ (.A(net229),
    .Y(_2545_));
 sky130_fd_sc_hd__inv_2 _2956_ (.A(net223),
    .Y(_2546_));
 sky130_fd_sc_hd__clkinv_2 _2957_ (.A(net10),
    .Y(_2547_));
 sky130_fd_sc_hd__inv_2 _2958_ (.A(net325),
    .Y(_2548_));
 sky130_fd_sc_hd__inv_2 _2959_ (.A(net350),
    .Y(_2549_));
 sky130_fd_sc_hd__inv_4 _2960_ (.A(net345),
    .Y(_2550_));
 sky130_fd_sc_hd__inv_2 _2961_ (.A(net341),
    .Y(_2551_));
 sky130_fd_sc_hd__clkinv_4 _2962_ (.A(net339),
    .Y(_2552_));
 sky130_fd_sc_hd__clkinv_4 _2963_ (.A(net335),
    .Y(_2553_));
 sky130_fd_sc_hd__clkinv_4 _2964_ (.A(net334),
    .Y(_2554_));
 sky130_fd_sc_hd__inv_2 _2965_ (.A(\as2650.holding_reg[5] ),
    .Y(_2555_));
 sky130_fd_sc_hd__inv_4 _2966_ (.A(net331),
    .Y(_2556_));
 sky130_fd_sc_hd__clkinv_2 _2967_ (.A(net296),
    .Y(_2557_));
 sky130_fd_sc_hd__nand2_1 _2968_ (.A(_2527_),
    .B(net217),
    .Y(_2558_));
 sky130_fd_sc_hd__or2_4 _2969_ (.A(_2529_),
    .B(net168),
    .X(_2559_));
 sky130_fd_sc_hd__nor2_8 _2970_ (.A(net293),
    .B(net347),
    .Y(_2560_));
 sky130_fd_sc_hd__or2_4 _2971_ (.A(net293),
    .B(net347),
    .X(_2561_));
 sky130_fd_sc_hd__nor4_2 _2972_ (.A(\as2650.cycle[5] ),
    .B(\as2650.cycle[4] ),
    .C(net288),
    .D(net289),
    .Y(_2562_));
 sky130_fd_sc_hd__or4_4 _2973_ (.A(\as2650.cycle[7] ),
    .B(\as2650.cycle[6] ),
    .C(\as2650.cycle[5] ),
    .D(\as2650.cycle[4] ),
    .X(_2563_));
 sky130_fd_sc_hd__nor3_4 _2974_ (.A(net288),
    .B(net289),
    .C(_2563_),
    .Y(_2564_));
 sky130_fd_sc_hd__or3_4 _2975_ (.A(net288),
    .B(net289),
    .C(_2563_),
    .X(_2565_));
 sky130_fd_sc_hd__nor2_4 _2976_ (.A(_2537_),
    .B(net290),
    .Y(_2566_));
 sky130_fd_sc_hd__nor2_2 _2977_ (.A(_2537_),
    .B(net164),
    .Y(_2567_));
 sky130_fd_sc_hd__nand2_4 _2978_ (.A(\as2650.cycle[1] ),
    .B(net165),
    .Y(_2568_));
 sky130_fd_sc_hd__nor2_1 _2979_ (.A(net291),
    .B(net148),
    .Y(_2569_));
 sky130_fd_sc_hd__nand2_4 _2980_ (.A(net165),
    .B(net163),
    .Y(_2570_));
 sky130_fd_sc_hd__nor2_8 _2981_ (.A(net299),
    .B(net298),
    .Y(_2571_));
 sky130_fd_sc_hd__nand2_8 _2982_ (.A(net226),
    .B(_2571_),
    .Y(_2572_));
 sky130_fd_sc_hd__nor2_1 _2983_ (.A(net300),
    .B(_2572_),
    .Y(_2573_));
 sky130_fd_sc_hd__or2_1 _2984_ (.A(net300),
    .B(_2572_),
    .X(_2574_));
 sky130_fd_sc_hd__nor2_1 _2985_ (.A(net303),
    .B(net231),
    .Y(_2575_));
 sky130_fd_sc_hd__or2_4 _2986_ (.A(net303),
    .B(net231),
    .X(_2576_));
 sky130_fd_sc_hd__and2b_4 _2987_ (.A_N(net304),
    .B(net306),
    .X(_2577_));
 sky130_fd_sc_hd__nand2_1 _2988_ (.A(_2543_),
    .B(net308),
    .Y(_2578_));
 sky130_fd_sc_hd__and3_4 _2989_ (.A(_2573_),
    .B(net201),
    .C(_2577_),
    .X(_2579_));
 sky130_fd_sc_hd__and2_4 _2990_ (.A(net78),
    .B(_2579_),
    .X(_2580_));
 sky130_fd_sc_hd__nand2_2 _2991_ (.A(_2560_),
    .B(_2580_),
    .Y(_2581_));
 sky130_fd_sc_hd__or2_4 _2992_ (.A(_2559_),
    .B(net49),
    .X(_2582_));
 sky130_fd_sc_hd__and2_4 _2993_ (.A(net304),
    .B(net306),
    .X(_2583_));
 sky130_fd_sc_hd__nand2_8 _2994_ (.A(net305),
    .B(net306),
    .Y(_2584_));
 sky130_fd_sc_hd__and2b_4 _2995_ (.A_N(\as2650.ins_reg[6] ),
    .B(net297),
    .X(_2585_));
 sky130_fd_sc_hd__nand2b_4 _2996_ (.A_N(net299),
    .B(net298),
    .Y(_2586_));
 sky130_fd_sc_hd__nor2_4 _2997_ (.A(net206),
    .B(net202),
    .Y(_2587_));
 sky130_fd_sc_hd__nand2_2 _2998_ (.A(net229),
    .B(net225),
    .Y(_2588_));
 sky130_fd_sc_hd__and3_1 _2999_ (.A(net196),
    .B(net195),
    .C(net162),
    .X(_2589_));
 sky130_fd_sc_hd__or3_4 _3000_ (.A(_2584_),
    .B(_2586_),
    .C(net194),
    .X(_2590_));
 sky130_fd_sc_hd__nor2_2 _3001_ (.A(net208),
    .B(_2590_),
    .Y(_2591_));
 sky130_fd_sc_hd__or2_2 _3002_ (.A(net208),
    .B(_2590_),
    .X(_2592_));
 sky130_fd_sc_hd__or2_4 _3003_ (.A(\as2650.cycle[1] ),
    .B(net290),
    .X(_2593_));
 sky130_fd_sc_hd__nor3b_4 _3004_ (.A(_2563_),
    .B(\as2650.cycle[3] ),
    .C_N(net289),
    .Y(_2594_));
 sky130_fd_sc_hd__or3b_4 _3005_ (.A(_2593_),
    .B(net288),
    .C_N(\as2650.cycle[2] ),
    .X(_2595_));
 sky130_fd_sc_hd__nor2_4 _3006_ (.A(_2563_),
    .B(_2595_),
    .Y(_2596_));
 sky130_fd_sc_hd__or2_4 _3007_ (.A(_2563_),
    .B(_2595_),
    .X(_2597_));
 sky130_fd_sc_hd__and3_4 _3008_ (.A(net300),
    .B(net136),
    .C(net130),
    .X(_2598_));
 sky130_fd_sc_hd__nand2_8 _3009_ (.A(net299),
    .B(net297),
    .Y(_2599_));
 sky130_fd_sc_hd__nand2_4 _3010_ (.A(net224),
    .B(net301),
    .Y(_2600_));
 sky130_fd_sc_hd__nor2_4 _3011_ (.A(net302),
    .B(_2590_),
    .Y(_2601_));
 sky130_fd_sc_hd__or2_4 _3012_ (.A(net302),
    .B(_2590_),
    .X(_2602_));
 sky130_fd_sc_hd__nor2_8 _3013_ (.A(net206),
    .B(net120),
    .Y(_2603_));
 sky130_fd_sc_hd__or2_2 _3014_ (.A(net206),
    .B(net120),
    .X(_2604_));
 sky130_fd_sc_hd__or3b_2 _3015_ (.A(_2600_),
    .B(_2604_),
    .C_N(_2599_),
    .X(_2605_));
 sky130_fd_sc_hd__and4bb_4 _3016_ (.A_N(\as2650.cycle[2] ),
    .B_N(_2563_),
    .C(_2537_),
    .D(net288),
    .X(_2606_));
 sky130_fd_sc_hd__nand2_8 _3017_ (.A(net291),
    .B(_2606_),
    .Y(_2607_));
 sky130_fd_sc_hd__nand2_8 _3018_ (.A(\as2650.cycle[1] ),
    .B(net290),
    .Y(_2608_));
 sky130_fd_sc_hd__nor4_4 _3019_ (.A(\as2650.cycle[3] ),
    .B(net289),
    .C(_2563_),
    .D(_2608_),
    .Y(_2609_));
 sky130_fd_sc_hd__or4_4 _3020_ (.A(net288),
    .B(net289),
    .C(_2563_),
    .D(_2608_),
    .X(_2610_));
 sky130_fd_sc_hd__nor2_2 _3021_ (.A(net324),
    .B(_2610_),
    .Y(_2611_));
 sky130_fd_sc_hd__nor2_8 _3022_ (.A(net164),
    .B(_2608_),
    .Y(_2612_));
 sky130_fd_sc_hd__or2_2 _3023_ (.A(net164),
    .B(_2608_),
    .X(_2613_));
 sky130_fd_sc_hd__o2bb2a_1 _3024_ (.A1_N(net208),
    .A2_N(_2611_),
    .B1(_2591_),
    .B2(_2607_),
    .X(_2614_));
 sky130_fd_sc_hd__nor2_4 _3025_ (.A(net294),
    .B(net123),
    .Y(_2615_));
 sky130_fd_sc_hd__or2_4 _3026_ (.A(net294),
    .B(net122),
    .X(_2616_));
 sky130_fd_sc_hd__a21oi_2 _3027_ (.A1(_2614_),
    .A2(_2616_),
    .B1(_2605_),
    .Y(_2617_));
 sky130_fd_sc_hd__o21ai_4 _3028_ (.A1(_2598_),
    .A2(_2617_),
    .B1(_2560_),
    .Y(_2618_));
 sky130_fd_sc_hd__o21ai_4 _3029_ (.A1(_2559_),
    .A2(_2618_),
    .B1(_2582_),
    .Y(_2619_));
 sky130_fd_sc_hd__nor2_1 _3030_ (.A(net300),
    .B(_2592_),
    .Y(_2620_));
 sky130_fd_sc_hd__o31a_1 _3031_ (.A1(net294),
    .A2(net124),
    .A3(_2620_),
    .B1(_2614_),
    .X(_2621_));
 sky130_fd_sc_hd__nor2_1 _3032_ (.A(_2605_),
    .B(_2621_),
    .Y(_2622_));
 sky130_fd_sc_hd__o21ai_4 _3033_ (.A1(_2598_),
    .A2(_2622_),
    .B1(_2560_),
    .Y(_2623_));
 sky130_fd_sc_hd__mux2_1 _3034_ (.A0(\as2650.r123[0][0] ),
    .A1(\as2650.r123_2[0][0] ),
    .S(net213),
    .X(_2624_));
 sky130_fd_sc_hd__mux2_8 _3035_ (.A0(net192),
    .A1(\as2650.pc[8] ),
    .S(net48),
    .X(_2625_));
 sky130_fd_sc_hd__nor2_2 _3036_ (.A(net302),
    .B(_2610_),
    .Y(_2626_));
 sky130_fd_sc_hd__nand2_8 _3037_ (.A(net208),
    .B(net161),
    .Y(_2627_));
 sky130_fd_sc_hd__o21a_1 _3038_ (.A1(net324),
    .A2(_2627_),
    .B1(_2607_),
    .X(_2628_));
 sky130_fd_sc_hd__o22a_1 _3039_ (.A1(_2616_),
    .A2(_2620_),
    .B1(_2628_),
    .B2(net136),
    .X(_2629_));
 sky130_fd_sc_hd__nor2_1 _3040_ (.A(_2605_),
    .B(_2629_),
    .Y(_2630_));
 sky130_fd_sc_hd__o21ai_4 _3041_ (.A1(_2598_),
    .A2(_2630_),
    .B1(_2560_),
    .Y(_2631_));
 sky130_fd_sc_hd__mux2_1 _3042_ (.A0(\as2650.stack[6][8] ),
    .A1(_2625_),
    .S(_2619_),
    .X(_0000_));
 sky130_fd_sc_hd__mux2_8 _3043_ (.A0(\as2650.r123[0][1] ),
    .A1(\as2650.r123_2[0][1] ),
    .S(net214),
    .X(_2632_));
 sky130_fd_sc_hd__mux2_8 _3044_ (.A0(_2632_),
    .A1(\as2650.pc[9] ),
    .S(net48),
    .X(_2633_));
 sky130_fd_sc_hd__mux2_1 _3045_ (.A0(\as2650.stack[6][9] ),
    .A1(_2633_),
    .S(_2619_),
    .X(_0001_));
 sky130_fd_sc_hd__mux2_8 _3046_ (.A0(\as2650.r123[0][2] ),
    .A1(\as2650.r123_2[0][2] ),
    .S(net212),
    .X(_2634_));
 sky130_fd_sc_hd__mux2_4 _3047_ (.A0(_2634_),
    .A1(net266),
    .S(net48),
    .X(_2635_));
 sky130_fd_sc_hd__mux2_1 _3048_ (.A0(\as2650.stack[6][10] ),
    .A1(_2635_),
    .S(_2619_),
    .X(_0002_));
 sky130_fd_sc_hd__mux2_8 _3049_ (.A0(\as2650.r123[0][3] ),
    .A1(\as2650.r123_2[0][3] ),
    .S(net210),
    .X(_2636_));
 sky130_fd_sc_hd__mux2_8 _3050_ (.A0(_2636_),
    .A1(net265),
    .S(net48),
    .X(_2637_));
 sky130_fd_sc_hd__mux2_1 _3051_ (.A0(\as2650.stack[6][11] ),
    .A1(_2637_),
    .S(_2619_),
    .X(_0003_));
 sky130_fd_sc_hd__mux2_8 _3052_ (.A0(\as2650.r123[0][4] ),
    .A1(\as2650.r123_2[0][4] ),
    .S(net212),
    .X(_2638_));
 sky130_fd_sc_hd__mux2_8 _3053_ (.A0(_2638_),
    .A1(net264),
    .S(net48),
    .X(_2639_));
 sky130_fd_sc_hd__mux2_1 _3054_ (.A0(\as2650.stack[6][12] ),
    .A1(_2639_),
    .S(_2619_),
    .X(_0004_));
 sky130_fd_sc_hd__mux2_2 _3055_ (.A0(\as2650.r123[0][5] ),
    .A1(\as2650.r123_2[0][5] ),
    .S(net210),
    .X(_2640_));
 sky130_fd_sc_hd__mux2_8 _3056_ (.A0(net182),
    .A1(\as2650.pc[13] ),
    .S(net49),
    .X(_2641_));
 sky130_fd_sc_hd__mux2_1 _3057_ (.A0(\as2650.stack[6][13] ),
    .A1(_2641_),
    .S(_2619_),
    .X(_0005_));
 sky130_fd_sc_hd__mux2_2 _3058_ (.A0(\as2650.r123[0][6] ),
    .A1(\as2650.r123_2[0][6] ),
    .S(net210),
    .X(_2642_));
 sky130_fd_sc_hd__mux2_8 _3059_ (.A0(net180),
    .A1(\as2650.pc[14] ),
    .S(net49),
    .X(_2643_));
 sky130_fd_sc_hd__mux2_1 _3060_ (.A0(\as2650.stack[6][14] ),
    .A1(_2643_),
    .S(_2619_),
    .X(_0006_));
 sky130_fd_sc_hd__nor2_2 _3061_ (.A(net305),
    .B(net306),
    .Y(_2644_));
 sky130_fd_sc_hd__or2_4 _3062_ (.A(net304),
    .B(net308),
    .X(_2645_));
 sky130_fd_sc_hd__nor2_8 _3063_ (.A(net212),
    .B(net144),
    .Y(_2646_));
 sky130_fd_sc_hd__nand2_8 _3064_ (.A(_2560_),
    .B(_2646_),
    .Y(_2647_));
 sky130_fd_sc_hd__or2_4 _3065_ (.A(net177),
    .B(_2647_),
    .X(_2648_));
 sky130_fd_sc_hd__nand2_4 _3066_ (.A(net224),
    .B(net299),
    .Y(_2649_));
 sky130_fd_sc_hd__nor2_4 _3067_ (.A(net204),
    .B(_2599_),
    .Y(_2650_));
 sky130_fd_sc_hd__nor2_2 _3068_ (.A(net300),
    .B(_2599_),
    .Y(_2651_));
 sky130_fd_sc_hd__or2_4 _3069_ (.A(net300),
    .B(_2599_),
    .X(_2652_));
 sky130_fd_sc_hd__nor2_8 _3070_ (.A(net204),
    .B(_2652_),
    .Y(_2653_));
 sky130_fd_sc_hd__nand2_2 _3071_ (.A(net224),
    .B(_2651_),
    .Y(_2654_));
 sky130_fd_sc_hd__nand2_8 _3072_ (.A(net201),
    .B(_2653_),
    .Y(_2655_));
 sky130_fd_sc_hd__nor2_4 _3073_ (.A(_2648_),
    .B(_2655_),
    .Y(_2656_));
 sky130_fd_sc_hd__or2_4 _3074_ (.A(_2648_),
    .B(_2655_),
    .X(_2657_));
 sky130_fd_sc_hd__and2b_4 _3075_ (.A_N(net298),
    .B(net299),
    .X(_2658_));
 sky130_fd_sc_hd__nand2b_4 _3076_ (.A_N(net298),
    .B(net299),
    .Y(_2659_));
 sky130_fd_sc_hd__nor2_2 _3077_ (.A(net301),
    .B(_2659_),
    .Y(_2660_));
 sky130_fd_sc_hd__or2_4 _3078_ (.A(net301),
    .B(_2659_),
    .X(_2661_));
 sky130_fd_sc_hd__and3_4 _3079_ (.A(net209),
    .B(net227),
    .C(_2660_),
    .X(_2662_));
 sky130_fd_sc_hd__or3_4 _3080_ (.A(net302),
    .B(net204),
    .C(_2661_),
    .X(_2663_));
 sky130_fd_sc_hd__nand2_8 _3081_ (.A(net207),
    .B(_2662_),
    .Y(_2664_));
 sky130_fd_sc_hd__nor2_4 _3082_ (.A(_2648_),
    .B(_2664_),
    .Y(_2665_));
 sky130_fd_sc_hd__or2_4 _3083_ (.A(_2648_),
    .B(_2664_),
    .X(_2666_));
 sky130_fd_sc_hd__nand2_8 _3084_ (.A(_2525_),
    .B(_2645_),
    .Y(_2667_));
 sky130_fd_sc_hd__and2_4 _3085_ (.A(_2537_),
    .B(net290),
    .X(_2668_));
 sky130_fd_sc_hd__nand2_2 _3086_ (.A(\as2650.cycle[6] ),
    .B(_2562_),
    .Y(_2669_));
 sky130_fd_sc_hd__or3b_4 _3087_ (.A(_2669_),
    .B(\as2650.cycle[1] ),
    .C_N(net290),
    .X(_2670_));
 sky130_fd_sc_hd__nor2_4 _3088_ (.A(_2536_),
    .B(_2670_),
    .Y(_2671_));
 sky130_fd_sc_hd__or2_1 _3089_ (.A(_2536_),
    .B(_2670_),
    .X(_2672_));
 sky130_fd_sc_hd__or2_4 _3090_ (.A(net294),
    .B(net72),
    .X(_2673_));
 sky130_fd_sc_hd__nand2_4 _3091_ (.A(net204),
    .B(_2560_),
    .Y(_2674_));
 sky130_fd_sc_hd__nor2_8 _3092_ (.A(\as2650.addr_buff[6] ),
    .B(\as2650.addr_buff[5] ),
    .Y(_2675_));
 sky130_fd_sc_hd__nor2_8 _3093_ (.A(net223),
    .B(_2675_),
    .Y(_2676_));
 sky130_fd_sc_hd__nand2_8 _3094_ (.A(_2560_),
    .B(_2676_),
    .Y(_2677_));
 sky130_fd_sc_hd__nor3_2 _3095_ (.A(_2667_),
    .B(_2673_),
    .C(_2677_),
    .Y(_2678_));
 sky130_fd_sc_hd__or2_4 _3096_ (.A(net303),
    .B(_2600_),
    .X(_2679_));
 sky130_fd_sc_hd__nor2_4 _3097_ (.A(net297),
    .B(_2679_),
    .Y(_2680_));
 sky130_fd_sc_hd__or2_4 _3098_ (.A(net297),
    .B(_2679_),
    .X(_2681_));
 sky130_fd_sc_hd__nand2_4 _3099_ (.A(net206),
    .B(net115),
    .Y(_2682_));
 sky130_fd_sc_hd__or3_4 _3100_ (.A(_2561_),
    .B(_2610_),
    .C(_2682_),
    .X(_2683_));
 sky130_fd_sc_hd__nor2_1 _3101_ (.A(\as2650.cycle[7] ),
    .B(_2670_),
    .Y(_2684_));
 sky130_fd_sc_hd__or2_4 _3102_ (.A(\as2650.cycle[7] ),
    .B(_2670_),
    .X(_2685_));
 sky130_fd_sc_hd__nor2_4 _3103_ (.A(\as2650.idx_ctrl[1] ),
    .B(\as2650.idx_ctrl[0] ),
    .Y(_2686_));
 sky130_fd_sc_hd__or2_4 _3104_ (.A(\as2650.idx_ctrl[1] ),
    .B(\as2650.idx_ctrl[0] ),
    .X(_2687_));
 sky130_fd_sc_hd__or3_4 _3105_ (.A(_2674_),
    .B(_2685_),
    .C(_2686_),
    .X(_2688_));
 sky130_fd_sc_hd__nor2_8 _3106_ (.A(net206),
    .B(net139),
    .Y(_2689_));
 sky130_fd_sc_hd__or2_4 _3107_ (.A(_2545_),
    .B(net143),
    .X(_2690_));
 sky130_fd_sc_hd__o311a_1 _3108_ (.A1(_2561_),
    .A2(_2649_),
    .A3(_2690_),
    .B1(_2688_),
    .C1(_2683_),
    .X(_2691_));
 sky130_fd_sc_hd__nand2_2 _3109_ (.A(net202),
    .B(_2651_),
    .Y(_2692_));
 sky130_fd_sc_hd__or2_4 _3110_ (.A(net197),
    .B(_2692_),
    .X(_2693_));
 sky130_fd_sc_hd__nor2_4 _3111_ (.A(_2648_),
    .B(_2693_),
    .Y(_2694_));
 sky130_fd_sc_hd__or2_4 _3112_ (.A(_2648_),
    .B(_2693_),
    .X(_2695_));
 sky130_fd_sc_hd__nand2_8 _3113_ (.A(net203),
    .B(net132),
    .Y(_2696_));
 sky130_fd_sc_hd__and3_2 _3114_ (.A(net301),
    .B(\as2650.ins_reg[6] ),
    .C(net297),
    .X(_2697_));
 sky130_fd_sc_hd__or4_4 _3115_ (.A(net201),
    .B(net177),
    .C(_2687_),
    .D(_2697_),
    .X(_2698_));
 sky130_fd_sc_hd__nor2_4 _3116_ (.A(_2667_),
    .B(_2683_),
    .Y(_2699_));
 sky130_fd_sc_hd__or2_2 _3117_ (.A(_2667_),
    .B(_2683_),
    .X(_2700_));
 sky130_fd_sc_hd__nand2_4 _3118_ (.A(net261),
    .B(net178),
    .Y(_2701_));
 sky130_fd_sc_hd__and2b_4 _3119_ (.A_N(net306),
    .B(net305),
    .X(_2702_));
 sky130_fd_sc_hd__mux2_8 _3120_ (.A0(\as2650.r123[2][0] ),
    .A1(\as2650.r123_2[2][0] ),
    .S(net211),
    .X(_2703_));
 sky130_fd_sc_hd__xor2_4 _3121_ (.A(net305),
    .B(net306),
    .X(_2704_));
 sky130_fd_sc_hd__mux4_2 _3122_ (.A0(\as2650.r123[1][0] ),
    .A1(\as2650.r123[0][0] ),
    .A2(\as2650.r123_2[1][0] ),
    .A3(\as2650.r123_2[0][0] ),
    .S0(net306),
    .S1(net213),
    .X(_2705_));
 sky130_fd_sc_hd__a22oi_4 _3123_ (.A1(net196),
    .A2(_2703_),
    .B1(_2704_),
    .B2(_2705_),
    .Y(_2706_));
 sky130_fd_sc_hd__and2_4 _3124_ (.A(_2701_),
    .B(_2706_),
    .X(_2707_));
 sky130_fd_sc_hd__nand2_2 _3125_ (.A(_2701_),
    .B(_2706_),
    .Y(_2708_));
 sky130_fd_sc_hd__xnor2_4 _3126_ (.A(_2650_),
    .B(_2707_),
    .Y(_2709_));
 sky130_fd_sc_hd__or3_4 _3127_ (.A(_2561_),
    .B(net117),
    .C(_2682_),
    .X(_2710_));
 sky130_fd_sc_hd__or2_2 _3128_ (.A(_2667_),
    .B(_2710_),
    .X(_2711_));
 sky130_fd_sc_hd__mux2_1 _3129_ (.A0(net350),
    .A1(_2709_),
    .S(_2700_),
    .X(_2712_));
 sky130_fd_sc_hd__or2_1 _3130_ (.A(_2665_),
    .B(_2712_),
    .X(_2713_));
 sky130_fd_sc_hd__mux4_1 _3131_ (.A0(\as2650.r123[1][1] ),
    .A1(\as2650.r123[0][1] ),
    .A2(\as2650.r123_2[1][1] ),
    .A3(\as2650.r123_2[0][1] ),
    .S0(net306),
    .S1(net214),
    .X(_2714_));
 sky130_fd_sc_hd__mux2_4 _3132_ (.A0(\as2650.r123[2][1] ),
    .A1(\as2650.r123_2[2][1] ),
    .S(net211),
    .X(_2715_));
 sky130_fd_sc_hd__and2_2 _3133_ (.A(net196),
    .B(_2715_),
    .X(_2716_));
 sky130_fd_sc_hd__a22o_2 _3134_ (.A1(net257),
    .A2(net178),
    .B1(_2704_),
    .B2(_2714_),
    .X(_2717_));
 sky130_fd_sc_hd__or2_4 _3135_ (.A(_2716_),
    .B(_2717_),
    .X(_2718_));
 sky130_fd_sc_hd__o211a_1 _3136_ (.A1(_2666_),
    .A2(_2718_),
    .B1(_2713_),
    .C1(_2657_),
    .X(_2719_));
 sky130_fd_sc_hd__nand2_4 _3137_ (.A(\as2650.psl[3] ),
    .B(_2526_),
    .Y(_2720_));
 sky130_fd_sc_hd__mux2_4 _3138_ (.A0(\as2650.r123[2][7] ),
    .A1(\as2650.r123_2[2][7] ),
    .S(net211),
    .X(_2721_));
 sky130_fd_sc_hd__mux2_4 _3139_ (.A0(\as2650.r123[0][7] ),
    .A1(\as2650.r123_2[0][7] ),
    .S(net211),
    .X(_2722_));
 sky130_fd_sc_hd__mux4_1 _3140_ (.A0(\as2650.r123[1][7] ),
    .A1(\as2650.r123[0][7] ),
    .A2(\as2650.r123_2[1][7] ),
    .A3(\as2650.r123_2[0][7] ),
    .S0(net307),
    .S1(net211),
    .X(_2723_));
 sky130_fd_sc_hd__a22o_1 _3141_ (.A1(net196),
    .A2(_2721_),
    .B1(_2723_),
    .B2(_2704_),
    .X(_2724_));
 sky130_fd_sc_hd__a21o_2 _3142_ (.A1(net234),
    .A2(net177),
    .B1(_2724_),
    .X(_2725_));
 sky130_fd_sc_hd__nand2_1 _3143_ (.A(\as2650.psl[3] ),
    .B(\as2650.carry ),
    .Y(_2726_));
 sky130_fd_sc_hd__o21a_2 _3144_ (.A1(\as2650.psl[3] ),
    .A2(net109),
    .B1(_2720_),
    .X(_2727_));
 sky130_fd_sc_hd__inv_2 _3145_ (.A(_2727_),
    .Y(_2728_));
 sky130_fd_sc_hd__a211o_1 _3146_ (.A1(_2656_),
    .A2(_2727_),
    .B1(_2719_),
    .C1(_2694_),
    .X(_2729_));
 sky130_fd_sc_hd__nor2_8 _3147_ (.A(_2667_),
    .B(_2688_),
    .Y(_2730_));
 sky130_fd_sc_hd__or2_1 _3148_ (.A(_2667_),
    .B(_2688_),
    .X(_2731_));
 sky130_fd_sc_hd__and2b_2 _3149_ (.A_N(\as2650.addr_buff[6] ),
    .B(\as2650.addr_buff[5] ),
    .X(_2732_));
 sky130_fd_sc_hd__nand2b_4 _3150_ (.A_N(\as2650.addr_buff[6] ),
    .B(\as2650.addr_buff[5] ),
    .Y(_2733_));
 sky130_fd_sc_hd__nand2b_4 _3151_ (.A_N(\as2650.addr_buff[5] ),
    .B(\as2650.addr_buff[6] ),
    .Y(_2734_));
 sky130_fd_sc_hd__nand2_8 _3152_ (.A(_2733_),
    .B(_2734_),
    .Y(_2735_));
 sky130_fd_sc_hd__xnor2_4 _3153_ (.A(_2707_),
    .B(_2735_),
    .Y(_2736_));
 sky130_fd_sc_hd__or3_4 _3154_ (.A(_2667_),
    .B(_2673_),
    .C(_2677_),
    .X(_2737_));
 sky130_fd_sc_hd__o21a_1 _3155_ (.A1(net262),
    .A2(_2695_),
    .B1(_2737_),
    .X(_2738_));
 sky130_fd_sc_hd__nor3_4 _3156_ (.A(_2667_),
    .B(_2673_),
    .C(_2677_),
    .Y(_2739_));
 sky130_fd_sc_hd__a22o_1 _3157_ (.A1(_2729_),
    .A2(_2738_),
    .B1(_2739_),
    .B2(_2736_),
    .X(_2740_));
 sky130_fd_sc_hd__or3_2 _3158_ (.A(_2674_),
    .B(_2685_),
    .C(_2686_),
    .X(_2741_));
 sky130_fd_sc_hd__and2b_4 _3159_ (.A_N(\as2650.idx_ctrl[1] ),
    .B(\as2650.idx_ctrl[0] ),
    .X(_2742_));
 sky130_fd_sc_hd__nand2b_4 _3160_ (.A_N(\as2650.idx_ctrl[1] ),
    .B(\as2650.idx_ctrl[0] ),
    .Y(_2743_));
 sky130_fd_sc_hd__nand2b_4 _3161_ (.A_N(\as2650.idx_ctrl[0] ),
    .B(\as2650.idx_ctrl[1] ),
    .Y(_2744_));
 sky130_fd_sc_hd__nand2_8 _3162_ (.A(_2743_),
    .B(_2744_),
    .Y(_2745_));
 sky130_fd_sc_hd__xnor2_4 _3163_ (.A(_2707_),
    .B(_2745_),
    .Y(_2746_));
 sky130_fd_sc_hd__or4_2 _3164_ (.A(net213),
    .B(_2561_),
    .C(_2696_),
    .D(_2698_),
    .X(_2747_));
 sky130_fd_sc_hd__mux2_1 _3165_ (.A0(_2740_),
    .A1(_2746_),
    .S(_2730_),
    .X(_2748_));
 sky130_fd_sc_hd__nor4_4 _3166_ (.A(net213),
    .B(_2597_),
    .C(_2674_),
    .D(_2698_),
    .Y(_2749_));
 sky130_fd_sc_hd__nor2_1 _3167_ (.A(\as2650.holding_reg[0] ),
    .B(net197),
    .Y(_2750_));
 sky130_fd_sc_hd__a31o_4 _3168_ (.A1(net197),
    .A2(_2701_),
    .A3(_2706_),
    .B1(_2750_),
    .X(_2751_));
 sky130_fd_sc_hd__inv_2 _3169_ (.A(_2751_),
    .Y(_2752_));
 sky130_fd_sc_hd__nor2_1 _3170_ (.A(\as2650.holding_reg[0] ),
    .B(net199),
    .Y(_2753_));
 sky130_fd_sc_hd__a31o_4 _3171_ (.A1(net199),
    .A2(_2701_),
    .A3(_2706_),
    .B1(_2753_),
    .X(_2754_));
 sky130_fd_sc_hd__nor2_1 _3172_ (.A(_2752_),
    .B(_2754_),
    .Y(_2755_));
 sky130_fd_sc_hd__and2_1 _3173_ (.A(\as2650.holding_reg[0] ),
    .B(net113),
    .X(_2756_));
 sky130_fd_sc_hd__or2_1 _3174_ (.A(_2751_),
    .B(_2756_),
    .X(_2757_));
 sky130_fd_sc_hd__xnor2_4 _3175_ (.A(_2751_),
    .B(_2754_),
    .Y(_2758_));
 sky130_fd_sc_hd__nor2_4 _3176_ (.A(net301),
    .B(_2586_),
    .Y(_2759_));
 sky130_fd_sc_hd__or2_4 _3177_ (.A(net301),
    .B(_2586_),
    .X(_2760_));
 sky130_fd_sc_hd__a21oi_1 _3178_ (.A1(_2726_),
    .A2(_2758_),
    .B1(_2760_),
    .Y(_2761_));
 sky130_fd_sc_hd__o21a_1 _3179_ (.A1(_2726_),
    .A2(_2758_),
    .B1(_2761_),
    .X(_2762_));
 sky130_fd_sc_hd__nand2_1 _3180_ (.A(_2720_),
    .B(_2758_),
    .Y(_2763_));
 sky130_fd_sc_hd__and2_2 _3181_ (.A(net301),
    .B(net195),
    .X(_2764_));
 sky130_fd_sc_hd__nand2_4 _3182_ (.A(net301),
    .B(net195),
    .Y(_2765_));
 sky130_fd_sc_hd__o2111a_1 _3183_ (.A1(_2720_),
    .A2(_2758_),
    .B1(_2763_),
    .C1(net195),
    .D1(\as2650.ins_reg[5] ),
    .X(_2766_));
 sky130_fd_sc_hd__o221a_1 _3184_ (.A1(_2659_),
    .A2(_2751_),
    .B1(_2754_),
    .B2(net195),
    .C1(net160),
    .X(_2767_));
 sky130_fd_sc_hd__or3b_1 _3185_ (.A(_2762_),
    .B(_2766_),
    .C_N(_2767_),
    .X(_2768_));
 sky130_fd_sc_hd__nand2_4 _3186_ (.A(\as2650.ins_reg[5] ),
    .B(_2571_),
    .Y(_2769_));
 sky130_fd_sc_hd__o21a_1 _3187_ (.A1(_2661_),
    .A2(_2756_),
    .B1(net159),
    .X(_2770_));
 sky130_fd_sc_hd__a2bb2o_4 _3188_ (.A1_N(_2758_),
    .A2_N(net159),
    .B1(_2770_),
    .B2(_2768_),
    .X(_2771_));
 sky130_fd_sc_hd__mux2_8 _3189_ (.A0(_2748_),
    .A1(_2771_),
    .S(net71),
    .X(_2772_));
 sky130_fd_sc_hd__nand2_1 _3190_ (.A(net226),
    .B(_2759_),
    .Y(_2773_));
 sky130_fd_sc_hd__and4_4 _3191_ (.A(net227),
    .B(net200),
    .C(_2577_),
    .D(_2759_),
    .X(_2774_));
 sky130_fd_sc_hd__or3_4 _3192_ (.A(net197),
    .B(_2578_),
    .C(_2773_),
    .X(_2775_));
 sky130_fd_sc_hd__nand2_4 _3193_ (.A(net201),
    .B(net177),
    .Y(_2776_));
 sky130_fd_sc_hd__nor2_1 _3194_ (.A(_2574_),
    .B(_2776_),
    .Y(_2777_));
 sky130_fd_sc_hd__or2_4 _3195_ (.A(_2574_),
    .B(_2776_),
    .X(_2778_));
 sky130_fd_sc_hd__nor2_1 _3196_ (.A(_2774_),
    .B(net69),
    .Y(_2779_));
 sky130_fd_sc_hd__nand2_4 _3197_ (.A(_2775_),
    .B(net66),
    .Y(_2780_));
 sky130_fd_sc_hd__nor2_2 _3198_ (.A(net293),
    .B(_2779_),
    .Y(_2781_));
 sky130_fd_sc_hd__or3_1 _3199_ (.A(_2561_),
    .B(_2649_),
    .C(_2690_),
    .X(_2782_));
 sky130_fd_sc_hd__and3_2 _3200_ (.A(_2683_),
    .B(_2741_),
    .C(_2782_),
    .X(_2783_));
 sky130_fd_sc_hd__and4_1 _3201_ (.A(_2657_),
    .B(_2666_),
    .C(_2695_),
    .D(_2737_),
    .X(_2784_));
 sky130_fd_sc_hd__o211a_4 _3202_ (.A1(_2667_),
    .A2(_2783_),
    .B1(_2784_),
    .C1(_2747_),
    .X(_2785_));
 sky130_fd_sc_hd__or2_2 _3203_ (.A(net305),
    .B(_2785_),
    .X(_2786_));
 sky130_fd_sc_hd__inv_6 _3204_ (.A(_2786_),
    .Y(_2787_));
 sky130_fd_sc_hd__a211oi_4 _3205_ (.A1(_2646_),
    .A2(_2781_),
    .B1(_2787_),
    .C1(net347),
    .Y(_2788_));
 sky130_fd_sc_hd__a211o_4 _3206_ (.A1(_2646_),
    .A2(_2781_),
    .B1(_2787_),
    .C1(net348),
    .X(_2789_));
 sky130_fd_sc_hd__nor2_1 _3207_ (.A(net215),
    .B(net218),
    .Y(_2790_));
 sky130_fd_sc_hd__or2_2 _3208_ (.A(net215),
    .B(net217),
    .X(_2791_));
 sky130_fd_sc_hd__nor2_2 _3209_ (.A(net219),
    .B(net172),
    .Y(_2792_));
 sky130_fd_sc_hd__nand2_8 _3210_ (.A(net220),
    .B(net172),
    .Y(_2793_));
 sky130_fd_sc_hd__and3_1 _3211_ (.A(net219),
    .B(\as2650.stack[3][8] ),
    .C(net173),
    .X(_2794_));
 sky130_fd_sc_hd__nand2_1 _3212_ (.A(net215),
    .B(_2528_),
    .Y(_2795_));
 sky130_fd_sc_hd__nor2_1 _3213_ (.A(_2527_),
    .B(_2528_),
    .Y(_2796_));
 sky130_fd_sc_hd__nand2_2 _3214_ (.A(net215),
    .B(net217),
    .Y(_2797_));
 sky130_fd_sc_hd__nor2_1 _3215_ (.A(net173),
    .B(_2796_),
    .Y(_2798_));
 sky130_fd_sc_hd__o22a_1 _3216_ (.A1(\as2650.stack[1][8] ),
    .A2(net167),
    .B1(net156),
    .B2(\as2650.stack[0][8] ),
    .X(_2799_));
 sky130_fd_sc_hd__and2b_4 _3217_ (.A_N(net158),
    .B(_2793_),
    .X(_2800_));
 sky130_fd_sc_hd__nand2b_4 _3218_ (.A_N(net158),
    .B(_2793_),
    .Y(_2801_));
 sky130_fd_sc_hd__o221a_1 _3219_ (.A1(net158),
    .A2(_2794_),
    .B1(_2797_),
    .B2(\as2650.stack[2][8] ),
    .C1(_2799_),
    .X(_2802_));
 sky130_fd_sc_hd__mux4_2 _3220_ (.A0(\as2650.stack[7][8] ),
    .A1(\as2650.stack[4][8] ),
    .A2(\as2650.stack[5][8] ),
    .A3(\as2650.stack[6][8] ),
    .S0(net215),
    .S1(net217),
    .X(_2803_));
 sky130_fd_sc_hd__a21o_4 _3221_ (.A1(net107),
    .A2(_2803_),
    .B1(_2802_),
    .X(_2804_));
 sky130_fd_sc_hd__or2_4 _3222_ (.A(_2773_),
    .B(_2776_),
    .X(_2805_));
 sky130_fd_sc_hd__or3_4 _3223_ (.A(net304),
    .B(net197),
    .C(_2773_),
    .X(_2806_));
 sky130_fd_sc_hd__and2_4 _3224_ (.A(net66),
    .B(_2806_),
    .X(_2807_));
 sky130_fd_sc_hd__nand2_1 _3225_ (.A(net66),
    .B(_2806_),
    .Y(_2808_));
 sky130_fd_sc_hd__nor2_8 _3226_ (.A(_2647_),
    .B(_2807_),
    .Y(_2809_));
 sky130_fd_sc_hd__nor2_4 _3227_ (.A(net143),
    .B(net66),
    .Y(_2810_));
 sky130_fd_sc_hd__or4b_1 _3228_ (.A(net212),
    .B(_2561_),
    .C(_2804_),
    .D_N(_2810_),
    .X(_2811_));
 sky130_fd_sc_hd__o211a_1 _3229_ (.A1(net260),
    .A2(net69),
    .B1(_2809_),
    .C1(_2811_),
    .X(_2812_));
 sky130_fd_sc_hd__a211o_1 _3230_ (.A1(_2772_),
    .A2(_2787_),
    .B1(_2788_),
    .C1(_2812_),
    .X(_2813_));
 sky130_fd_sc_hd__o21a_1 _3231_ (.A1(\as2650.r123[0][0] ),
    .A2(_2789_),
    .B1(_2813_),
    .X(_0007_));
 sky130_fd_sc_hd__or2_1 _3232_ (.A(net254),
    .B(net69),
    .X(_2814_));
 sky130_fd_sc_hd__mux4_1 _3233_ (.A0(\as2650.stack[7][9] ),
    .A1(\as2650.stack[4][9] ),
    .A2(\as2650.stack[5][9] ),
    .A3(\as2650.stack[6][9] ),
    .S0(net215),
    .S1(net217),
    .X(_2815_));
 sky130_fd_sc_hd__o22a_1 _3234_ (.A1(\as2650.stack[1][9] ),
    .A2(net166),
    .B1(net156),
    .B2(\as2650.stack[0][9] ),
    .X(_2816_));
 sky130_fd_sc_hd__o221a_1 _3235_ (.A1(\as2650.stack[3][9] ),
    .A2(net171),
    .B1(_2797_),
    .B2(\as2650.stack[2][9] ),
    .C1(_2816_),
    .X(_2817_));
 sky130_fd_sc_hd__mux2_4 _3236_ (.A0(_2815_),
    .A1(_2817_),
    .S(_2801_),
    .X(_2818_));
 sky130_fd_sc_hd__o211a_1 _3237_ (.A1(net66),
    .A2(_2818_),
    .B1(_2814_),
    .C1(_2809_),
    .X(_2819_));
 sky130_fd_sc_hd__nor2_4 _3238_ (.A(_2599_),
    .B(_2600_),
    .Y(_2820_));
 sky130_fd_sc_hd__mux2_4 _3239_ (.A0(_2653_),
    .A1(_2820_),
    .S(_2707_),
    .X(_2821_));
 sky130_fd_sc_hd__xor2_4 _3240_ (.A(net112),
    .B(_2821_),
    .X(_2822_));
 sky130_fd_sc_hd__mux2_4 _3241_ (.A0(\as2650.r123[2][2] ),
    .A1(\as2650.r123_2[2][2] ),
    .S(net210),
    .X(_2823_));
 sky130_fd_sc_hd__mux4_1 _3242_ (.A0(\as2650.r123[1][2] ),
    .A1(\as2650.r123[0][2] ),
    .A2(\as2650.r123_2[1][2] ),
    .A3(\as2650.r123_2[0][2] ),
    .S0(net307),
    .S1(net212),
    .X(_2824_));
 sky130_fd_sc_hd__a22o_1 _3243_ (.A1(net196),
    .A2(_2823_),
    .B1(_2824_),
    .B2(_2704_),
    .X(_2825_));
 sky130_fd_sc_hd__a21o_4 _3244_ (.A1(net251),
    .A2(net177),
    .B1(_2825_),
    .X(_2826_));
 sky130_fd_sc_hd__a221o_1 _3245_ (.A1(net345),
    .A2(_2699_),
    .B1(_2711_),
    .B2(_2822_),
    .C1(_2665_),
    .X(_2827_));
 sky130_fd_sc_hd__o21a_1 _3246_ (.A1(_2666_),
    .A2(net105),
    .B1(_2657_),
    .X(_2828_));
 sky130_fd_sc_hd__a221o_1 _3247_ (.A1(_2656_),
    .A2(net113),
    .B1(_2827_),
    .B2(_2828_),
    .C1(_2694_),
    .X(_2829_));
 sky130_fd_sc_hd__o2bb2a_4 _3248_ (.A1_N(_2701_),
    .A2_N(_2706_),
    .B1(_2716_),
    .B2(_2717_),
    .X(_2830_));
 sky130_fd_sc_hd__nor2_1 _3249_ (.A(net113),
    .B(net112),
    .Y(_2831_));
 sky130_fd_sc_hd__xnor2_4 _3250_ (.A(net113),
    .B(net112),
    .Y(_2832_));
 sky130_fd_sc_hd__o21ai_4 _3251_ (.A1(_2707_),
    .A2(_2732_),
    .B1(_2734_),
    .Y(_2833_));
 sky130_fd_sc_hd__xnor2_4 _3252_ (.A(_2832_),
    .B(_2833_),
    .Y(_2834_));
 sky130_fd_sc_hd__o21a_1 _3253_ (.A1(net258),
    .A2(_2695_),
    .B1(_2737_),
    .X(_2835_));
 sky130_fd_sc_hd__a22o_1 _3254_ (.A1(_2739_),
    .A2(_2834_),
    .B1(_2835_),
    .B2(_2829_),
    .X(_2836_));
 sky130_fd_sc_hd__o21ai_4 _3255_ (.A1(_2707_),
    .A2(_2742_),
    .B1(_2744_),
    .Y(_2837_));
 sky130_fd_sc_hd__xnor2_4 _3256_ (.A(_2832_),
    .B(_2837_),
    .Y(_2838_));
 sky130_fd_sc_hd__mux2_1 _3257_ (.A0(_2836_),
    .A1(_2838_),
    .S(_2730_),
    .X(_2839_));
 sky130_fd_sc_hd__and2_1 _3258_ (.A(\as2650.holding_reg[1] ),
    .B(net111),
    .X(_2840_));
 sky130_fd_sc_hd__or2_1 _3259_ (.A(\as2650.holding_reg[1] ),
    .B(net111),
    .X(_2841_));
 sky130_fd_sc_hd__and2b_4 _3260_ (.A_N(_2840_),
    .B(_2841_),
    .X(_2842_));
 sky130_fd_sc_hd__o21bai_2 _3261_ (.A1(_2726_),
    .A2(_2758_),
    .B1_N(_2756_),
    .Y(_2843_));
 sky130_fd_sc_hd__xor2_1 _3262_ (.A(_2842_),
    .B(_2843_),
    .X(_2844_));
 sky130_fd_sc_hd__a21oi_2 _3263_ (.A1(_2757_),
    .A2(_2763_),
    .B1(_2842_),
    .Y(_2845_));
 sky130_fd_sc_hd__and3_1 _3264_ (.A(_2757_),
    .B(_2763_),
    .C(_2842_),
    .X(_2846_));
 sky130_fd_sc_hd__o21ai_1 _3265_ (.A1(_2845_),
    .A2(_2846_),
    .B1(_2764_),
    .Y(_2847_));
 sky130_fd_sc_hd__mux2_1 _3266_ (.A0(\as2650.holding_reg[1] ),
    .A1(net111),
    .S(net199),
    .X(_2848_));
 sky130_fd_sc_hd__o221a_1 _3267_ (.A1(_2760_),
    .A2(_2844_),
    .B1(_2848_),
    .B2(net195),
    .C1(_2847_),
    .X(_2849_));
 sky130_fd_sc_hd__or2_1 _3268_ (.A(net160),
    .B(_2840_),
    .X(_2850_));
 sky130_fd_sc_hd__nand2_8 _3269_ (.A(\as2650.ins_reg[5] ),
    .B(_2658_),
    .Y(_2851_));
 sky130_fd_sc_hd__o221a_4 _3270_ (.A1(_2658_),
    .A2(_2849_),
    .B1(_2851_),
    .B2(_2841_),
    .C1(_2850_),
    .X(_2852_));
 sky130_fd_sc_hd__or2_1 _3271_ (.A(\as2650.holding_reg[1] ),
    .B(net197),
    .X(_2853_));
 sky130_fd_sc_hd__o21ai_2 _3272_ (.A1(net199),
    .A2(net111),
    .B1(_2853_),
    .Y(_2854_));
 sky130_fd_sc_hd__or2_4 _3273_ (.A(net159),
    .B(_2854_),
    .X(_2855_));
 sky130_fd_sc_hd__xnor2_4 _3274_ (.A(_2852_),
    .B(_2855_),
    .Y(_2856_));
 sky130_fd_sc_hd__mux2_8 _3275_ (.A0(_2839_),
    .A1(_2856_),
    .S(net71),
    .X(_2857_));
 sky130_fd_sc_hd__a211o_1 _3276_ (.A1(_2787_),
    .A2(_2857_),
    .B1(_2819_),
    .C1(_2788_),
    .X(_2858_));
 sky130_fd_sc_hd__o21a_1 _3277_ (.A1(\as2650.r123[0][1] ),
    .A2(_2789_),
    .B1(_2858_),
    .X(_0008_));
 sky130_fd_sc_hd__or2_1 _3278_ (.A(net251),
    .B(net68),
    .X(_2859_));
 sky130_fd_sc_hd__and3_1 _3279_ (.A(net221),
    .B(\as2650.stack[3][10] ),
    .C(net173),
    .X(_2860_));
 sky130_fd_sc_hd__o22a_1 _3280_ (.A1(\as2650.stack[1][10] ),
    .A2(net167),
    .B1(net155),
    .B2(\as2650.stack[0][10] ),
    .X(_2861_));
 sky130_fd_sc_hd__o221a_1 _3281_ (.A1(\as2650.stack[2][10] ),
    .A2(net169),
    .B1(_2860_),
    .B2(net158),
    .C1(_2861_),
    .X(_2862_));
 sky130_fd_sc_hd__o22a_1 _3282_ (.A1(\as2650.stack[4][10] ),
    .A2(net156),
    .B1(net170),
    .B2(\as2650.stack[6][10] ),
    .X(_2863_));
 sky130_fd_sc_hd__o22a_1 _3283_ (.A1(\as2650.stack[5][10] ),
    .A2(net167),
    .B1(net171),
    .B2(\as2650.stack[7][10] ),
    .X(_2864_));
 sky130_fd_sc_hd__a31o_2 _3284_ (.A1(net108),
    .A2(_2863_),
    .A3(_2864_),
    .B1(_2862_),
    .X(_2865_));
 sky130_fd_sc_hd__o211a_1 _3285_ (.A1(net67),
    .A2(_2865_),
    .B1(_2859_),
    .C1(_2809_),
    .X(_2866_));
 sky130_fd_sc_hd__a22o_2 _3286_ (.A1(_2653_),
    .A2(_2830_),
    .B1(_2831_),
    .B2(_2820_),
    .X(_2867_));
 sky130_fd_sc_hd__nor3_2 _3287_ (.A(net113),
    .B(net112),
    .C(net104),
    .Y(_2868_));
 sky130_fd_sc_hd__and3_1 _3288_ (.A(_2653_),
    .B(net104),
    .C(_2830_),
    .X(_2869_));
 sky130_fd_sc_hd__xor2_4 _3289_ (.A(net105),
    .B(_2867_),
    .X(_2870_));
 sky130_fd_sc_hd__mux2_4 _3290_ (.A0(\as2650.r123[2][3] ),
    .A1(\as2650.r123_2[2][3] ),
    .S(net210),
    .X(_2871_));
 sky130_fd_sc_hd__mux4_1 _3291_ (.A0(\as2650.r123[1][3] ),
    .A1(\as2650.r123[0][3] ),
    .A2(\as2650.r123_2[1][3] ),
    .A3(\as2650.r123_2[0][3] ),
    .S0(net307),
    .S1(net210),
    .X(_2872_));
 sky130_fd_sc_hd__a22o_1 _3292_ (.A1(net247),
    .A2(net178),
    .B1(_2704_),
    .B2(_2872_),
    .X(_2873_));
 sky130_fd_sc_hd__a21o_4 _3293_ (.A1(net196),
    .A2(_2871_),
    .B1(_2873_),
    .X(_2874_));
 sky130_fd_sc_hd__a221o_1 _3294_ (.A1(net342),
    .A2(_2699_),
    .B1(_2711_),
    .B2(_2870_),
    .C1(_2665_),
    .X(_2875_));
 sky130_fd_sc_hd__o211a_1 _3295_ (.A1(_2666_),
    .A2(_2874_),
    .B1(_2875_),
    .C1(_2657_),
    .X(_2876_));
 sky130_fd_sc_hd__a211o_1 _3296_ (.A1(_2656_),
    .A2(net111),
    .B1(_2876_),
    .C1(_2694_),
    .X(_2877_));
 sky130_fd_sc_hd__xor2_1 _3297_ (.A(net104),
    .B(_2830_),
    .X(_2878_));
 sky130_fd_sc_hd__or2_1 _3298_ (.A(_2733_),
    .B(_2878_),
    .X(_2879_));
 sky130_fd_sc_hd__o21a_1 _3299_ (.A1(net113),
    .A2(net112),
    .B1(net104),
    .X(_2880_));
 sky130_fd_sc_hd__or2_2 _3300_ (.A(_2868_),
    .B(_2880_),
    .X(_2881_));
 sky130_fd_sc_hd__o221a_4 _3301_ (.A1(_2735_),
    .A2(net104),
    .B1(_2881_),
    .B2(_2734_),
    .C1(_2879_),
    .X(_2882_));
 sky130_fd_sc_hd__o21a_1 _3302_ (.A1(net253),
    .A2(_2695_),
    .B1(_2737_),
    .X(_2883_));
 sky130_fd_sc_hd__a22o_1 _3303_ (.A1(_2739_),
    .A2(_2882_),
    .B1(_2883_),
    .B2(_2877_),
    .X(_2884_));
 sky130_fd_sc_hd__or2_1 _3304_ (.A(_2743_),
    .B(_2878_),
    .X(_2885_));
 sky130_fd_sc_hd__o221a_4 _3305_ (.A1(_2745_),
    .A2(net104),
    .B1(_2881_),
    .B2(_2744_),
    .C1(_2885_),
    .X(_2886_));
 sky130_fd_sc_hd__mux2_1 _3306_ (.A0(_2884_),
    .A1(_2886_),
    .S(_2730_),
    .X(_2887_));
 sky130_fd_sc_hd__or2_2 _3307_ (.A(\as2650.holding_reg[2] ),
    .B(net106),
    .X(_2888_));
 sky130_fd_sc_hd__nand2_2 _3308_ (.A(\as2650.holding_reg[2] ),
    .B(net106),
    .Y(_2889_));
 sky130_fd_sc_hd__and2_2 _3309_ (.A(_2888_),
    .B(_2889_),
    .X(_2890_));
 sky130_fd_sc_hd__a21o_1 _3310_ (.A1(_2842_),
    .A2(_2843_),
    .B1(_2840_),
    .X(_2891_));
 sky130_fd_sc_hd__nand2_1 _3311_ (.A(_2890_),
    .B(_2891_),
    .Y(_2892_));
 sky130_fd_sc_hd__or2_1 _3312_ (.A(_2890_),
    .B(_2891_),
    .X(_2893_));
 sky130_fd_sc_hd__a21o_1 _3313_ (.A1(_2892_),
    .A2(_2893_),
    .B1(_2760_),
    .X(_2894_));
 sky130_fd_sc_hd__nor2_1 _3314_ (.A(_2840_),
    .B(_2854_),
    .Y(_2895_));
 sky130_fd_sc_hd__o21bai_2 _3315_ (.A1(_2845_),
    .A2(_2895_),
    .B1_N(_2890_),
    .Y(_2896_));
 sky130_fd_sc_hd__or3b_1 _3316_ (.A(_2845_),
    .B(_2895_),
    .C_N(_2890_),
    .X(_2897_));
 sky130_fd_sc_hd__and2_1 _3317_ (.A(_2896_),
    .B(_2897_),
    .X(_2898_));
 sky130_fd_sc_hd__mux2_1 _3318_ (.A0(\as2650.holding_reg[2] ),
    .A1(net106),
    .S(net199),
    .X(_2899_));
 sky130_fd_sc_hd__o221a_1 _3319_ (.A1(_2765_),
    .A2(_2898_),
    .B1(_2899_),
    .B2(net195),
    .C1(_2894_),
    .X(_2900_));
 sky130_fd_sc_hd__nand2_1 _3320_ (.A(_2660_),
    .B(_2889_),
    .Y(_2901_));
 sky130_fd_sc_hd__o221a_1 _3321_ (.A1(_2851_),
    .A2(_2888_),
    .B1(_2900_),
    .B2(_2658_),
    .C1(_2901_),
    .X(_2902_));
 sky130_fd_sc_hd__mux2_8 _3322_ (.A0(_2890_),
    .A1(_2902_),
    .S(_2769_),
    .X(_2903_));
 sky130_fd_sc_hd__mux2_8 _3323_ (.A0(_2887_),
    .A1(_2903_),
    .S(net71),
    .X(_2904_));
 sky130_fd_sc_hd__a211o_1 _3324_ (.A1(_2787_),
    .A2(_2904_),
    .B1(_2866_),
    .C1(_2788_),
    .X(_2905_));
 sky130_fd_sc_hd__o21a_1 _3325_ (.A1(\as2650.r123[0][2] ),
    .A2(_2789_),
    .B1(_2905_),
    .X(_0009_));
 sky130_fd_sc_hd__or2_1 _3326_ (.A(net247),
    .B(net68),
    .X(_2906_));
 sky130_fd_sc_hd__mux4_2 _3327_ (.A0(\as2650.stack[7][11] ),
    .A1(\as2650.stack[4][11] ),
    .A2(\as2650.stack[5][11] ),
    .A3(\as2650.stack[6][11] ),
    .S0(net215),
    .S1(net217),
    .X(_2907_));
 sky130_fd_sc_hd__o22a_1 _3328_ (.A1(\as2650.stack[3][11] ),
    .A2(net171),
    .B1(net170),
    .B2(\as2650.stack[2][11] ),
    .X(_2908_));
 sky130_fd_sc_hd__o221a_2 _3329_ (.A1(\as2650.stack[1][11] ),
    .A2(net167),
    .B1(net156),
    .B2(\as2650.stack[0][11] ),
    .C1(_2801_),
    .X(_2909_));
 sky130_fd_sc_hd__a22oi_4 _3330_ (.A1(net108),
    .A2(_2907_),
    .B1(_2908_),
    .B2(_2909_),
    .Y(_2910_));
 sky130_fd_sc_hd__nand2_1 _3331_ (.A(net68),
    .B(_2910_),
    .Y(_2911_));
 sky130_fd_sc_hd__a31o_1 _3332_ (.A1(_2809_),
    .A2(_2906_),
    .A3(_2911_),
    .B1(_2788_),
    .X(_2912_));
 sky130_fd_sc_hd__a21oi_4 _3333_ (.A1(_2820_),
    .A2(_2868_),
    .B1(_2869_),
    .Y(_2913_));
 sky130_fd_sc_hd__xnor2_4 _3334_ (.A(net102),
    .B(_2913_),
    .Y(_2914_));
 sky130_fd_sc_hd__or2_1 _3335_ (.A(_2699_),
    .B(_2914_),
    .X(_2915_));
 sky130_fd_sc_hd__o211a_1 _3336_ (.A1(net339),
    .A2(_2700_),
    .B1(_2915_),
    .C1(_2666_),
    .X(_2916_));
 sky130_fd_sc_hd__or2_1 _3337_ (.A(net214),
    .B(\as2650.r123[1][4] ),
    .X(_2917_));
 sky130_fd_sc_hd__nand2b_1 _3338_ (.A_N(\as2650.r123_2[1][4] ),
    .B(net214),
    .Y(_2918_));
 sky130_fd_sc_hd__a32o_1 _3339_ (.A1(_2702_),
    .A2(_2917_),
    .A3(_2918_),
    .B1(net184),
    .B2(_2577_),
    .X(_2919_));
 sky130_fd_sc_hd__mux2_4 _3340_ (.A0(\as2650.r123[2][4] ),
    .A1(\as2650.r123_2[2][4] ),
    .S(net210),
    .X(_2920_));
 sky130_fd_sc_hd__a221o_2 _3341_ (.A1(net245),
    .A2(net178),
    .B1(_2920_),
    .B2(_2583_),
    .C1(_2919_),
    .X(_2921_));
 sky130_fd_sc_hd__a211o_1 _3342_ (.A1(_2665_),
    .A2(net99),
    .B1(_2916_),
    .C1(_2656_),
    .X(_2922_));
 sky130_fd_sc_hd__o211a_1 _3343_ (.A1(_2657_),
    .A2(net105),
    .B1(_2922_),
    .C1(_2695_),
    .X(_2923_));
 sky130_fd_sc_hd__a211o_1 _3344_ (.A1(net246),
    .A2(_2694_),
    .B1(_2923_),
    .C1(_2678_),
    .X(_2924_));
 sky130_fd_sc_hd__nor4_4 _3345_ (.A(net113),
    .B(net112),
    .C(net104),
    .D(net102),
    .Y(_2925_));
 sky130_fd_sc_hd__o31a_1 _3346_ (.A1(net113),
    .A2(net112),
    .A3(net104),
    .B1(net102),
    .X(_2926_));
 sky130_fd_sc_hd__or3_2 _3347_ (.A(_2734_),
    .B(_2925_),
    .C(_2926_),
    .X(_2927_));
 sky130_fd_sc_hd__and3_4 _3348_ (.A(net104),
    .B(_2830_),
    .C(net102),
    .X(_2928_));
 sky130_fd_sc_hd__a21oi_1 _3349_ (.A1(net104),
    .A2(_2830_),
    .B1(net102),
    .Y(_2929_));
 sky130_fd_sc_hd__nor2_2 _3350_ (.A(_2928_),
    .B(_2929_),
    .Y(_2930_));
 sky130_fd_sc_hd__or2_2 _3351_ (.A(_2735_),
    .B(net102),
    .X(_2931_));
 sky130_fd_sc_hd__o211a_2 _3352_ (.A1(_2733_),
    .A2(_2930_),
    .B1(_2931_),
    .C1(_2927_),
    .X(_2932_));
 sky130_fd_sc_hd__o211ai_4 _3353_ (.A1(_2733_),
    .A2(_2930_),
    .B1(_2931_),
    .C1(_2927_),
    .Y(_0284_));
 sky130_fd_sc_hd__a21oi_1 _3354_ (.A1(_2678_),
    .A2(_0284_),
    .B1(_2730_),
    .Y(_0285_));
 sky130_fd_sc_hd__or3_1 _3355_ (.A(_2744_),
    .B(_2925_),
    .C(_2926_),
    .X(_0286_));
 sky130_fd_sc_hd__or2_1 _3356_ (.A(_2745_),
    .B(net102),
    .X(_0287_));
 sky130_fd_sc_hd__o211a_4 _3357_ (.A1(_2743_),
    .A2(_2930_),
    .B1(_0286_),
    .C1(_0287_),
    .X(_0288_));
 sky130_fd_sc_hd__a22o_1 _3358_ (.A1(_2924_),
    .A2(_0285_),
    .B1(_0288_),
    .B2(_2730_),
    .X(_0289_));
 sky130_fd_sc_hd__and2_2 _3359_ (.A(\as2650.holding_reg[3] ),
    .B(net103),
    .X(_0290_));
 sky130_fd_sc_hd__nand2_2 _3360_ (.A(\as2650.holding_reg[3] ),
    .B(net103),
    .Y(_0291_));
 sky130_fd_sc_hd__nor2_4 _3361_ (.A(\as2650.holding_reg[3] ),
    .B(net103),
    .Y(_0292_));
 sky130_fd_sc_hd__nor2_4 _3362_ (.A(_0290_),
    .B(_0292_),
    .Y(_0293_));
 sky130_fd_sc_hd__nand2_1 _3363_ (.A(\as2650.holding_reg[2] ),
    .B(net199),
    .Y(_0294_));
 sky130_fd_sc_hd__nand2_1 _3364_ (.A(net197),
    .B(net106),
    .Y(_0295_));
 sky130_fd_sc_hd__nand2b_1 _3365_ (.A_N(_2899_),
    .B(_2888_),
    .Y(_0296_));
 sky130_fd_sc_hd__a21o_2 _3366_ (.A1(_2896_),
    .A2(_0296_),
    .B1(_0293_),
    .X(_0297_));
 sky130_fd_sc_hd__and3_1 _3367_ (.A(_2896_),
    .B(_0293_),
    .C(_0296_),
    .X(_0298_));
 sky130_fd_sc_hd__or3b_1 _3368_ (.A(_0298_),
    .B(_2765_),
    .C_N(_0297_),
    .X(_0299_));
 sky130_fd_sc_hd__nand2_2 _3369_ (.A(_2888_),
    .B(_2891_),
    .Y(_0300_));
 sky130_fd_sc_hd__and2_1 _3370_ (.A(_2889_),
    .B(_0300_),
    .X(_0301_));
 sky130_fd_sc_hd__xor2_1 _3371_ (.A(_0293_),
    .B(_0301_),
    .X(_0302_));
 sky130_fd_sc_hd__or2_2 _3372_ (.A(\as2650.holding_reg[3] ),
    .B(net198),
    .X(_0303_));
 sky130_fd_sc_hd__o21ai_4 _3373_ (.A1(net199),
    .A2(net103),
    .B1(_0303_),
    .Y(_0304_));
 sky130_fd_sc_hd__mux2_1 _3374_ (.A0(\as2650.holding_reg[3] ),
    .A1(_2874_),
    .S(net199),
    .X(_0305_));
 sky130_fd_sc_hd__a21oi_1 _3375_ (.A1(_2586_),
    .A2(_0305_),
    .B1(_2660_),
    .Y(_0306_));
 sky130_fd_sc_hd__o221a_1 _3376_ (.A1(_2760_),
    .A2(_0302_),
    .B1(_0304_),
    .B2(_2659_),
    .C1(_0306_),
    .X(_0307_));
 sky130_fd_sc_hd__o2bb2a_1 _3377_ (.A1_N(_0299_),
    .A2_N(_0307_),
    .B1(net160),
    .B2(_0290_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_8 _3378_ (.A0(_0293_),
    .A1(_0308_),
    .S(net159),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_8 _3379_ (.A0(_0289_),
    .A1(_0309_),
    .S(net71),
    .X(_0310_));
 sky130_fd_sc_hd__a21o_1 _3380_ (.A1(_2787_),
    .A2(_0310_),
    .B1(_2912_),
    .X(_0311_));
 sky130_fd_sc_hd__o21a_1 _3381_ (.A1(\as2650.r123[0][3] ),
    .A2(_2789_),
    .B1(_0311_),
    .X(_0010_));
 sky130_fd_sc_hd__or2_1 _3382_ (.A(net243),
    .B(net68),
    .X(_0312_));
 sky130_fd_sc_hd__and3_1 _3383_ (.A(net219),
    .B(\as2650.stack[3][12] ),
    .C(net172),
    .X(_0313_));
 sky130_fd_sc_hd__o22a_1 _3384_ (.A1(\as2650.stack[1][12] ),
    .A2(net166),
    .B1(net155),
    .B2(\as2650.stack[0][12] ),
    .X(_0314_));
 sky130_fd_sc_hd__o221a_1 _3385_ (.A1(\as2650.stack[2][12] ),
    .A2(net169),
    .B1(_0313_),
    .B2(net158),
    .C1(_0314_),
    .X(_0315_));
 sky130_fd_sc_hd__mux4_2 _3386_ (.A0(\as2650.stack[7][12] ),
    .A1(\as2650.stack[4][12] ),
    .A2(\as2650.stack[5][12] ),
    .A3(\as2650.stack[6][12] ),
    .S0(net215),
    .S1(net217),
    .X(_0316_));
 sky130_fd_sc_hd__a21oi_4 _3387_ (.A1(net108),
    .A2(_0316_),
    .B1(_0315_),
    .Y(_0317_));
 sky130_fd_sc_hd__nand2_1 _3388_ (.A(net68),
    .B(_0317_),
    .Y(_0318_));
 sky130_fd_sc_hd__a31o_1 _3389_ (.A1(_2809_),
    .A2(_0312_),
    .A3(_0318_),
    .B1(_2788_),
    .X(_0319_));
 sky130_fd_sc_hd__a22o_2 _3390_ (.A1(_2820_),
    .A2(_2925_),
    .B1(_2928_),
    .B2(_2653_),
    .X(_0320_));
 sky130_fd_sc_hd__xor2_4 _3391_ (.A(net98),
    .B(_0320_),
    .X(_0321_));
 sky130_fd_sc_hd__or2_1 _3392_ (.A(_2699_),
    .B(_0321_),
    .X(_0322_));
 sky130_fd_sc_hd__o211a_1 _3393_ (.A1(net335),
    .A2(_2700_),
    .B1(_0322_),
    .C1(_2666_),
    .X(_0323_));
 sky130_fd_sc_hd__nand2b_1 _3394_ (.A_N(\as2650.r123_2[1][5] ),
    .B(net214),
    .Y(_0324_));
 sky130_fd_sc_hd__or2_1 _3395_ (.A(net214),
    .B(\as2650.r123[1][5] ),
    .X(_0325_));
 sky130_fd_sc_hd__a32o_1 _3396_ (.A1(_2702_),
    .A2(_0324_),
    .A3(_0325_),
    .B1(net182),
    .B2(_2577_),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_4 _3397_ (.A0(\as2650.r123[2][5] ),
    .A1(\as2650.r123_2[2][5] ),
    .S(net210),
    .X(_0327_));
 sky130_fd_sc_hd__a221o_4 _3398_ (.A1(net242),
    .A2(net178),
    .B1(_0327_),
    .B2(_2583_),
    .C1(_0326_),
    .X(_0328_));
 sky130_fd_sc_hd__clkinv_4 _3399_ (.A(net97),
    .Y(_0329_));
 sky130_fd_sc_hd__a21o_1 _3400_ (.A1(_2665_),
    .A2(net96),
    .B1(_2656_),
    .X(_0330_));
 sky130_fd_sc_hd__o22a_1 _3401_ (.A1(_2657_),
    .A2(net102),
    .B1(_0323_),
    .B2(_0330_),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _3402_ (.A0(net245),
    .A1(_0331_),
    .S(_2695_),
    .X(_0332_));
 sky130_fd_sc_hd__and2b_1 _3403_ (.A_N(net98),
    .B(_2925_),
    .X(_0333_));
 sky130_fd_sc_hd__xor2_2 _3404_ (.A(net98),
    .B(_2925_),
    .X(_0334_));
 sky130_fd_sc_hd__xnor2_4 _3405_ (.A(net98),
    .B(_2928_),
    .Y(_0335_));
 sky130_fd_sc_hd__nand2_1 _3406_ (.A(_2732_),
    .B(_0335_),
    .Y(_0336_));
 sky130_fd_sc_hd__o221a_4 _3407_ (.A1(_2735_),
    .A2(net98),
    .B1(_0334_),
    .B2(_2734_),
    .C1(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _3408_ (.A0(_0332_),
    .A1(_0337_),
    .S(_2739_),
    .X(_0338_));
 sky130_fd_sc_hd__o22a_1 _3409_ (.A1(_2745_),
    .A2(net98),
    .B1(_0334_),
    .B2(_2744_),
    .X(_0339_));
 sky130_fd_sc_hd__a21boi_4 _3410_ (.A1(_2742_),
    .A2(_0335_),
    .B1_N(_0339_),
    .Y(_0340_));
 sky130_fd_sc_hd__a21bo_4 _3411_ (.A1(_2742_),
    .A2(_0335_),
    .B1_N(_0339_),
    .X(_0341_));
 sky130_fd_sc_hd__mux2_2 _3412_ (.A0(_0338_),
    .A1(_0340_),
    .S(_2730_),
    .X(_0342_));
 sky130_fd_sc_hd__and2_2 _3413_ (.A(\as2650.holding_reg[4] ),
    .B(net101),
    .X(_0343_));
 sky130_fd_sc_hd__nor2_1 _3414_ (.A(\as2650.holding_reg[4] ),
    .B(net101),
    .Y(_0344_));
 sky130_fd_sc_hd__or2_4 _3415_ (.A(_0343_),
    .B(_0344_),
    .X(_0345_));
 sky130_fd_sc_hd__or2_2 _3416_ (.A(_0290_),
    .B(_0304_),
    .X(_0346_));
 sky130_fd_sc_hd__a21boi_4 _3417_ (.A1(_0297_),
    .A2(_0346_),
    .B1_N(_0345_),
    .Y(_0347_));
 sky130_fd_sc_hd__and3b_1 _3418_ (.A_N(_0345_),
    .B(_0346_),
    .C(_0297_),
    .X(_0348_));
 sky130_fd_sc_hd__nor3_1 _3419_ (.A(_2765_),
    .B(_0347_),
    .C(_0348_),
    .Y(_0349_));
 sky130_fd_sc_hd__o211a_1 _3420_ (.A1(_0292_),
    .A2(_0301_),
    .B1(_0345_),
    .C1(_0291_),
    .X(_0350_));
 sky130_fd_sc_hd__a311oi_4 _3421_ (.A1(_2889_),
    .A2(_0291_),
    .A3(_0300_),
    .B1(_0345_),
    .C1(_0292_),
    .Y(_0351_));
 sky130_fd_sc_hd__or3_1 _3422_ (.A(_2760_),
    .B(_0350_),
    .C(_0351_),
    .X(_0352_));
 sky130_fd_sc_hd__or2_2 _3423_ (.A(\as2650.holding_reg[4] ),
    .B(net198),
    .X(_0353_));
 sky130_fd_sc_hd__o21ai_4 _3424_ (.A1(net199),
    .A2(net101),
    .B1(_0353_),
    .Y(_0354_));
 sky130_fd_sc_hd__mux2_1 _3425_ (.A0(\as2650.holding_reg[4] ),
    .A1(net101),
    .S(net199),
    .X(_0355_));
 sky130_fd_sc_hd__inv_2 _3426_ (.A(_0355_),
    .Y(_0356_));
 sky130_fd_sc_hd__o221a_1 _3427_ (.A1(_2659_),
    .A2(_0354_),
    .B1(_0356_),
    .B2(net195),
    .C1(net160),
    .X(_0357_));
 sky130_fd_sc_hd__and3b_1 _3428_ (.A_N(_0349_),
    .B(_0352_),
    .C(_0357_),
    .X(_0358_));
 sky130_fd_sc_hd__o21ai_1 _3429_ (.A1(net160),
    .A2(_0343_),
    .B1(net159),
    .Y(_0359_));
 sky130_fd_sc_hd__o22a_4 _3430_ (.A1(net159),
    .A2(_0345_),
    .B1(_0358_),
    .B2(_0359_),
    .X(_0360_));
 sky130_fd_sc_hd__inv_2 _3431_ (.A(_0360_),
    .Y(_0361_));
 sky130_fd_sc_hd__mux2_8 _3432_ (.A0(_0342_),
    .A1(_0361_),
    .S(net71),
    .X(_0362_));
 sky130_fd_sc_hd__a21o_1 _3433_ (.A1(_2787_),
    .A2(_0362_),
    .B1(_0319_),
    .X(_0363_));
 sky130_fd_sc_hd__o21a_1 _3434_ (.A1(\as2650.r123[0][4] ),
    .A2(_2789_),
    .B1(_0363_),
    .X(_0011_));
 sky130_fd_sc_hd__or2_1 _3435_ (.A(net242),
    .B(net68),
    .X(_0364_));
 sky130_fd_sc_hd__o22a_1 _3436_ (.A1(\as2650.stack[7][13] ),
    .A2(_2791_),
    .B1(net169),
    .B2(\as2650.stack[6][13] ),
    .X(_0365_));
 sky130_fd_sc_hd__o22a_1 _3437_ (.A1(\as2650.stack[5][13] ),
    .A2(net166),
    .B1(net155),
    .B2(\as2650.stack[4][13] ),
    .X(_0366_));
 sky130_fd_sc_hd__and3_1 _3438_ (.A(net108),
    .B(_0365_),
    .C(_0366_),
    .X(_0367_));
 sky130_fd_sc_hd__o22a_1 _3439_ (.A1(\as2650.stack[1][13] ),
    .A2(net166),
    .B1(net155),
    .B2(\as2650.stack[0][13] ),
    .X(_0368_));
 sky130_fd_sc_hd__o221a_2 _3440_ (.A1(\as2650.stack[3][13] ),
    .A2(net171),
    .B1(net169),
    .B2(\as2650.stack[2][13] ),
    .C1(_0368_),
    .X(_0369_));
 sky130_fd_sc_hd__a21oi_4 _3441_ (.A1(_2801_),
    .A2(_0369_),
    .B1(_0367_),
    .Y(_0370_));
 sky130_fd_sc_hd__nand2_1 _3442_ (.A(net68),
    .B(_0370_),
    .Y(_0371_));
 sky130_fd_sc_hd__a31o_1 _3443_ (.A1(_2809_),
    .A2(_0364_),
    .A3(_0371_),
    .B1(_2788_),
    .X(_0372_));
 sky130_fd_sc_hd__nor2_1 _3444_ (.A(net98),
    .B(net96),
    .Y(_0373_));
 sky130_fd_sc_hd__and2_4 _3445_ (.A(_2925_),
    .B(_0373_),
    .X(_0374_));
 sky130_fd_sc_hd__inv_2 _3446_ (.A(_0374_),
    .Y(_0375_));
 sky130_fd_sc_hd__and3_1 _3447_ (.A(_2820_),
    .B(_2925_),
    .C(_0373_),
    .X(_0376_));
 sky130_fd_sc_hd__and3_4 _3448_ (.A(net98),
    .B(_2928_),
    .C(net96),
    .X(_0377_));
 sky130_fd_sc_hd__and2_1 _3449_ (.A(_2653_),
    .B(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__a21oi_2 _3450_ (.A1(net98),
    .A2(_2928_),
    .B1(net96),
    .Y(_0379_));
 sky130_fd_sc_hd__a221o_1 _3451_ (.A1(_2654_),
    .A2(_0329_),
    .B1(_0333_),
    .B2(_2820_),
    .C1(_0379_),
    .X(_0380_));
 sky130_fd_sc_hd__o21ba_2 _3452_ (.A1(_0378_),
    .A2(_0380_),
    .B1_N(_0376_),
    .X(_0381_));
 sky130_fd_sc_hd__mux2_4 _3453_ (.A0(\as2650.r123[2][6] ),
    .A1(\as2650.r123_2[2][6] ),
    .S(net210),
    .X(_0382_));
 sky130_fd_sc_hd__mux4_1 _3454_ (.A0(\as2650.r123[1][6] ),
    .A1(\as2650.r123[0][6] ),
    .A2(\as2650.r123_2[1][6] ),
    .A3(\as2650.r123_2[0][6] ),
    .S0(net307),
    .S1(net210),
    .X(_0383_));
 sky130_fd_sc_hd__a22o_1 _3455_ (.A1(_2583_),
    .A2(_0382_),
    .B1(_0383_),
    .B2(_2704_),
    .X(_0384_));
 sky130_fd_sc_hd__a21o_2 _3456_ (.A1(net239),
    .A2(net178),
    .B1(_0384_),
    .X(_0385_));
 sky130_fd_sc_hd__nand2_1 _3457_ (.A(_2700_),
    .B(_0381_),
    .Y(_0386_));
 sky130_fd_sc_hd__o211a_1 _3458_ (.A1(net332),
    .A2(_2700_),
    .B1(_0386_),
    .C1(_2666_),
    .X(_0387_));
 sky130_fd_sc_hd__a211o_1 _3459_ (.A1(_2665_),
    .A2(net94),
    .B1(_0387_),
    .C1(_2656_),
    .X(_0388_));
 sky130_fd_sc_hd__o21a_1 _3460_ (.A1(_2657_),
    .A2(net99),
    .B1(_2695_),
    .X(_0389_));
 sky130_fd_sc_hd__a22o_1 _3461_ (.A1(net240),
    .A2(_2694_),
    .B1(_0388_),
    .B2(_0389_),
    .X(_0390_));
 sky130_fd_sc_hd__o21ai_1 _3462_ (.A1(_0377_),
    .A2(_0379_),
    .B1(_2732_),
    .Y(_0391_));
 sky130_fd_sc_hd__nor2_1 _3463_ (.A(_0329_),
    .B(_0333_),
    .Y(_0392_));
 sky130_fd_sc_hd__or2_2 _3464_ (.A(_0374_),
    .B(_0392_),
    .X(_0393_));
 sky130_fd_sc_hd__o221a_4 _3465_ (.A1(_2735_),
    .A2(net96),
    .B1(_0393_),
    .B2(_2734_),
    .C1(_0391_),
    .X(_0394_));
 sky130_fd_sc_hd__o21ai_1 _3466_ (.A1(_0377_),
    .A2(_0379_),
    .B1(_2742_),
    .Y(_0395_));
 sky130_fd_sc_hd__o221a_4 _3467_ (.A1(_2745_),
    .A2(net96),
    .B1(_0393_),
    .B2(_2744_),
    .C1(_0395_),
    .X(_0396_));
 sky130_fd_sc_hd__mux2_1 _3468_ (.A0(_0390_),
    .A1(_0394_),
    .S(_2739_),
    .X(_0397_));
 sky130_fd_sc_hd__mux2_1 _3469_ (.A0(_0396_),
    .A1(_0397_),
    .S(_2731_),
    .X(_0398_));
 sky130_fd_sc_hd__nor2_2 _3470_ (.A(_2555_),
    .B(_0329_),
    .Y(_0399_));
 sky130_fd_sc_hd__nor2_1 _3471_ (.A(\as2650.holding_reg[5] ),
    .B(net97),
    .Y(_0400_));
 sky130_fd_sc_hd__or2_4 _3472_ (.A(_0399_),
    .B(_0400_),
    .X(_0401_));
 sky130_fd_sc_hd__nor2_1 _3473_ (.A(_0343_),
    .B(_0354_),
    .Y(_0402_));
 sky130_fd_sc_hd__o21ai_2 _3474_ (.A1(_0347_),
    .A2(_0402_),
    .B1(_0401_),
    .Y(_0403_));
 sky130_fd_sc_hd__or3_1 _3475_ (.A(_0347_),
    .B(_0401_),
    .C(_0402_),
    .X(_0404_));
 sky130_fd_sc_hd__or3b_1 _3476_ (.A(_0343_),
    .B(_0351_),
    .C_N(_0401_),
    .X(_0405_));
 sky130_fd_sc_hd__o21ba_1 _3477_ (.A1(_0343_),
    .A2(_0351_),
    .B1_N(_0401_),
    .X(_0406_));
 sky130_fd_sc_hd__and3b_1 _3478_ (.A_N(_0406_),
    .B(_2759_),
    .C(_0405_),
    .X(_0407_));
 sky130_fd_sc_hd__mux2_2 _3479_ (.A0(_2555_),
    .A1(_0329_),
    .S(net198),
    .X(_0408_));
 sky130_fd_sc_hd__mux2_1 _3480_ (.A0(\as2650.holding_reg[5] ),
    .A1(net97),
    .S(net200),
    .X(_0409_));
 sky130_fd_sc_hd__a21oi_1 _3481_ (.A1(\as2650.ins_reg[5] ),
    .A2(_0408_),
    .B1(_2659_),
    .Y(_0410_));
 sky130_fd_sc_hd__a31o_1 _3482_ (.A1(_2764_),
    .A2(_0403_),
    .A3(_0404_),
    .B1(_0410_),
    .X(_0411_));
 sky130_fd_sc_hd__a211o_1 _3483_ (.A1(_2586_),
    .A2(_0409_),
    .B1(_0411_),
    .C1(_0407_),
    .X(_0412_));
 sky130_fd_sc_hd__o21a_1 _3484_ (.A1(net160),
    .A2(_0399_),
    .B1(_2769_),
    .X(_0413_));
 sky130_fd_sc_hd__a2bb2o_4 _3485_ (.A1_N(net159),
    .A2_N(_0401_),
    .B1(_0412_),
    .B2(_0413_),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_8 _3486_ (.A0(_0398_),
    .A1(_0414_),
    .S(_2749_),
    .X(_0415_));
 sky130_fd_sc_hd__a21o_1 _3487_ (.A1(_2787_),
    .A2(_0415_),
    .B1(_0372_),
    .X(_0416_));
 sky130_fd_sc_hd__o21a_1 _3488_ (.A1(\as2650.r123[0][5] ),
    .A2(_2789_),
    .B1(_0416_),
    .X(_0012_));
 sky130_fd_sc_hd__or2_1 _3489_ (.A(net237),
    .B(net68),
    .X(_0417_));
 sky130_fd_sc_hd__and3_1 _3490_ (.A(net219),
    .B(\as2650.stack[3][14] ),
    .C(net172),
    .X(_0418_));
 sky130_fd_sc_hd__o22a_1 _3491_ (.A1(\as2650.stack[1][14] ),
    .A2(net166),
    .B1(net155),
    .B2(\as2650.stack[0][14] ),
    .X(_0419_));
 sky130_fd_sc_hd__o221a_1 _3492_ (.A1(\as2650.stack[2][14] ),
    .A2(net169),
    .B1(_0418_),
    .B2(_2792_),
    .C1(_0419_),
    .X(_0420_));
 sky130_fd_sc_hd__mux4_1 _3493_ (.A0(\as2650.stack[7][14] ),
    .A1(\as2650.stack[4][14] ),
    .A2(\as2650.stack[5][14] ),
    .A3(\as2650.stack[6][14] ),
    .S0(net215),
    .S1(net217),
    .X(_0421_));
 sky130_fd_sc_hd__a21o_2 _3494_ (.A1(net108),
    .A2(_0421_),
    .B1(_0420_),
    .X(_0422_));
 sky130_fd_sc_hd__or2_1 _3495_ (.A(net67),
    .B(_0422_),
    .X(_0423_));
 sky130_fd_sc_hd__a31o_1 _3496_ (.A1(_2809_),
    .A2(_0417_),
    .A3(_0423_),
    .B1(_2788_),
    .X(_0424_));
 sky130_fd_sc_hd__nor2_2 _3497_ (.A(_0376_),
    .B(_0378_),
    .Y(_0425_));
 sky130_fd_sc_hd__xnor2_4 _3498_ (.A(net93),
    .B(_0425_),
    .Y(_0426_));
 sky130_fd_sc_hd__a221o_1 _3499_ (.A1(net331),
    .A2(_2699_),
    .B1(_2711_),
    .B2(_0426_),
    .C1(_2665_),
    .X(_0427_));
 sky130_fd_sc_hd__o211a_1 _3500_ (.A1(_2666_),
    .A2(net109),
    .B1(_0427_),
    .C1(_2657_),
    .X(_0428_));
 sky130_fd_sc_hd__a211o_1 _3501_ (.A1(_2656_),
    .A2(net96),
    .B1(_0428_),
    .C1(_2694_),
    .X(_0429_));
 sky130_fd_sc_hd__o211a_1 _3502_ (.A1(net238),
    .A2(_2695_),
    .B1(_2737_),
    .C1(_0429_),
    .X(_0430_));
 sky130_fd_sc_hd__nor2_4 _3503_ (.A(_0375_),
    .B(net93),
    .Y(_0431_));
 sky130_fd_sc_hd__xor2_1 _3504_ (.A(_0374_),
    .B(net93),
    .X(_0432_));
 sky130_fd_sc_hd__nand2_1 _3505_ (.A(_0377_),
    .B(net93),
    .Y(_0433_));
 sky130_fd_sc_hd__xor2_2 _3506_ (.A(_0377_),
    .B(net93),
    .X(_0434_));
 sky130_fd_sc_hd__o22a_1 _3507_ (.A1(_2734_),
    .A2(_0432_),
    .B1(_0434_),
    .B2(_2733_),
    .X(_0435_));
 sky130_fd_sc_hd__o21a_4 _3508_ (.A1(_2735_),
    .A2(net93),
    .B1(_0435_),
    .X(_0436_));
 sky130_fd_sc_hd__a211o_1 _3509_ (.A1(_2678_),
    .A2(_0436_),
    .B1(_0430_),
    .C1(_2730_),
    .X(_0437_));
 sky130_fd_sc_hd__or2_1 _3510_ (.A(_2744_),
    .B(_0432_),
    .X(_0438_));
 sky130_fd_sc_hd__o221a_4 _3511_ (.A1(_2745_),
    .A2(net93),
    .B1(_0434_),
    .B2(_2743_),
    .C1(_0438_),
    .X(_0439_));
 sky130_fd_sc_hd__o211a_1 _3512_ (.A1(_2731_),
    .A2(_0439_),
    .B1(_0437_),
    .C1(_2747_),
    .X(_0440_));
 sky130_fd_sc_hd__and2_2 _3513_ (.A(\as2650.holding_reg[6] ),
    .B(net95),
    .X(_0441_));
 sky130_fd_sc_hd__nor2_1 _3514_ (.A(\as2650.holding_reg[6] ),
    .B(net95),
    .Y(_0442_));
 sky130_fd_sc_hd__nor2_4 _3515_ (.A(_0441_),
    .B(_0442_),
    .Y(_0443_));
 sky130_fd_sc_hd__inv_2 _3516_ (.A(_0443_),
    .Y(_0444_));
 sky130_fd_sc_hd__o21a_1 _3517_ (.A1(_0399_),
    .A2(_0406_),
    .B1(_0443_),
    .X(_0445_));
 sky130_fd_sc_hd__nor2_1 _3518_ (.A(_2760_),
    .B(_0445_),
    .Y(_0446_));
 sky130_fd_sc_hd__o31a_1 _3519_ (.A1(_0399_),
    .A2(_0406_),
    .A3(_0443_),
    .B1(_0446_),
    .X(_0447_));
 sky130_fd_sc_hd__or2_1 _3520_ (.A(_0399_),
    .B(_0408_),
    .X(_0448_));
 sky130_fd_sc_hd__a21oi_1 _3521_ (.A1(_0403_),
    .A2(_0448_),
    .B1(_0443_),
    .Y(_0449_));
 sky130_fd_sc_hd__a31o_1 _3522_ (.A1(_0403_),
    .A2(_0443_),
    .A3(_0448_),
    .B1(_2765_),
    .X(_0450_));
 sky130_fd_sc_hd__or2_2 _3523_ (.A(\as2650.holding_reg[6] ),
    .B(net198),
    .X(_0451_));
 sky130_fd_sc_hd__o21ai_4 _3524_ (.A1(net200),
    .A2(net95),
    .B1(_0451_),
    .Y(_0452_));
 sky130_fd_sc_hd__mux2_1 _3525_ (.A0(\as2650.holding_reg[6] ),
    .A1(net95),
    .S(net200),
    .X(_0453_));
 sky130_fd_sc_hd__inv_2 _3526_ (.A(_0453_),
    .Y(_0454_));
 sky130_fd_sc_hd__o221a_1 _3527_ (.A1(_2659_),
    .A2(_0452_),
    .B1(_0454_),
    .B2(net195),
    .C1(net160),
    .X(_0455_));
 sky130_fd_sc_hd__o21ai_1 _3528_ (.A1(_0449_),
    .A2(_0450_),
    .B1(_0455_),
    .Y(_0456_));
 sky130_fd_sc_hd__o22a_1 _3529_ (.A1(net160),
    .A2(_0441_),
    .B1(_0447_),
    .B2(_0456_),
    .X(_0457_));
 sky130_fd_sc_hd__mux2_8 _3530_ (.A0(_0443_),
    .A1(_0457_),
    .S(net159),
    .X(_0458_));
 sky130_fd_sc_hd__a21o_4 _3531_ (.A1(_2749_),
    .A2(_0458_),
    .B1(_0440_),
    .X(_0459_));
 sky130_fd_sc_hd__a21o_1 _3532_ (.A1(_2787_),
    .A2(_0459_),
    .B1(_0424_),
    .X(_0460_));
 sky130_fd_sc_hd__o21a_1 _3533_ (.A1(\as2650.r123[0][6] ),
    .A2(_2789_),
    .B1(_0460_),
    .X(_0013_));
 sky130_fd_sc_hd__a31o_1 _3534_ (.A1(net234),
    .A2(net67),
    .A3(_2809_),
    .B1(_2788_),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_4 _3535_ (.A0(_0376_),
    .A1(_0378_),
    .S(net93),
    .X(_0462_));
 sky130_fd_sc_hd__xor2_4 _3536_ (.A(net110),
    .B(_0462_),
    .X(_0463_));
 sky130_fd_sc_hd__nand2_1 _3537_ (.A(net312),
    .B(_2699_),
    .Y(_0464_));
 sky130_fd_sc_hd__o211a_1 _3538_ (.A1(_2699_),
    .A2(_0463_),
    .B1(_0464_),
    .C1(_2666_),
    .X(_0465_));
 sky130_fd_sc_hd__o21a_1 _3539_ (.A1(\as2650.psl[3] ),
    .A2(net114),
    .B1(_2720_),
    .X(_0466_));
 sky130_fd_sc_hd__o21ai_1 _3540_ (.A1(\as2650.psl[3] ),
    .A2(net114),
    .B1(_2720_),
    .Y(_0467_));
 sky130_fd_sc_hd__a21o_1 _3541_ (.A1(_2665_),
    .A2(_0466_),
    .B1(_2656_),
    .X(_0468_));
 sky130_fd_sc_hd__o22a_1 _3542_ (.A1(_2657_),
    .A2(net94),
    .B1(_0465_),
    .B2(_0468_),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _3543_ (.A0(net235),
    .A1(_0469_),
    .S(_2695_),
    .X(_0470_));
 sky130_fd_sc_hd__xnor2_1 _3544_ (.A(net110),
    .B(_0433_),
    .Y(_0471_));
 sky130_fd_sc_hd__or2_1 _3545_ (.A(_2733_),
    .B(_0471_),
    .X(_0472_));
 sky130_fd_sc_hd__xor2_4 _3546_ (.A(net110),
    .B(_0431_),
    .X(_0473_));
 sky130_fd_sc_hd__o221a_4 _3547_ (.A1(net110),
    .A2(_2735_),
    .B1(_0473_),
    .B2(_2734_),
    .C1(_0472_),
    .X(_0474_));
 sky130_fd_sc_hd__mux2_1 _3548_ (.A0(_0470_),
    .A1(_0474_),
    .S(_2739_),
    .X(_0475_));
 sky130_fd_sc_hd__or2_1 _3549_ (.A(_2743_),
    .B(_0471_),
    .X(_0476_));
 sky130_fd_sc_hd__o221a_4 _3550_ (.A1(net110),
    .A2(_2745_),
    .B1(_0473_),
    .B2(_2744_),
    .C1(_0476_),
    .X(_0477_));
 sky130_fd_sc_hd__mux2_1 _3551_ (.A0(_0475_),
    .A1(_0477_),
    .S(_2730_),
    .X(_0478_));
 sky130_fd_sc_hd__nand2_1 _3552_ (.A(\as2650.holding_reg[7] ),
    .B(net109),
    .Y(_0479_));
 sky130_fd_sc_hd__or2_2 _3553_ (.A(\as2650.holding_reg[7] ),
    .B(net109),
    .X(_0480_));
 sky130_fd_sc_hd__and2_2 _3554_ (.A(_0479_),
    .B(_0480_),
    .X(_0481_));
 sky130_fd_sc_hd__nand2_2 _3555_ (.A(_0479_),
    .B(_0480_),
    .Y(_0482_));
 sky130_fd_sc_hd__nor2_1 _3556_ (.A(_0441_),
    .B(_0452_),
    .Y(_0483_));
 sky130_fd_sc_hd__nor2_1 _3557_ (.A(_0449_),
    .B(_0483_),
    .Y(_0484_));
 sky130_fd_sc_hd__xnor2_1 _3558_ (.A(_0481_),
    .B(_0484_),
    .Y(_0485_));
 sky130_fd_sc_hd__nor2_1 _3559_ (.A(_0441_),
    .B(_0445_),
    .Y(_0486_));
 sky130_fd_sc_hd__xnor2_1 _3560_ (.A(_0482_),
    .B(_0486_),
    .Y(_0487_));
 sky130_fd_sc_hd__mux2_1 _3561_ (.A0(\as2650.holding_reg[7] ),
    .A1(net109),
    .S(net200),
    .X(_0488_));
 sky130_fd_sc_hd__inv_2 _3562_ (.A(_0488_),
    .Y(_0489_));
 sky130_fd_sc_hd__o221a_1 _3563_ (.A1(_2760_),
    .A2(_0487_),
    .B1(_0489_),
    .B2(_2585_),
    .C1(_2851_),
    .X(_0490_));
 sky130_fd_sc_hd__o21ai_1 _3564_ (.A1(_2765_),
    .A2(_0485_),
    .B1(_0490_),
    .Y(_0491_));
 sky130_fd_sc_hd__o211a_1 _3565_ (.A1(_2659_),
    .A2(_0480_),
    .B1(_0491_),
    .C1(net160),
    .X(_0492_));
 sky130_fd_sc_hd__o21ai_1 _3566_ (.A1(net160),
    .A2(_0479_),
    .B1(net159),
    .Y(_0493_));
 sky130_fd_sc_hd__o22a_4 _3567_ (.A1(net159),
    .A2(_0481_),
    .B1(_0492_),
    .B2(_0493_),
    .X(_0494_));
 sky130_fd_sc_hd__mux2_4 _3568_ (.A0(_0478_),
    .A1(_0494_),
    .S(_2749_),
    .X(_0495_));
 sky130_fd_sc_hd__a21o_1 _3569_ (.A1(_2787_),
    .A2(_0495_),
    .B1(_0461_),
    .X(_0496_));
 sky130_fd_sc_hd__o21a_1 _3570_ (.A1(\as2650.r123[0][7] ),
    .A2(_2789_),
    .B1(_0496_),
    .X(_0014_));
 sky130_fd_sc_hd__or2_4 _3571_ (.A(_2529_),
    .B(net157),
    .X(_0497_));
 sky130_fd_sc_hd__or2_4 _3572_ (.A(net49),
    .B(_0497_),
    .X(_0498_));
 sky130_fd_sc_hd__or2_1 _3573_ (.A(_2631_),
    .B(_0497_),
    .X(_0499_));
 sky130_fd_sc_hd__and2_4 _3574_ (.A(_0498_),
    .B(_0499_),
    .X(_0500_));
 sky130_fd_sc_hd__mux2_1 _3575_ (.A0(_2625_),
    .A1(\as2650.stack[5][8] ),
    .S(_0500_),
    .X(_0015_));
 sky130_fd_sc_hd__mux2_1 _3576_ (.A0(_2633_),
    .A1(\as2650.stack[5][9] ),
    .S(_0500_),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_1 _3577_ (.A0(_2635_),
    .A1(\as2650.stack[5][10] ),
    .S(_0500_),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _3578_ (.A0(_2637_),
    .A1(\as2650.stack[5][11] ),
    .S(_0500_),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _3579_ (.A0(_2639_),
    .A1(\as2650.stack[5][12] ),
    .S(_0500_),
    .X(_0019_));
 sky130_fd_sc_hd__mux2_1 _3580_ (.A0(_2641_),
    .A1(\as2650.stack[5][13] ),
    .S(_0500_),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_1 _3581_ (.A0(_2643_),
    .A1(\as2650.stack[5][14] ),
    .S(_0500_),
    .X(_0021_));
 sky130_fd_sc_hd__nor2_8 _3582_ (.A(net47),
    .B(_0497_),
    .Y(_0501_));
 sky130_fd_sc_hd__mux2_1 _3583_ (.A0(net286),
    .A1(\as2650.stack[5][0] ),
    .S(_0499_),
    .X(_0502_));
 sky130_fd_sc_hd__mux2_1 _3584_ (.A0(net259),
    .A1(_0502_),
    .S(_2582_),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_1 _3585_ (.A0(\as2650.stack[5][1] ),
    .A1(net282),
    .S(_0501_),
    .X(_0503_));
 sky130_fd_sc_hd__mux2_1 _3586_ (.A0(net254),
    .A1(_0503_),
    .S(_2582_),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_1 _3587_ (.A0(\as2650.stack[5][2] ),
    .A1(net280),
    .S(_0501_),
    .X(_0504_));
 sky130_fd_sc_hd__mux2_1 _3588_ (.A0(net250),
    .A1(_0504_),
    .S(_2582_),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_1 _3589_ (.A0(\as2650.stack[5][3] ),
    .A1(net277),
    .S(_0501_),
    .X(_0505_));
 sky130_fd_sc_hd__mux2_1 _3590_ (.A0(net246),
    .A1(_0505_),
    .S(_2582_),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_1 _3591_ (.A0(\as2650.stack[5][4] ),
    .A1(net276),
    .S(_0501_),
    .X(_0506_));
 sky130_fd_sc_hd__mux2_1 _3592_ (.A0(net243),
    .A1(_0506_),
    .S(_2582_),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_1 _3593_ (.A0(\as2650.stack[5][5] ),
    .A1(net273),
    .S(_0501_),
    .X(_0507_));
 sky130_fd_sc_hd__mux2_1 _3594_ (.A0(net240),
    .A1(_0507_),
    .S(_2582_),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _3595_ (.A0(\as2650.stack[5][6] ),
    .A1(net271),
    .S(_0501_),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_1 _3596_ (.A0(net237),
    .A1(_0508_),
    .S(_2582_),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _3597_ (.A0(\as2650.stack[5][7] ),
    .A1(net269),
    .S(_0501_),
    .X(_0509_));
 sky130_fd_sc_hd__mux2_1 _3598_ (.A0(net232),
    .A1(_0509_),
    .S(_2582_),
    .X(_0029_));
 sky130_fd_sc_hd__or2_4 _3599_ (.A(net49),
    .B(_2793_),
    .X(_0510_));
 sky130_fd_sc_hd__or2_1 _3600_ (.A(_2631_),
    .B(_2793_),
    .X(_0511_));
 sky130_fd_sc_hd__and2_4 _3601_ (.A(_0510_),
    .B(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__mux2_1 _3602_ (.A0(_2625_),
    .A1(\as2650.stack[4][8] ),
    .S(_0512_),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _3603_ (.A0(_2633_),
    .A1(\as2650.stack[4][9] ),
    .S(_0512_),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _3604_ (.A0(_2635_),
    .A1(\as2650.stack[4][10] ),
    .S(_0512_),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _3605_ (.A0(_2637_),
    .A1(\as2650.stack[4][11] ),
    .S(_0512_),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _3606_ (.A0(_2639_),
    .A1(\as2650.stack[4][12] ),
    .S(_0512_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _3607_ (.A0(_2641_),
    .A1(\as2650.stack[4][13] ),
    .S(_0512_),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _3608_ (.A0(_2643_),
    .A1(\as2650.stack[4][14] ),
    .S(_0512_),
    .X(_0036_));
 sky130_fd_sc_hd__nand2_1 _3609_ (.A(net213),
    .B(_2560_),
    .Y(_0513_));
 sky130_fd_sc_hd__or2_4 _3610_ (.A(net145),
    .B(_0513_),
    .X(_0514_));
 sky130_fd_sc_hd__or2_4 _3611_ (.A(net177),
    .B(_0514_),
    .X(_0515_));
 sky130_fd_sc_hd__nor2_4 _3612_ (.A(_2664_),
    .B(_0515_),
    .Y(_0516_));
 sky130_fd_sc_hd__or2_4 _3613_ (.A(_2664_),
    .B(_0515_),
    .X(_0517_));
 sky130_fd_sc_hd__nor2_4 _3614_ (.A(_2693_),
    .B(_0515_),
    .Y(_0518_));
 sky130_fd_sc_hd__or2_4 _3615_ (.A(_2693_),
    .B(_0515_),
    .X(_0519_));
 sky130_fd_sc_hd__nand2_2 _3616_ (.A(net213),
    .B(_2645_),
    .Y(_0520_));
 sky130_fd_sc_hd__nor3_4 _3617_ (.A(_2673_),
    .B(_2677_),
    .C(net154),
    .Y(_0521_));
 sky130_fd_sc_hd__or3_4 _3618_ (.A(_2673_),
    .B(_2677_),
    .C(net154),
    .X(_0522_));
 sky130_fd_sc_hd__nor2_4 _3619_ (.A(_2655_),
    .B(_0515_),
    .Y(_0523_));
 sky130_fd_sc_hd__or2_4 _3620_ (.A(_2655_),
    .B(_0515_),
    .X(_0524_));
 sky130_fd_sc_hd__or4_4 _3621_ (.A(_2525_),
    .B(_2561_),
    .C(_2696_),
    .D(_2698_),
    .X(_0525_));
 sky130_fd_sc_hd__o211a_1 _3622_ (.A1(_2691_),
    .A2(net154),
    .B1(_0524_),
    .C1(_0525_),
    .X(_0526_));
 sky130_fd_sc_hd__and4_4 _3623_ (.A(_0517_),
    .B(_0519_),
    .C(_0522_),
    .D(_0526_),
    .X(_0527_));
 sky130_fd_sc_hd__nor2_1 _3624_ (.A(net305),
    .B(_0527_),
    .Y(_0528_));
 sky130_fd_sc_hd__nor2_4 _3625_ (.A(_2683_),
    .B(net154),
    .Y(_0529_));
 sky130_fd_sc_hd__or2_2 _3626_ (.A(_2683_),
    .B(_0520_),
    .X(_0530_));
 sky130_fd_sc_hd__or2_1 _3627_ (.A(_2710_),
    .B(_0520_),
    .X(_0531_));
 sky130_fd_sc_hd__a221o_1 _3628_ (.A1(net350),
    .A2(_0529_),
    .B1(_0531_),
    .B2(_2709_),
    .C1(_0516_),
    .X(_0532_));
 sky130_fd_sc_hd__o211a_1 _3629_ (.A1(_2718_),
    .A2(_0517_),
    .B1(_0524_),
    .C1(_0532_),
    .X(_0533_));
 sky130_fd_sc_hd__a21o_1 _3630_ (.A1(_2727_),
    .A2(_0523_),
    .B1(_0518_),
    .X(_0534_));
 sky130_fd_sc_hd__o22a_1 _3631_ (.A1(net262),
    .A2(_0519_),
    .B1(_0533_),
    .B2(_0534_),
    .X(_0535_));
 sky130_fd_sc_hd__or3_1 _3632_ (.A(_2673_),
    .B(_2677_),
    .C(net154),
    .X(_0536_));
 sky130_fd_sc_hd__or3_1 _3633_ (.A(_2673_),
    .B(_2677_),
    .C(net154),
    .X(_0537_));
 sky130_fd_sc_hd__nor2_2 _3634_ (.A(_2688_),
    .B(net154),
    .Y(_0538_));
 sky130_fd_sc_hd__or2_4 _3635_ (.A(_2688_),
    .B(net154),
    .X(_0539_));
 sky130_fd_sc_hd__or2_1 _3636_ (.A(_2736_),
    .B(_0522_),
    .X(_0540_));
 sky130_fd_sc_hd__nor2_2 _3637_ (.A(_2741_),
    .B(net154),
    .Y(_0541_));
 sky130_fd_sc_hd__o211a_1 _3638_ (.A1(_0521_),
    .A2(_0535_),
    .B1(_0539_),
    .C1(_0540_),
    .X(_0542_));
 sky130_fd_sc_hd__or3_4 _3639_ (.A(_2696_),
    .B(_2698_),
    .C(_0513_),
    .X(_0543_));
 sky130_fd_sc_hd__inv_2 _3640_ (.A(_0543_),
    .Y(_0544_));
 sky130_fd_sc_hd__or4_1 _3641_ (.A(_2525_),
    .B(net126),
    .C(_2674_),
    .D(_2698_),
    .X(_0545_));
 sky130_fd_sc_hd__a211o_1 _3642_ (.A1(_2746_),
    .A2(_0541_),
    .B1(_0542_),
    .C1(_0544_),
    .X(_0546_));
 sky130_fd_sc_hd__o21a_4 _3643_ (.A1(_2771_),
    .A2(_0525_),
    .B1(_0546_),
    .X(_0547_));
 sky130_fd_sc_hd__o41a_4 _3644_ (.A1(_2525_),
    .A2(net293),
    .A3(net144),
    .A4(_2779_),
    .B1(net319),
    .X(_0548_));
 sky130_fd_sc_hd__and4_1 _3645_ (.A(_0517_),
    .B(_0524_),
    .C(_0536_),
    .D(_0543_),
    .X(_0549_));
 sky130_fd_sc_hd__o211a_4 _3646_ (.A1(_2783_),
    .A2(net154),
    .B1(_0549_),
    .C1(_0519_),
    .X(_0550_));
 sky130_fd_sc_hd__a311o_1 _3647_ (.A1(_2688_),
    .A2(_2710_),
    .A3(_2782_),
    .B1(net177),
    .C1(_2525_),
    .X(_0551_));
 sky130_fd_sc_hd__a311o_1 _3648_ (.A1(_2655_),
    .A2(_2664_),
    .A3(_2693_),
    .B1(_0514_),
    .C1(net177),
    .X(_0552_));
 sky130_fd_sc_hd__a41o_4 _3649_ (.A1(_0537_),
    .A2(_0545_),
    .A3(_0551_),
    .A4(_0552_),
    .B1(net304),
    .X(_0553_));
 sky130_fd_sc_hd__o21ai_4 _3650_ (.A1(net305),
    .A2(_0527_),
    .B1(_0548_),
    .Y(_0554_));
 sky130_fd_sc_hd__inv_2 _3651_ (.A(_0554_),
    .Y(_0555_));
 sky130_fd_sc_hd__nor2_1 _3652_ (.A(net67),
    .B(_0514_),
    .Y(_0556_));
 sky130_fd_sc_hd__or2_1 _3653_ (.A(net67),
    .B(_0514_),
    .X(_0557_));
 sky130_fd_sc_hd__nor2_8 _3654_ (.A(_2807_),
    .B(_0514_),
    .Y(_0558_));
 sky130_fd_sc_hd__o221a_1 _3655_ (.A1(net263),
    .A2(net69),
    .B1(_2804_),
    .B2(_0557_),
    .C1(_0558_),
    .X(_0559_));
 sky130_fd_sc_hd__and2_1 _3656_ (.A(_0554_),
    .B(_0559_),
    .X(_0560_));
 sky130_fd_sc_hd__a221o_1 _3657_ (.A1(_0528_),
    .A2(_0547_),
    .B1(_0555_),
    .B2(\as2650.r123_2[0][0] ),
    .C1(_0560_),
    .X(_0037_));
 sky130_fd_sc_hd__o211a_1 _3658_ (.A1(_2818_),
    .A2(_0557_),
    .B1(_0558_),
    .C1(_2814_),
    .X(_0561_));
 sky130_fd_sc_hd__or2_1 _3659_ (.A(_2822_),
    .B(_0529_),
    .X(_0562_));
 sky130_fd_sc_hd__o211a_1 _3660_ (.A1(net345),
    .A2(_0530_),
    .B1(_0562_),
    .C1(_0517_),
    .X(_0563_));
 sky130_fd_sc_hd__a21o_1 _3661_ (.A1(net106),
    .A2(_0516_),
    .B1(_0523_),
    .X(_0564_));
 sky130_fd_sc_hd__o22a_1 _3662_ (.A1(net114),
    .A2(_0524_),
    .B1(_0563_),
    .B2(_0564_),
    .X(_0565_));
 sky130_fd_sc_hd__mux2_1 _3663_ (.A0(net258),
    .A1(_0565_),
    .S(_0519_),
    .X(_0566_));
 sky130_fd_sc_hd__or2_1 _3664_ (.A(_2834_),
    .B(_0522_),
    .X(_0567_));
 sky130_fd_sc_hd__o211a_1 _3665_ (.A1(_0521_),
    .A2(_0566_),
    .B1(_0567_),
    .C1(_0539_),
    .X(_0568_));
 sky130_fd_sc_hd__a211o_1 _3666_ (.A1(_2838_),
    .A2(_0541_),
    .B1(_0544_),
    .C1(_0568_),
    .X(_0569_));
 sky130_fd_sc_hd__o21a_4 _3667_ (.A1(_2856_),
    .A2(_0525_),
    .B1(_0569_),
    .X(_0570_));
 sky130_fd_sc_hd__a211o_1 _3668_ (.A1(_0528_),
    .A2(_0570_),
    .B1(_0561_),
    .C1(_0555_),
    .X(_0571_));
 sky130_fd_sc_hd__o21a_1 _3669_ (.A1(\as2650.r123_2[0][1] ),
    .A2(_0554_),
    .B1(_0571_),
    .X(_0038_));
 sky130_fd_sc_hd__or2_1 _3670_ (.A(_2865_),
    .B(_0557_),
    .X(_0572_));
 sky130_fd_sc_hd__a31o_1 _3671_ (.A1(_2859_),
    .A2(_0558_),
    .A3(_0572_),
    .B1(_0548_),
    .X(_0573_));
 sky130_fd_sc_hd__or2_1 _3672_ (.A(_2870_),
    .B(_0529_),
    .X(_0574_));
 sky130_fd_sc_hd__o211a_1 _3673_ (.A1(net342),
    .A2(_0530_),
    .B1(_0574_),
    .C1(_0517_),
    .X(_0575_));
 sky130_fd_sc_hd__a21o_1 _3674_ (.A1(net103),
    .A2(_0516_),
    .B1(_0523_),
    .X(_0576_));
 sky130_fd_sc_hd__o22a_1 _3675_ (.A1(net111),
    .A2(_0524_),
    .B1(_0575_),
    .B2(_0576_),
    .X(_0577_));
 sky130_fd_sc_hd__mux2_1 _3676_ (.A0(net253),
    .A1(_0577_),
    .S(_0519_),
    .X(_0578_));
 sky130_fd_sc_hd__or2_1 _3677_ (.A(_2882_),
    .B(_0522_),
    .X(_0579_));
 sky130_fd_sc_hd__o211a_1 _3678_ (.A1(_0521_),
    .A2(_0578_),
    .B1(_0579_),
    .C1(_0539_),
    .X(_0580_));
 sky130_fd_sc_hd__a21o_1 _3679_ (.A1(_2886_),
    .A2(_0538_),
    .B1(_0580_),
    .X(_0581_));
 sky130_fd_sc_hd__mux2_8 _3680_ (.A0(_2903_),
    .A1(_0581_),
    .S(_0525_),
    .X(_0582_));
 sky130_fd_sc_hd__o221a_1 _3681_ (.A1(\as2650.r123_2[0][2] ),
    .A2(_0554_),
    .B1(_0582_),
    .B2(_0553_),
    .C1(_0573_),
    .X(_0039_));
 sky130_fd_sc_hd__nand2_1 _3682_ (.A(_2910_),
    .B(_0556_),
    .Y(_0583_));
 sky130_fd_sc_hd__a31o_1 _3683_ (.A1(_2906_),
    .A2(_0558_),
    .A3(_0583_),
    .B1(_0548_),
    .X(_0584_));
 sky130_fd_sc_hd__or2_1 _3684_ (.A(_2914_),
    .B(_0529_),
    .X(_0585_));
 sky130_fd_sc_hd__o211a_1 _3685_ (.A1(net339),
    .A2(_0530_),
    .B1(_0585_),
    .C1(_0517_),
    .X(_0586_));
 sky130_fd_sc_hd__a211o_1 _3686_ (.A1(net99),
    .A2(_0516_),
    .B1(_0523_),
    .C1(_0586_),
    .X(_0587_));
 sky130_fd_sc_hd__o21a_1 _3687_ (.A1(net106),
    .A2(_0524_),
    .B1(_0519_),
    .X(_0588_));
 sky130_fd_sc_hd__a221o_1 _3688_ (.A1(net246),
    .A2(_0518_),
    .B1(_0587_),
    .B2(_0588_),
    .C1(_0521_),
    .X(_0589_));
 sky130_fd_sc_hd__o211a_1 _3689_ (.A1(_2932_),
    .A2(_0522_),
    .B1(_0539_),
    .C1(_0589_),
    .X(_0590_));
 sky130_fd_sc_hd__a21o_1 _3690_ (.A1(_0288_),
    .A2(_0538_),
    .B1(_0590_),
    .X(_0591_));
 sky130_fd_sc_hd__mux2_8 _3691_ (.A0(_0309_),
    .A1(_0591_),
    .S(_0525_),
    .X(_0592_));
 sky130_fd_sc_hd__o221a_1 _3692_ (.A1(\as2650.r123_2[0][3] ),
    .A2(_0554_),
    .B1(_0592_),
    .B2(_0553_),
    .C1(_0584_),
    .X(_0040_));
 sky130_fd_sc_hd__nand2_1 _3693_ (.A(_0317_),
    .B(_0556_),
    .Y(_0593_));
 sky130_fd_sc_hd__a31o_1 _3694_ (.A1(_0312_),
    .A2(_0558_),
    .A3(_0593_),
    .B1(_0548_),
    .X(_0594_));
 sky130_fd_sc_hd__and2_1 _3695_ (.A(_0321_),
    .B(_0530_),
    .X(_0595_));
 sky130_fd_sc_hd__a21o_1 _3696_ (.A1(net335),
    .A2(_0529_),
    .B1(_0516_),
    .X(_0596_));
 sky130_fd_sc_hd__o221a_1 _3697_ (.A1(net96),
    .A2(_0517_),
    .B1(_0595_),
    .B2(_0596_),
    .C1(_0524_),
    .X(_0597_));
 sky130_fd_sc_hd__a211o_1 _3698_ (.A1(net103),
    .A2(_0523_),
    .B1(_0597_),
    .C1(_0518_),
    .X(_0598_));
 sky130_fd_sc_hd__o21ai_1 _3699_ (.A1(net245),
    .A2(_0519_),
    .B1(_0598_),
    .Y(_0599_));
 sky130_fd_sc_hd__nor2_1 _3700_ (.A(_0337_),
    .B(_0522_),
    .Y(_0600_));
 sky130_fd_sc_hd__a211o_1 _3701_ (.A1(_0522_),
    .A2(_0599_),
    .B1(_0600_),
    .C1(_0538_),
    .X(_0601_));
 sky130_fd_sc_hd__o21ai_2 _3702_ (.A1(_0341_),
    .A2(_0539_),
    .B1(_0601_),
    .Y(_0602_));
 sky130_fd_sc_hd__mux2_8 _3703_ (.A0(_0361_),
    .A1(_0602_),
    .S(_0525_),
    .X(_0603_));
 sky130_fd_sc_hd__o221a_1 _3704_ (.A1(\as2650.r123_2[0][4] ),
    .A2(_0554_),
    .B1(_0603_),
    .B2(_0553_),
    .C1(_0594_),
    .X(_0041_));
 sky130_fd_sc_hd__nor2_1 _3705_ (.A(_0381_),
    .B(_0529_),
    .Y(_0604_));
 sky130_fd_sc_hd__a211o_1 _3706_ (.A1(net332),
    .A2(_0529_),
    .B1(_0604_),
    .C1(_0516_),
    .X(_0605_));
 sky130_fd_sc_hd__o211a_1 _3707_ (.A1(net94),
    .A2(_0517_),
    .B1(_0524_),
    .C1(_0605_),
    .X(_0606_));
 sky130_fd_sc_hd__a211o_1 _3708_ (.A1(net99),
    .A2(_0523_),
    .B1(_0606_),
    .C1(_0518_),
    .X(_0607_));
 sky130_fd_sc_hd__o211a_1 _3709_ (.A1(net242),
    .A2(_0519_),
    .B1(_0522_),
    .C1(_0607_),
    .X(_0608_));
 sky130_fd_sc_hd__a21o_1 _3710_ (.A1(_0394_),
    .A2(_0521_),
    .B1(_0538_),
    .X(_0609_));
 sky130_fd_sc_hd__o22a_1 _3711_ (.A1(_0396_),
    .A2(_0539_),
    .B1(_0608_),
    .B2(_0609_),
    .X(_0610_));
 sky130_fd_sc_hd__mux2_8 _3712_ (.A0(_0414_),
    .A1(_0610_),
    .S(_0543_),
    .X(_0611_));
 sky130_fd_sc_hd__a31o_1 _3713_ (.A1(_0364_),
    .A2(_0371_),
    .A3(_0558_),
    .B1(_0548_),
    .X(_0612_));
 sky130_fd_sc_hd__o221a_1 _3714_ (.A1(\as2650.r123_2[0][5] ),
    .A2(_0554_),
    .B1(_0611_),
    .B2(_0553_),
    .C1(_0612_),
    .X(_0042_));
 sky130_fd_sc_hd__a31o_1 _3715_ (.A1(_0417_),
    .A2(_0423_),
    .A3(_0558_),
    .B1(_0548_),
    .X(_0613_));
 sky130_fd_sc_hd__a221o_1 _3716_ (.A1(net331),
    .A2(_0529_),
    .B1(_0531_),
    .B2(_0426_),
    .C1(_0516_),
    .X(_0614_));
 sky130_fd_sc_hd__o211a_1 _3717_ (.A1(net109),
    .A2(_0517_),
    .B1(_0524_),
    .C1(_0614_),
    .X(_0615_));
 sky130_fd_sc_hd__a211o_1 _3718_ (.A1(net96),
    .A2(_0523_),
    .B1(_0615_),
    .C1(_0518_),
    .X(_0616_));
 sky130_fd_sc_hd__o211a_1 _3719_ (.A1(net238),
    .A2(_0519_),
    .B1(_0522_),
    .C1(_0616_),
    .X(_0617_));
 sky130_fd_sc_hd__a211o_1 _3720_ (.A1(_0436_),
    .A2(_0521_),
    .B1(_0538_),
    .C1(_0617_),
    .X(_0618_));
 sky130_fd_sc_hd__o211a_1 _3721_ (.A1(_0439_),
    .A2(_0539_),
    .B1(_0543_),
    .C1(_0618_),
    .X(_0619_));
 sky130_fd_sc_hd__a21o_4 _3722_ (.A1(_0458_),
    .A2(_0544_),
    .B1(_0619_),
    .X(_0620_));
 sky130_fd_sc_hd__o221a_1 _3723_ (.A1(\as2650.r123_2[0][6] ),
    .A2(_0554_),
    .B1(_0620_),
    .B2(_0553_),
    .C1(_0613_),
    .X(_0043_));
 sky130_fd_sc_hd__a21o_1 _3724_ (.A1(net327),
    .A2(_0529_),
    .B1(_0516_),
    .X(_0621_));
 sky130_fd_sc_hd__a21o_1 _3725_ (.A1(_0463_),
    .A2(_0530_),
    .B1(_0621_),
    .X(_0622_));
 sky130_fd_sc_hd__o211a_1 _3726_ (.A1(_0466_),
    .A2(_0517_),
    .B1(_0524_),
    .C1(_0622_),
    .X(_0623_));
 sky130_fd_sc_hd__a211o_1 _3727_ (.A1(net94),
    .A2(_0523_),
    .B1(_0623_),
    .C1(_0518_),
    .X(_0624_));
 sky130_fd_sc_hd__o211a_1 _3728_ (.A1(net234),
    .A2(_0519_),
    .B1(_0522_),
    .C1(_0624_),
    .X(_0625_));
 sky130_fd_sc_hd__a21o_1 _3729_ (.A1(_0474_),
    .A2(_0521_),
    .B1(_0625_),
    .X(_0626_));
 sky130_fd_sc_hd__mux2_1 _3730_ (.A0(_0626_),
    .A1(_0477_),
    .S(_0541_),
    .X(_0627_));
 sky130_fd_sc_hd__mux2_4 _3731_ (.A0(_0494_),
    .A1(_0627_),
    .S(_0543_),
    .X(_0628_));
 sky130_fd_sc_hd__a32o_1 _3732_ (.A1(net234),
    .A2(net67),
    .A3(_0558_),
    .B1(_0628_),
    .B2(_0528_),
    .X(_0629_));
 sky130_fd_sc_hd__mux2_1 _3733_ (.A0(\as2650.r123_2[0][7] ),
    .A1(_0629_),
    .S(_0554_),
    .X(_0044_));
 sky130_fd_sc_hd__nor2_4 _3734_ (.A(net303),
    .B(_2654_),
    .Y(_0630_));
 sky130_fd_sc_hd__nand2_8 _3735_ (.A(net209),
    .B(_2653_),
    .Y(_0631_));
 sky130_fd_sc_hd__nor2_1 _3736_ (.A(_2662_),
    .B(_0630_),
    .Y(_0632_));
 sky130_fd_sc_hd__nand2_4 _3737_ (.A(_2663_),
    .B(_0631_),
    .Y(_0633_));
 sky130_fd_sc_hd__and3_2 _3738_ (.A(_2663_),
    .B(_2679_),
    .C(_0631_),
    .X(_0634_));
 sky130_fd_sc_hd__nand2_1 _3739_ (.A(_2679_),
    .B(net55),
    .Y(_0635_));
 sky130_fd_sc_hd__nor2_8 _3740_ (.A(net208),
    .B(_2572_),
    .Y(_0636_));
 sky130_fd_sc_hd__or2_4 _3741_ (.A(net208),
    .B(_2572_),
    .X(_0637_));
 sky130_fd_sc_hd__nor2_4 _3742_ (.A(net231),
    .B(net204),
    .Y(_0638_));
 sky130_fd_sc_hd__nand2_2 _3743_ (.A(net207),
    .B(net228),
    .Y(_0639_));
 sky130_fd_sc_hd__nor3_4 _3744_ (.A(net209),
    .B(_2851_),
    .C(net151),
    .Y(_0640_));
 sky130_fd_sc_hd__or3_4 _3745_ (.A(net209),
    .B(_2851_),
    .C(net152),
    .X(_0641_));
 sky130_fd_sc_hd__o211a_2 _3746_ (.A1(net196),
    .A2(_0641_),
    .B1(net92),
    .C1(_0634_),
    .X(_0642_));
 sky130_fd_sc_hd__inv_2 _3747_ (.A(_0642_),
    .Y(_0643_));
 sky130_fd_sc_hd__nor2_2 _3748_ (.A(_2578_),
    .B(_0641_),
    .Y(_0644_));
 sky130_fd_sc_hd__nand2_4 _3749_ (.A(_2577_),
    .B(_0640_),
    .Y(_0645_));
 sky130_fd_sc_hd__o21ai_1 _3750_ (.A1(_0642_),
    .A2(_0644_),
    .B1(_2609_),
    .Y(_0646_));
 sky130_fd_sc_hd__nor2_1 _3751_ (.A(_2579_),
    .B(net69),
    .Y(_0647_));
 sky130_fd_sc_hd__nor2_2 _3752_ (.A(_2579_),
    .B(_2808_),
    .Y(_0648_));
 sky130_fd_sc_hd__and3_1 _3753_ (.A(_2573_),
    .B(net201),
    .C(net196),
    .X(_0649_));
 sky130_fd_sc_hd__and3_1 _3754_ (.A(_2573_),
    .B(net201),
    .C(_2702_),
    .X(_0650_));
 sky130_fd_sc_hd__or2_2 _3755_ (.A(_0649_),
    .B(net65),
    .X(_0651_));
 sky130_fd_sc_hd__nand2_1 _3756_ (.A(net81),
    .B(_0651_),
    .Y(_0652_));
 sky130_fd_sc_hd__and4_2 _3757_ (.A(net226),
    .B(net201),
    .C(_2702_),
    .D(_2759_),
    .X(_0653_));
 sky130_fd_sc_hd__nor2_1 _3758_ (.A(_0649_),
    .B(_0653_),
    .Y(_0654_));
 sky130_fd_sc_hd__nor2_1 _3759_ (.A(_2579_),
    .B(net64),
    .Y(_0655_));
 sky130_fd_sc_hd__or2_1 _3760_ (.A(_2579_),
    .B(_0651_),
    .X(_0656_));
 sky130_fd_sc_hd__nor2_1 _3761_ (.A(_0653_),
    .B(_0656_),
    .Y(_0657_));
 sky130_fd_sc_hd__nand2_1 _3762_ (.A(_0648_),
    .B(_0657_),
    .Y(_0658_));
 sky130_fd_sc_hd__or2_1 _3763_ (.A(net291),
    .B(_0636_),
    .X(_0659_));
 sky130_fd_sc_hd__and3_4 _3764_ (.A(net79),
    .B(_2679_),
    .C(_0637_),
    .X(_0660_));
 sky130_fd_sc_hd__or3b_1 _3765_ (.A(_0633_),
    .B(_0658_),
    .C_N(_0660_),
    .X(_0661_));
 sky130_fd_sc_hd__or2_1 _3766_ (.A(\as2650.psl[6] ),
    .B(net308),
    .X(_0662_));
 sky130_fd_sc_hd__nand2_1 _3767_ (.A(\as2650.psl[6] ),
    .B(net308),
    .Y(_0663_));
 sky130_fd_sc_hd__or2_1 _3768_ (.A(\as2650.psl[7] ),
    .B(net304),
    .X(_0664_));
 sky130_fd_sc_hd__nand2_1 _3769_ (.A(\as2650.psl[7] ),
    .B(net304),
    .Y(_0665_));
 sky130_fd_sc_hd__a22o_1 _3770_ (.A1(_0662_),
    .A2(_0663_),
    .B1(_0664_),
    .B2(_0665_),
    .X(_0666_));
 sky130_fd_sc_hd__nand2_1 _3771_ (.A(_2584_),
    .B(_0666_),
    .Y(_0667_));
 sky130_fd_sc_hd__and3_1 _3772_ (.A(net165),
    .B(net163),
    .C(_0667_),
    .X(_0668_));
 sky130_fd_sc_hd__a21oi_1 _3773_ (.A1(net300),
    .A2(_0668_),
    .B1(_0637_),
    .Y(_0669_));
 sky130_fd_sc_hd__or4b_1 _3774_ (.A(\as2650.halted ),
    .B(net148),
    .C(_0635_),
    .D_N(_0648_),
    .X(_0670_));
 sky130_fd_sc_hd__or3_1 _3775_ (.A(net152),
    .B(_0669_),
    .C(_0670_),
    .X(_0671_));
 sky130_fd_sc_hd__and4b_1 _3776_ (.A_N(_0671_),
    .B(_0661_),
    .C(_0652_),
    .D(_0646_),
    .X(_0672_));
 sky130_fd_sc_hd__and3_2 _3777_ (.A(net242),
    .B(net165),
    .C(net163),
    .X(_0673_));
 sky130_fd_sc_hd__nor2_4 _3778_ (.A(_2645_),
    .B(_0641_),
    .Y(_0674_));
 sky130_fd_sc_hd__nand2_1 _3779_ (.A(net332),
    .B(_0674_),
    .Y(_0675_));
 sky130_fd_sc_hd__o211a_1 _3780_ (.A1(\as2650.psu[5] ),
    .A2(net333),
    .B1(net144),
    .C1(_0675_),
    .X(_0676_));
 sky130_fd_sc_hd__o21ai_1 _3781_ (.A1(_0673_),
    .A2(_0676_),
    .B1(net92),
    .Y(_0677_));
 sky130_fd_sc_hd__o21ai_1 _3782_ (.A1(\as2650.psu[5] ),
    .A2(_0672_),
    .B1(net319),
    .Y(_0678_));
 sky130_fd_sc_hd__a21oi_1 _3783_ (.A1(_0672_),
    .A2(_0677_),
    .B1(_0678_),
    .Y(_0045_));
 sky130_fd_sc_hd__or2_4 _3784_ (.A(net221),
    .B(net169),
    .X(_0679_));
 sky130_fd_sc_hd__or2_4 _3785_ (.A(net48),
    .B(_0679_),
    .X(_0680_));
 sky130_fd_sc_hd__o21a_4 _3786_ (.A1(_2631_),
    .A2(_0679_),
    .B1(_0680_),
    .X(_0681_));
 sky130_fd_sc_hd__mux2_1 _3787_ (.A0(_2625_),
    .A1(\as2650.stack[3][8] ),
    .S(_0681_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _3788_ (.A0(_2633_),
    .A1(\as2650.stack[3][9] ),
    .S(_0681_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _3789_ (.A0(_2635_),
    .A1(\as2650.stack[3][10] ),
    .S(_0681_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _3790_ (.A0(_2637_),
    .A1(\as2650.stack[3][11] ),
    .S(_0681_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _3791_ (.A0(_2639_),
    .A1(\as2650.stack[3][12] ),
    .S(_0681_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _3792_ (.A0(_2641_),
    .A1(\as2650.stack[3][13] ),
    .S(_0681_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _3793_ (.A0(_2643_),
    .A1(\as2650.stack[3][14] ),
    .S(_0681_),
    .X(_0052_));
 sky130_fd_sc_hd__nor2_1 _3794_ (.A(_2593_),
    .B(_2669_),
    .Y(_0682_));
 sky130_fd_sc_hd__or2_4 _3795_ (.A(_2593_),
    .B(_2669_),
    .X(_0683_));
 sky130_fd_sc_hd__nor2_8 _3796_ (.A(\as2650.cycle[7] ),
    .B(_0683_),
    .Y(_0684_));
 sky130_fd_sc_hd__inv_2 _3797_ (.A(_0684_),
    .Y(_0685_));
 sky130_fd_sc_hd__nor2_8 _3798_ (.A(net74),
    .B(_0684_),
    .Y(_0686_));
 sky130_fd_sc_hd__or2_4 _3799_ (.A(net74),
    .B(_0684_),
    .X(_0687_));
 sky130_fd_sc_hd__or4b_4 _3800_ (.A(_2536_),
    .B(\as2650.cycle[1] ),
    .C(net290),
    .D_N(_2562_),
    .X(_0688_));
 sky130_fd_sc_hd__inv_2 _3801_ (.A(_0688_),
    .Y(_0689_));
 sky130_fd_sc_hd__or4_4 _3802_ (.A(net131),
    .B(_2606_),
    .C(_2612_),
    .D(_0689_),
    .X(_0690_));
 sky130_fd_sc_hd__or3_1 _3803_ (.A(_2684_),
    .B(_0687_),
    .C(_0690_),
    .X(_0691_));
 sky130_fd_sc_hd__or3_2 _3804_ (.A(net223),
    .B(net150),
    .C(_0691_),
    .X(_0692_));
 sky130_fd_sc_hd__nor2_2 _3805_ (.A(net223),
    .B(net80),
    .Y(_0693_));
 sky130_fd_sc_hd__nand2_8 _3806_ (.A(net202),
    .B(net140),
    .Y(_0694_));
 sky130_fd_sc_hd__nor2_2 _3807_ (.A(_0685_),
    .B(_0694_),
    .Y(_0695_));
 sky130_fd_sc_hd__nor2_4 _3808_ (.A(\as2650.cycle[1] ),
    .B(net164),
    .Y(_0696_));
 sky130_fd_sc_hd__nand2_8 _3809_ (.A(_2537_),
    .B(net165),
    .Y(_0697_));
 sky130_fd_sc_hd__nor2_2 _3810_ (.A(net164),
    .B(_2593_),
    .Y(_0698_));
 sky130_fd_sc_hd__or2_4 _3811_ (.A(net164),
    .B(_2593_),
    .X(_0699_));
 sky130_fd_sc_hd__nor2_1 _3812_ (.A(net222),
    .B(net90),
    .Y(_0700_));
 sky130_fd_sc_hd__nand2_2 _3813_ (.A(net203),
    .B(net88),
    .Y(_0701_));
 sky130_fd_sc_hd__nor2_2 _3814_ (.A(\as2650.cycle[6] ),
    .B(_0688_),
    .Y(_0702_));
 sky130_fd_sc_hd__or2_2 _3815_ (.A(\as2650.cycle[6] ),
    .B(_0688_),
    .X(_0703_));
 sky130_fd_sc_hd__nand2_1 _3816_ (.A(net326),
    .B(net87),
    .Y(_0704_));
 sky130_fd_sc_hd__nor2_1 _3817_ (.A(_0701_),
    .B(_0704_),
    .Y(_0705_));
 sky130_fd_sc_hd__nor2_1 _3818_ (.A(_0695_),
    .B(_0705_),
    .Y(_0706_));
 sky130_fd_sc_hd__nand2_1 _3819_ (.A(net294),
    .B(net74),
    .Y(_0707_));
 sky130_fd_sc_hd__nor2_1 _3820_ (.A(net222),
    .B(_0707_),
    .Y(_0708_));
 sky130_fd_sc_hd__nand2b_2 _3821_ (.A_N(\as2650.cycle[0] ),
    .B(_2606_),
    .Y(_0709_));
 sky130_fd_sc_hd__or2_4 _3822_ (.A(net224),
    .B(_0709_),
    .X(_0710_));
 sky130_fd_sc_hd__and2_4 _3823_ (.A(net165),
    .B(_2668_),
    .X(_0711_));
 sky130_fd_sc_hd__nand2_8 _3824_ (.A(net165),
    .B(_2668_),
    .Y(_0712_));
 sky130_fd_sc_hd__nor2_2 _3825_ (.A(net222),
    .B(_2610_),
    .Y(_0713_));
 sky130_fd_sc_hd__nor2_2 _3826_ (.A(_0711_),
    .B(_0713_),
    .Y(_0714_));
 sky130_fd_sc_hd__or3b_4 _3827_ (.A(_2600_),
    .B(net303),
    .C_N(net298),
    .X(_0715_));
 sky130_fd_sc_hd__nor2_2 _3828_ (.A(net224),
    .B(_2607_),
    .Y(_0716_));
 sky130_fd_sc_hd__nor2_8 _3829_ (.A(net231),
    .B(net92),
    .Y(_0717_));
 sky130_fd_sc_hd__nand2_4 _3830_ (.A(net207),
    .B(_0636_),
    .Y(_0718_));
 sky130_fd_sc_hd__nor4_2 _3831_ (.A(_2536_),
    .B(net222),
    .C(_2593_),
    .D(_2669_),
    .Y(_0719_));
 sky130_fd_sc_hd__nand2_4 _3832_ (.A(\as2650.cycle[6] ),
    .B(_0689_),
    .Y(_0720_));
 sky130_fd_sc_hd__or4_1 _3833_ (.A(net292),
    .B(_0716_),
    .C(_0717_),
    .D(_0719_),
    .X(_0721_));
 sky130_fd_sc_hd__nor2_4 _3834_ (.A(net223),
    .B(net141),
    .Y(_0722_));
 sky130_fd_sc_hd__or2_2 _3835_ (.A(net224),
    .B(net142),
    .X(_0723_));
 sky130_fd_sc_hd__nor2_1 _3836_ (.A(net89),
    .B(net62),
    .Y(_0724_));
 sky130_fd_sc_hd__nor2_8 _3837_ (.A(\as2650.ins_reg[3] ),
    .B(_0636_),
    .Y(_0725_));
 sky130_fd_sc_hd__nand2_1 _3838_ (.A(_2545_),
    .B(_0637_),
    .Y(_0726_));
 sky130_fd_sc_hd__and3_2 _3839_ (.A(_2679_),
    .B(net92),
    .C(net153),
    .X(_0727_));
 sky130_fd_sc_hd__inv_2 _3840_ (.A(_0727_),
    .Y(_0728_));
 sky130_fd_sc_hd__and3_1 _3841_ (.A(_2696_),
    .B(net52),
    .C(_0728_),
    .X(_0729_));
 sky130_fd_sc_hd__mux2_8 _3842_ (.A0(net113),
    .A1(net262),
    .S(_2676_),
    .X(_0730_));
 sky130_fd_sc_hd__nand2_1 _3843_ (.A(_0710_),
    .B(_0712_),
    .Y(_0731_));
 sky130_fd_sc_hd__o221ai_2 _3844_ (.A1(net224),
    .A2(net118),
    .B1(_0715_),
    .B2(net79),
    .C1(_2682_),
    .Y(_0732_));
 sky130_fd_sc_hd__a211o_1 _3845_ (.A1(_2692_),
    .A2(net151),
    .B1(net62),
    .C1(_0727_),
    .X(_0733_));
 sky130_fd_sc_hd__or4_1 _3846_ (.A(_0708_),
    .B(_0731_),
    .C(_0732_),
    .D(_0733_),
    .X(_0734_));
 sky130_fd_sc_hd__and4b_1 _3847_ (.A_N(_0734_),
    .B(net88),
    .C(_2696_),
    .D(_0706_),
    .X(_0735_));
 sky130_fd_sc_hd__and3b_4 _3848_ (.A_N(_0721_),
    .B(_0735_),
    .C(_0692_),
    .X(_0736_));
 sky130_fd_sc_hd__mux2_1 _3849_ (.A0(net12),
    .A1(_0730_),
    .S(_0736_),
    .X(_0737_));
 sky130_fd_sc_hd__and2_1 _3850_ (.A(net313),
    .B(_0737_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_4 _3851_ (.A0(net112),
    .A1(net258),
    .S(_2676_),
    .X(_0738_));
 sky130_fd_sc_hd__mux2_1 _3852_ (.A0(net23),
    .A1(_0738_),
    .S(_0736_),
    .X(_0739_));
 sky130_fd_sc_hd__and2_1 _3853_ (.A(net313),
    .B(_0739_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_4 _3854_ (.A0(_2826_),
    .A1(net250),
    .S(_2676_),
    .X(_0740_));
 sky130_fd_sc_hd__mux2_1 _3855_ (.A0(net31),
    .A1(_0740_),
    .S(_0736_),
    .X(_0741_));
 sky130_fd_sc_hd__and2_1 _3856_ (.A(net313),
    .B(_0741_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_2 _3857_ (.A0(net102),
    .A1(net246),
    .S(_2676_),
    .X(_0742_));
 sky130_fd_sc_hd__mux2_1 _3858_ (.A0(net32),
    .A1(_0742_),
    .S(_0736_),
    .X(_0743_));
 sky130_fd_sc_hd__and2_1 _3859_ (.A(net313),
    .B(_0743_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_4 _3860_ (.A0(net100),
    .A1(net243),
    .S(_2676_),
    .X(_0744_));
 sky130_fd_sc_hd__mux2_1 _3861_ (.A0(net33),
    .A1(_0744_),
    .S(_0736_),
    .X(_0745_));
 sky130_fd_sc_hd__and2_1 _3862_ (.A(net313),
    .B(_0745_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_2 _3863_ (.A0(net96),
    .A1(\as2650.r0[5] ),
    .S(_2676_),
    .X(_0746_));
 sky130_fd_sc_hd__mux2_1 _3864_ (.A0(net34),
    .A1(_0746_),
    .S(_0736_),
    .X(_0747_));
 sky130_fd_sc_hd__and2_1 _3865_ (.A(net313),
    .B(_0747_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_2 _3866_ (.A0(net95),
    .A1(net238),
    .S(_2676_),
    .X(_0748_));
 sky130_fd_sc_hd__mux2_1 _3867_ (.A0(net35),
    .A1(_0748_),
    .S(_0736_),
    .X(_0749_));
 sky130_fd_sc_hd__and2_1 _3868_ (.A(net313),
    .B(_0749_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_2 _3869_ (.A0(net110),
    .A1(net232),
    .S(_2676_),
    .X(_0750_));
 sky130_fd_sc_hd__mux2_1 _3870_ (.A0(net36),
    .A1(_0750_),
    .S(_0736_),
    .X(_0751_));
 sky130_fd_sc_hd__and2_1 _3871_ (.A(net313),
    .B(_0751_),
    .X(_0060_));
 sky130_fd_sc_hd__or3_4 _3872_ (.A(net219),
    .B(net166),
    .C(net48),
    .X(_0752_));
 sky130_fd_sc_hd__or3_4 _3873_ (.A(net219),
    .B(net167),
    .C(_2631_),
    .X(_0753_));
 sky130_fd_sc_hd__nand2_8 _3874_ (.A(_0752_),
    .B(_0753_),
    .Y(_0754_));
 sky130_fd_sc_hd__mux2_1 _3875_ (.A0(\as2650.stack[2][8] ),
    .A1(_2625_),
    .S(_0754_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _3876_ (.A0(\as2650.stack[2][9] ),
    .A1(_2633_),
    .S(_0754_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _3877_ (.A0(\as2650.stack[2][10] ),
    .A1(_2635_),
    .S(_0754_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _3878_ (.A0(\as2650.stack[2][11] ),
    .A1(_2637_),
    .S(_0754_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _3879_ (.A0(\as2650.stack[2][12] ),
    .A1(_2639_),
    .S(_0754_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _3880_ (.A0(\as2650.stack[2][13] ),
    .A1(_2641_),
    .S(_0754_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _3881_ (.A0(\as2650.stack[2][14] ),
    .A1(_2643_),
    .S(_0754_),
    .X(_0067_));
 sky130_fd_sc_hd__or2_1 _3882_ (.A(\as2650.holding_reg[7] ),
    .B(net198),
    .X(_0755_));
 sky130_fd_sc_hd__o21ai_2 _3883_ (.A1(net200),
    .A2(net109),
    .B1(_0755_),
    .Y(_0756_));
 sky130_fd_sc_hd__o21ba_1 _3884_ (.A1(_2755_),
    .A2(_2842_),
    .B1_N(_2895_),
    .X(_0757_));
 sky130_fd_sc_hd__o21a_1 _3885_ (.A1(_2890_),
    .A2(_0757_),
    .B1(_0296_),
    .X(_0758_));
 sky130_fd_sc_hd__o21ai_1 _3886_ (.A1(_0293_),
    .A2(_0758_),
    .B1(_0346_),
    .Y(_0759_));
 sky130_fd_sc_hd__a21o_1 _3887_ (.A1(_0345_),
    .A2(_0759_),
    .B1(_0402_),
    .X(_0760_));
 sky130_fd_sc_hd__a21bo_1 _3888_ (.A1(_0401_),
    .A2(_0760_),
    .B1_N(_0448_),
    .X(_0761_));
 sky130_fd_sc_hd__a32o_1 _3889_ (.A1(_0444_),
    .A2(_0482_),
    .A3(_0761_),
    .B1(_0489_),
    .B2(_0480_),
    .X(_0762_));
 sky130_fd_sc_hd__nor2_1 _3890_ (.A(\as2650.psl[1] ),
    .B(_0482_),
    .Y(_0763_));
 sky130_fd_sc_hd__a211o_1 _3891_ (.A1(_0482_),
    .A2(_0483_),
    .B1(_0762_),
    .C1(_0763_),
    .X(_0764_));
 sky130_fd_sc_hd__nand2_1 _3892_ (.A(_0762_),
    .B(_0763_),
    .Y(_0765_));
 sky130_fd_sc_hd__a31o_1 _3893_ (.A1(_2697_),
    .A2(_0764_),
    .A3(_0765_),
    .B1(net82),
    .X(_0766_));
 sky130_fd_sc_hd__nand3b_1 _3894_ (.A_N(_2890_),
    .B(_0345_),
    .C(_0401_),
    .Y(_0767_));
 sky130_fd_sc_hd__or4_1 _3895_ (.A(net82),
    .B(_2842_),
    .C(_0443_),
    .D(_0481_),
    .X(_0768_));
 sky130_fd_sc_hd__or4b_1 _3896_ (.A(_0293_),
    .B(_0767_),
    .C(_0768_),
    .D_N(_2758_),
    .X(_0769_));
 sky130_fd_sc_hd__or4_1 _3897_ (.A(_2771_),
    .B(_2856_),
    .C(_2903_),
    .D(_0309_),
    .X(_0770_));
 sky130_fd_sc_hd__or4_1 _3898_ (.A(_0361_),
    .B(_0414_),
    .C(_0458_),
    .D(_0770_),
    .X(_0771_));
 sky130_fd_sc_hd__nor2_1 _3899_ (.A(_2697_),
    .B(_0494_),
    .Y(_0772_));
 sky130_fd_sc_hd__a22o_1 _3900_ (.A1(_0766_),
    .A2(_0769_),
    .B1(_0771_),
    .B2(_0772_),
    .X(_0773_));
 sky130_fd_sc_hd__or4_4 _3901_ (.A(net226),
    .B(net301),
    .C(net299),
    .D(net298),
    .X(_0774_));
 sky130_fd_sc_hd__inv_2 _3902_ (.A(_0774_),
    .Y(_0775_));
 sky130_fd_sc_hd__or2_1 _3903_ (.A(net109),
    .B(_0774_),
    .X(_0776_));
 sky130_fd_sc_hd__or4_1 _3904_ (.A(net238),
    .B(\as2650.r0[5] ),
    .C(net245),
    .D(net249),
    .X(_0777_));
 sky130_fd_sc_hd__o41a_1 _3905_ (.A1(net253),
    .A2(net258),
    .A3(net262),
    .A4(_0777_),
    .B1(_2530_),
    .X(_0778_));
 sky130_fd_sc_hd__a2bb2o_1 _3906_ (.A1_N(_0431_),
    .A2_N(_0776_),
    .B1(_0778_),
    .B2(_0774_),
    .X(_0779_));
 sky130_fd_sc_hd__o211a_1 _3907_ (.A1(net146),
    .A2(_0779_),
    .B1(_0773_),
    .C1(net204),
    .X(_0780_));
 sky130_fd_sc_hd__and3_1 _3908_ (.A(net148),
    .B(_0634_),
    .C(_0725_),
    .X(_0781_));
 sky130_fd_sc_hd__and4_1 _3909_ (.A(net226),
    .B(net201),
    .C(net196),
    .D(_2759_),
    .X(_0782_));
 sky130_fd_sc_hd__or2_1 _3910_ (.A(_0658_),
    .B(_0782_),
    .X(_0783_));
 sky130_fd_sc_hd__nor2_1 _3911_ (.A(_2571_),
    .B(net152),
    .Y(_0784_));
 sky130_fd_sc_hd__and4_4 _3912_ (.A(_2806_),
    .B(net55),
    .C(_0660_),
    .D(_0784_),
    .X(_0785_));
 sky130_fd_sc_hd__inv_2 _3913_ (.A(_0785_),
    .Y(_0786_));
 sky130_fd_sc_hd__o2bb2a_1 _3914_ (.A1_N(net226),
    .A2_N(_0781_),
    .B1(_0783_),
    .B2(_0786_),
    .X(_0787_));
 sky130_fd_sc_hd__and3_1 _3915_ (.A(net148),
    .B(net115),
    .C(net153),
    .X(_0788_));
 sky130_fd_sc_hd__nor2_1 _3916_ (.A(net80),
    .B(_2664_),
    .Y(_0789_));
 sky130_fd_sc_hd__nor2_2 _3917_ (.A(net197),
    .B(_2600_),
    .Y(_0790_));
 sky130_fd_sc_hd__nor2_1 _3918_ (.A(net230),
    .B(_0715_),
    .Y(_0791_));
 sky130_fd_sc_hd__nor2_1 _3919_ (.A(_0789_),
    .B(_0791_),
    .Y(_0792_));
 sky130_fd_sc_hd__nand2_4 _3920_ (.A(net143),
    .B(_0725_),
    .Y(_0793_));
 sky130_fd_sc_hd__inv_2 _3921_ (.A(_0793_),
    .Y(_0794_));
 sky130_fd_sc_hd__nand2_1 _3922_ (.A(net226),
    .B(net146),
    .Y(_0795_));
 sky130_fd_sc_hd__nor2_1 _3923_ (.A(_2692_),
    .B(_2776_),
    .Y(_0796_));
 sky130_fd_sc_hd__or2_1 _3924_ (.A(net197),
    .B(_0796_),
    .X(_0797_));
 sky130_fd_sc_hd__o2bb2a_1 _3925_ (.A1_N(net62),
    .A2_N(_0797_),
    .B1(_0793_),
    .B2(_0631_),
    .X(_0798_));
 sky130_fd_sc_hd__or3_4 _3926_ (.A(net131),
    .B(_2612_),
    .C(_0694_),
    .X(_0799_));
 sky130_fd_sc_hd__or3_2 _3927_ (.A(net308),
    .B(net118),
    .C(_0641_),
    .X(_0800_));
 sky130_fd_sc_hd__o31a_1 _3928_ (.A1(net308),
    .A2(_2610_),
    .A3(_0641_),
    .B1(_0714_),
    .X(_0801_));
 sky130_fd_sc_hd__or3_4 _3929_ (.A(net226),
    .B(_2661_),
    .C(_2776_),
    .X(_0802_));
 sky130_fd_sc_hd__nor2_4 _3930_ (.A(net142),
    .B(_0802_),
    .Y(_0803_));
 sky130_fd_sc_hd__nor2_2 _3931_ (.A(net292),
    .B(_0803_),
    .Y(_0804_));
 sky130_fd_sc_hd__or2_2 _3932_ (.A(net230),
    .B(net142),
    .X(_0805_));
 sky130_fd_sc_hd__nand2_2 _3933_ (.A(net81),
    .B(_0653_),
    .Y(_0806_));
 sky130_fd_sc_hd__nand3_2 _3934_ (.A(_2693_),
    .B(_0774_),
    .C(_0802_),
    .Y(_0807_));
 sky130_fd_sc_hd__o32a_1 _3935_ (.A1(net300),
    .A2(net118),
    .A3(_0643_),
    .B1(_2681_),
    .B2(net150),
    .X(_0808_));
 sky130_fd_sc_hd__o221a_1 _3936_ (.A1(_0723_),
    .A2(_0807_),
    .B1(_0808_),
    .B2(net152),
    .C1(_0801_),
    .X(_0809_));
 sky130_fd_sc_hd__and3_1 _3937_ (.A(_0799_),
    .B(_0804_),
    .C(_0809_),
    .X(_0810_));
 sky130_fd_sc_hd__and4_1 _3938_ (.A(net194),
    .B(net92),
    .C(_0648_),
    .D(net88),
    .X(_0811_));
 sky130_fd_sc_hd__o2111a_1 _3939_ (.A1(net142),
    .A2(_2682_),
    .B1(_0792_),
    .C1(_0806_),
    .D1(_0811_),
    .X(_0812_));
 sky130_fd_sc_hd__and4_2 _3940_ (.A(_0787_),
    .B(_0798_),
    .C(_0810_),
    .D(_0812_),
    .X(_0813_));
 sky130_fd_sc_hd__a211o_1 _3941_ (.A1(_2728_),
    .A2(_0374_),
    .B1(net94),
    .C1(_0631_),
    .X(_0814_));
 sky130_fd_sc_hd__or4_1 _3942_ (.A(net111),
    .B(net109),
    .C(_2826_),
    .D(net103),
    .X(_0815_));
 sky130_fd_sc_hd__or4_1 _3943_ (.A(net100),
    .B(net97),
    .C(net93),
    .D(_0815_),
    .X(_0816_));
 sky130_fd_sc_hd__or4_1 _3944_ (.A(net304),
    .B(net209),
    .C(net231),
    .D(_2556_),
    .X(_0817_));
 sky130_fd_sc_hd__mux2_1 _3945_ (.A0(net238),
    .A1(_0778_),
    .S(_0651_),
    .X(_0818_));
 sky130_fd_sc_hd__o2111a_1 _3946_ (.A1(\as2650.psl[6] ),
    .A2(net331),
    .B1(net146),
    .C1(_0817_),
    .D1(net308),
    .X(_0819_));
 sky130_fd_sc_hd__a22o_1 _3947_ (.A1(net82),
    .A2(_0818_),
    .B1(_0819_),
    .B2(_0640_),
    .X(_0820_));
 sky130_fd_sc_hd__a32o_1 _3948_ (.A1(_2662_),
    .A2(_0467_),
    .A3(_0816_),
    .B1(_0820_),
    .B2(net55),
    .X(_0821_));
 sky130_fd_sc_hd__or3b_1 _3949_ (.A(net115),
    .B(_0821_),
    .C_N(_0814_),
    .X(_0822_));
 sky130_fd_sc_hd__a21oi_1 _3950_ (.A1(net327),
    .A2(net115),
    .B1(net204),
    .Y(_0823_));
 sky130_fd_sc_hd__or4_1 _3951_ (.A(net350),
    .B(net345),
    .C(net343),
    .D(net339),
    .X(_0824_));
 sky130_fd_sc_hd__or4_1 _3952_ (.A(net335),
    .B(net333),
    .C(net331),
    .D(_0824_),
    .X(_0825_));
 sky130_fd_sc_hd__o211a_1 _3953_ (.A1(_2681_),
    .A2(_0825_),
    .B1(_0823_),
    .C1(_0822_),
    .X(_0826_));
 sky130_fd_sc_hd__or3b_1 _3954_ (.A(_0780_),
    .B(_0826_),
    .C_N(_0813_),
    .X(_0827_));
 sky130_fd_sc_hd__o211a_1 _3955_ (.A1(\as2650.psl[6] ),
    .A2(_0813_),
    .B1(_0827_),
    .C1(net320),
    .X(_0068_));
 sky130_fd_sc_hd__and3_1 _3956_ (.A(net303),
    .B(_2764_),
    .C(_0638_),
    .X(_0828_));
 sky130_fd_sc_hd__o22a_1 _3957_ (.A1(_2550_),
    .A2(net111),
    .B1(_2826_),
    .B2(_2551_),
    .X(_0829_));
 sky130_fd_sc_hd__o221a_1 _3958_ (.A1(_2553_),
    .A2(net101),
    .B1(net95),
    .B2(_2556_),
    .C1(_0829_),
    .X(_0830_));
 sky130_fd_sc_hd__o22a_1 _3959_ (.A1(_2552_),
    .A2(net103),
    .B1(net97),
    .B2(_2554_),
    .X(_0831_));
 sky130_fd_sc_hd__o221a_1 _3960_ (.A1(_2549_),
    .A2(net114),
    .B1(net110),
    .B2(net312),
    .C1(_0831_),
    .X(_0832_));
 sky130_fd_sc_hd__a21oi_1 _3961_ (.A1(_0830_),
    .A2(_0832_),
    .B1(_0828_),
    .Y(_0833_));
 sky130_fd_sc_hd__o22a_1 _3962_ (.A1(\as2650.psu[3] ),
    .A2(_2552_),
    .B1(_2553_),
    .B2(\as2650.psu[4] ),
    .X(_0834_));
 sky130_fd_sc_hd__o221a_1 _3963_ (.A1(\as2650.psu[0] ),
    .A2(_2549_),
    .B1(_2556_),
    .B2(net30),
    .C1(_0834_),
    .X(_0835_));
 sky130_fd_sc_hd__o221a_1 _3964_ (.A1(\as2650.psu[7] ),
    .A2(net311),
    .B1(_2554_),
    .B2(\as2650.psu[5] ),
    .C1(_0835_),
    .X(_0836_));
 sky130_fd_sc_hd__o221a_1 _3965_ (.A1(\as2650.psu[1] ),
    .A2(_2550_),
    .B1(_2551_),
    .B2(net221),
    .C1(_0836_),
    .X(_0837_));
 sky130_fd_sc_hd__or4_1 _3966_ (.A(net306),
    .B(net209),
    .C(_2765_),
    .D(net152),
    .X(_0838_));
 sky130_fd_sc_hd__nand2_1 _3967_ (.A(net196),
    .B(_0640_),
    .Y(_0839_));
 sky130_fd_sc_hd__nand2_1 _3968_ (.A(net306),
    .B(_0828_),
    .Y(_0840_));
 sky130_fd_sc_hd__o22a_1 _3969_ (.A1(\as2650.carry ),
    .A2(_2549_),
    .B1(_2554_),
    .B2(\as2650.psl[5] ),
    .X(_0841_));
 sky130_fd_sc_hd__o221a_1 _3970_ (.A1(\as2650.psl[7] ),
    .A2(net312),
    .B1(_2552_),
    .B2(\as2650.psl[3] ),
    .C1(_0841_),
    .X(_0842_));
 sky130_fd_sc_hd__o22a_1 _3971_ (.A1(\as2650.psl[1] ),
    .A2(_2550_),
    .B1(_2556_),
    .B2(\as2650.psl[6] ),
    .X(_0843_));
 sky130_fd_sc_hd__o22a_1 _3972_ (.A1(\as2650.overflow ),
    .A2(_2551_),
    .B1(_2553_),
    .B2(net213),
    .X(_0844_));
 sky130_fd_sc_hd__and3_1 _3973_ (.A(_0842_),
    .B(_0843_),
    .C(_0844_),
    .X(_0845_));
 sky130_fd_sc_hd__o221ai_1 _3974_ (.A1(_0837_),
    .A2(_0838_),
    .B1(_0840_),
    .B2(_0845_),
    .C1(_0839_),
    .Y(_0846_));
 sky130_fd_sc_hd__or2_1 _3975_ (.A(_0833_),
    .B(_0846_),
    .X(_0847_));
 sky130_fd_sc_hd__or4_1 _3976_ (.A(\as2650.psl[7] ),
    .B(net327),
    .C(_2584_),
    .D(_0641_),
    .X(_0848_));
 sky130_fd_sc_hd__and3_1 _3977_ (.A(_0645_),
    .B(_0847_),
    .C(_0848_),
    .X(_0849_));
 sky130_fd_sc_hd__a31o_1 _3978_ (.A1(\as2650.psl[7] ),
    .A2(net312),
    .A3(_0644_),
    .B1(_0849_),
    .X(_0850_));
 sky130_fd_sc_hd__mux2_1 _3979_ (.A0(net234),
    .A1(_0850_),
    .S(net146),
    .X(_0851_));
 sky130_fd_sc_hd__nand2_1 _3980_ (.A(net55),
    .B(_0851_),
    .Y(_0852_));
 sky130_fd_sc_hd__o2bb2a_1 _3981_ (.A1_N(net94),
    .A2_N(_0630_),
    .B1(_0467_),
    .B2(_2663_),
    .X(_0853_));
 sky130_fd_sc_hd__a21o_1 _3982_ (.A1(_0852_),
    .A2(_0853_),
    .B1(net115),
    .X(_0854_));
 sky130_fd_sc_hd__o211a_1 _3983_ (.A1(net232),
    .A2(_0775_),
    .B1(_0776_),
    .C1(net81),
    .X(_0855_));
 sky130_fd_sc_hd__o21ba_1 _3984_ (.A1(_0766_),
    .A2(_0772_),
    .B1_N(_0855_),
    .X(_0856_));
 sky130_fd_sc_hd__a22o_1 _3985_ (.A1(_0823_),
    .A2(_0854_),
    .B1(_0856_),
    .B2(net205),
    .X(_0857_));
 sky130_fd_sc_hd__nand2_1 _3986_ (.A(_0813_),
    .B(_0857_),
    .Y(_0858_));
 sky130_fd_sc_hd__o211a_1 _3987_ (.A1(\as2650.psl[7] ),
    .A2(_0813_),
    .B1(_0858_),
    .C1(net320),
    .X(_0069_));
 sky130_fd_sc_hd__or3_4 _3988_ (.A(net219),
    .B(net48),
    .C(net156),
    .X(_0859_));
 sky130_fd_sc_hd__o31ai_4 _3989_ (.A1(net219),
    .A2(_2618_),
    .A3(net155),
    .B1(_0859_),
    .Y(_0860_));
 sky130_fd_sc_hd__mux2_1 _3990_ (.A0(\as2650.stack[1][8] ),
    .A1(_2625_),
    .S(_0860_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _3991_ (.A0(\as2650.stack[1][9] ),
    .A1(_2633_),
    .S(_0860_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _3992_ (.A0(\as2650.stack[1][10] ),
    .A1(_2635_),
    .S(_0860_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _3993_ (.A0(\as2650.stack[1][11] ),
    .A1(_2637_),
    .S(_0860_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _3994_ (.A0(\as2650.stack[1][12] ),
    .A1(_2639_),
    .S(_0860_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _3995_ (.A0(\as2650.stack[1][13] ),
    .A1(_2641_),
    .S(_0860_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _3996_ (.A0(\as2650.stack[1][14] ),
    .A1(_2643_),
    .S(_0860_),
    .X(_0076_));
 sky130_fd_sc_hd__nand2_1 _3997_ (.A(net291),
    .B(_2560_),
    .Y(_0861_));
 sky130_fd_sc_hd__a2111o_4 _3998_ (.A1(_2602_),
    .A2(_0712_),
    .B1(_0861_),
    .C1(_2611_),
    .D1(net164),
    .X(_0862_));
 sky130_fd_sc_hd__and2_1 _3999_ (.A(net308),
    .B(_0862_),
    .X(_0863_));
 sky130_fd_sc_hd__nor2_1 _4000_ (.A(net194),
    .B(_0711_),
    .Y(_0864_));
 sky130_fd_sc_hd__nor2_4 _4001_ (.A(_0712_),
    .B(_0862_),
    .Y(_0865_));
 sky130_fd_sc_hd__and2b_1 _4002_ (.A_N(_0862_),
    .B(_0864_),
    .X(_0866_));
 sky130_fd_sc_hd__a211o_1 _4003_ (.A1(net349),
    .A2(_0865_),
    .B1(_0866_),
    .C1(_0863_),
    .X(_0077_));
 sky130_fd_sc_hd__and2_1 _4004_ (.A(net304),
    .B(_0862_),
    .X(_0867_));
 sky130_fd_sc_hd__a211o_1 _4005_ (.A1(net344),
    .A2(_0865_),
    .B1(_0866_),
    .C1(_0867_),
    .X(_0078_));
 sky130_fd_sc_hd__a22o_1 _4006_ (.A1(net302),
    .A2(_0862_),
    .B1(_0865_),
    .B2(net341),
    .X(_0079_));
 sky130_fd_sc_hd__a211o_1 _4007_ (.A1(net334),
    .A2(_0711_),
    .B1(_0862_),
    .C1(_0864_),
    .X(_0868_));
 sky130_fd_sc_hd__o21a_1 _4008_ (.A1(net300),
    .A2(_0865_),
    .B1(_0868_),
    .X(_0080_));
 sky130_fd_sc_hd__a22o_1 _4009_ (.A1(net299),
    .A2(_0862_),
    .B1(_0865_),
    .B2(net330),
    .X(_0081_));
 sky130_fd_sc_hd__a22o_1 _4010_ (.A1(net297),
    .A2(_0862_),
    .B1(_0865_),
    .B2(net325),
    .X(_0082_));
 sky130_fd_sc_hd__or3_4 _4011_ (.A(net219),
    .B(net48),
    .C(net171),
    .X(_0869_));
 sky130_fd_sc_hd__o31ai_4 _4012_ (.A1(net219),
    .A2(_2618_),
    .A3(net171),
    .B1(_0869_),
    .Y(_0870_));
 sky130_fd_sc_hd__mux2_1 _4013_ (.A0(\as2650.stack[0][8] ),
    .A1(_2625_),
    .S(_0870_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _4014_ (.A0(\as2650.stack[0][9] ),
    .A1(_2633_),
    .S(_0870_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _4015_ (.A0(\as2650.stack[0][10] ),
    .A1(_2635_),
    .S(_0870_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _4016_ (.A0(\as2650.stack[0][11] ),
    .A1(_2637_),
    .S(_0870_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _4017_ (.A0(\as2650.stack[0][12] ),
    .A1(_2639_),
    .S(_0870_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _4018_ (.A0(\as2650.stack[0][13] ),
    .A1(_2641_),
    .S(_0870_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _4019_ (.A0(\as2650.stack[0][14] ),
    .A1(_2643_),
    .S(_0870_),
    .X(_0089_));
 sky130_fd_sc_hd__nor2_2 _4020_ (.A(net293),
    .B(_2805_),
    .Y(_0871_));
 sky130_fd_sc_hd__a31o_4 _4021_ (.A1(net212),
    .A2(net81),
    .A3(_0871_),
    .B1(net348),
    .X(_0872_));
 sky130_fd_sc_hd__nor2_8 _4022_ (.A(net307),
    .B(_0550_),
    .Y(_0873_));
 sky130_fd_sc_hd__nor2_8 _4023_ (.A(_0872_),
    .B(_0873_),
    .Y(_0874_));
 sky130_fd_sc_hd__o21a_2 _4024_ (.A1(_0872_),
    .A2(_0873_),
    .B1(_0558_),
    .X(_0875_));
 sky130_fd_sc_hd__or3_2 _4025_ (.A(_2807_),
    .B(_0514_),
    .C(_0874_),
    .X(_0876_));
 sky130_fd_sc_hd__a22o_1 _4026_ (.A1(_0547_),
    .A2(_0873_),
    .B1(_0874_),
    .B2(\as2650.r123_2[1][0] ),
    .X(_0877_));
 sky130_fd_sc_hd__a31o_1 _4027_ (.A1(net260),
    .A2(net192),
    .A3(_0875_),
    .B1(_0877_),
    .X(_0090_));
 sky130_fd_sc_hd__a22oi_1 _4028_ (.A1(net256),
    .A2(net192),
    .B1(net189),
    .B2(net260),
    .Y(_0878_));
 sky130_fd_sc_hd__and4_1 _4029_ (.A(net256),
    .B(net260),
    .C(net192),
    .D(net189),
    .X(_0879_));
 sky130_fd_sc_hd__or2_1 _4030_ (.A(_0878_),
    .B(_0879_),
    .X(_0880_));
 sky130_fd_sc_hd__a22oi_1 _4031_ (.A1(_0570_),
    .A2(_0873_),
    .B1(_0874_),
    .B2(\as2650.r123_2[1][1] ),
    .Y(_0881_));
 sky130_fd_sc_hd__o21ai_1 _4032_ (.A1(net43),
    .A2(_0880_),
    .B1(_0881_),
    .Y(_0091_));
 sky130_fd_sc_hd__and4_2 _4033_ (.A(net256),
    .B(net261),
    .C(net189),
    .D(net187),
    .X(_0882_));
 sky130_fd_sc_hd__inv_2 _4034_ (.A(_0882_),
    .Y(_0883_));
 sky130_fd_sc_hd__a22o_1 _4035_ (.A1(net256),
    .A2(net189),
    .B1(net187),
    .B2(net261),
    .X(_0884_));
 sky130_fd_sc_hd__nand2_1 _4036_ (.A(net252),
    .B(net191),
    .Y(_0885_));
 sky130_fd_sc_hd__or3b_2 _4037_ (.A(_0882_),
    .B(_0885_),
    .C_N(_0884_),
    .X(_0886_));
 sky130_fd_sc_hd__a21bo_1 _4038_ (.A1(_0883_),
    .A2(_0884_),
    .B1_N(_0885_),
    .X(_0887_));
 sky130_fd_sc_hd__nand3_1 _4039_ (.A(_0879_),
    .B(_0886_),
    .C(_0887_),
    .Y(_0888_));
 sky130_fd_sc_hd__a21o_1 _4040_ (.A1(_0886_),
    .A2(_0887_),
    .B1(_0879_),
    .X(_0889_));
 sky130_fd_sc_hd__nand2_1 _4041_ (.A(_0888_),
    .B(_0889_),
    .Y(_0890_));
 sky130_fd_sc_hd__nor2_1 _4042_ (.A(net43),
    .B(_0890_),
    .Y(_0891_));
 sky130_fd_sc_hd__a221o_1 _4043_ (.A1(_0582_),
    .A2(_0873_),
    .B1(_0874_),
    .B2(\as2650.r123_2[1][2] ),
    .C1(_0891_),
    .X(_0092_));
 sky130_fd_sc_hd__nand2_2 _4044_ (.A(net248),
    .B(net191),
    .Y(_0892_));
 sky130_fd_sc_hd__xnor2_1 _4045_ (.A(_0882_),
    .B(_0892_),
    .Y(_0893_));
 sky130_fd_sc_hd__and4_1 _4046_ (.A(net256),
    .B(net260),
    .C(net187),
    .D(net186),
    .X(_0894_));
 sky130_fd_sc_hd__a22oi_1 _4047_ (.A1(net257),
    .A2(net187),
    .B1(net185),
    .B2(net260),
    .Y(_0895_));
 sky130_fd_sc_hd__a22o_1 _4048_ (.A1(net257),
    .A2(net187),
    .B1(net185),
    .B2(net260),
    .X(_0896_));
 sky130_fd_sc_hd__and4b_1 _4049_ (.A_N(_0894_),
    .B(_0896_),
    .C(net252),
    .D(net189),
    .X(_0897_));
 sky130_fd_sc_hd__o2bb2a_1 _4050_ (.A1_N(net252),
    .A2_N(net189),
    .B1(_0894_),
    .B2(_0895_),
    .X(_0898_));
 sky130_fd_sc_hd__or3b_4 _4051_ (.A(_0897_),
    .B(_0898_),
    .C_N(_0893_),
    .X(_0899_));
 sky130_fd_sc_hd__o21bai_1 _4052_ (.A1(_0897_),
    .A2(_0898_),
    .B1_N(_0893_),
    .Y(_0900_));
 sky130_fd_sc_hd__nand2_1 _4053_ (.A(_0899_),
    .B(_0900_),
    .Y(_0901_));
 sky130_fd_sc_hd__and3_1 _4054_ (.A(_0886_),
    .B(_0888_),
    .C(_0901_),
    .X(_0902_));
 sky130_fd_sc_hd__nor2_1 _4055_ (.A(_0886_),
    .B(_0901_),
    .Y(_0903_));
 sky130_fd_sc_hd__inv_2 _4056_ (.A(_0903_),
    .Y(_0904_));
 sky130_fd_sc_hd__nor2_1 _4057_ (.A(_0888_),
    .B(_0901_),
    .Y(_0905_));
 sky130_fd_sc_hd__inv_2 _4058_ (.A(_0905_),
    .Y(_0906_));
 sky130_fd_sc_hd__or3_1 _4059_ (.A(_0902_),
    .B(_0903_),
    .C(_0905_),
    .X(_0907_));
 sky130_fd_sc_hd__nor2_1 _4060_ (.A(net43),
    .B(_0907_),
    .Y(_0908_));
 sky130_fd_sc_hd__a221o_1 _4061_ (.A1(_0592_),
    .A2(_0873_),
    .B1(_0874_),
    .B2(\as2650.r123_2[1][3] ),
    .C1(_0908_),
    .X(_0093_));
 sky130_fd_sc_hd__nand2_1 _4062_ (.A(net260),
    .B(net184),
    .Y(_0909_));
 sky130_fd_sc_hd__a22o_1 _4063_ (.A1(net253),
    .A2(net187),
    .B1(net186),
    .B2(net256),
    .X(_0910_));
 sky130_fd_sc_hd__and4_2 _4064_ (.A(net252),
    .B(net256),
    .C(net187),
    .D(net185),
    .X(_0911_));
 sky130_fd_sc_hd__nand4_2 _4065_ (.A(net253),
    .B(net256),
    .C(net187),
    .D(net186),
    .Y(_0912_));
 sky130_fd_sc_hd__and4_2 _4066_ (.A(net248),
    .B(net189),
    .C(_0910_),
    .D(_0912_),
    .X(_0913_));
 sky130_fd_sc_hd__nand4_1 _4067_ (.A(net248),
    .B(net189),
    .C(_0910_),
    .D(_0912_),
    .Y(_0914_));
 sky130_fd_sc_hd__a22o_1 _4068_ (.A1(net248),
    .A2(net189),
    .B1(_0910_),
    .B2(_0912_),
    .X(_0915_));
 sky130_fd_sc_hd__or3b_2 _4069_ (.A(_0909_),
    .B(_0913_),
    .C_N(_0915_),
    .X(_0916_));
 sky130_fd_sc_hd__a21bo_1 _4070_ (.A1(_0914_),
    .A2(_0915_),
    .B1_N(_0909_),
    .X(_0917_));
 sky130_fd_sc_hd__a31o_1 _4071_ (.A1(net252),
    .A2(net189),
    .A3(_0896_),
    .B1(_0894_),
    .X(_0918_));
 sky130_fd_sc_hd__nand2_1 _4072_ (.A(net245),
    .B(net191),
    .Y(_0919_));
 sky130_fd_sc_hd__xnor2_1 _4073_ (.A(_0918_),
    .B(_0919_),
    .Y(_0920_));
 sky130_fd_sc_hd__and3_1 _4074_ (.A(_0916_),
    .B(_0917_),
    .C(_0920_),
    .X(_0921_));
 sky130_fd_sc_hd__a21oi_1 _4075_ (.A1(_0916_),
    .A2(_0917_),
    .B1(_0920_),
    .Y(_0922_));
 sky130_fd_sc_hd__or2_2 _4076_ (.A(_0921_),
    .B(_0922_),
    .X(_0923_));
 sky130_fd_sc_hd__o21ai_4 _4077_ (.A1(_0883_),
    .A2(_0892_),
    .B1(_0899_),
    .Y(_0924_));
 sky130_fd_sc_hd__and2b_1 _4078_ (.A_N(_0923_),
    .B(_0924_),
    .X(_0925_));
 sky130_fd_sc_hd__xor2_2 _4079_ (.A(_0923_),
    .B(_0924_),
    .X(_0926_));
 sky130_fd_sc_hd__nor2_1 _4080_ (.A(_0904_),
    .B(_0926_),
    .Y(_0927_));
 sky130_fd_sc_hd__xnor2_1 _4081_ (.A(_0904_),
    .B(_0926_),
    .Y(_0928_));
 sky130_fd_sc_hd__nor2_1 _4082_ (.A(_0906_),
    .B(_0928_),
    .Y(_0929_));
 sky130_fd_sc_hd__and2_1 _4083_ (.A(_0906_),
    .B(_0928_),
    .X(_0930_));
 sky130_fd_sc_hd__nor2_1 _4084_ (.A(_0929_),
    .B(_0930_),
    .Y(_0931_));
 sky130_fd_sc_hd__and2_1 _4085_ (.A(_0875_),
    .B(_0931_),
    .X(_0932_));
 sky130_fd_sc_hd__a221o_1 _4086_ (.A1(_0603_),
    .A2(_0873_),
    .B1(_0874_),
    .B2(\as2650.r123_2[1][4] ),
    .C1(_0932_),
    .X(_0094_));
 sky130_fd_sc_hd__a22oi_2 _4087_ (.A1(net256),
    .A2(net184),
    .B1(net181),
    .B2(net261),
    .Y(_0933_));
 sky130_fd_sc_hd__and4_2 _4088_ (.A(net256),
    .B(net261),
    .C(net184),
    .D(net182),
    .X(_0934_));
 sky130_fd_sc_hd__nor2_2 _4089_ (.A(_0933_),
    .B(_0934_),
    .Y(_0935_));
 sky130_fd_sc_hd__nand2_1 _4090_ (.A(net247),
    .B(net188),
    .Y(_0936_));
 sky130_fd_sc_hd__a22o_2 _4091_ (.A1(net249),
    .A2(net187),
    .B1(net186),
    .B2(net252),
    .X(_0937_));
 sky130_fd_sc_hd__and4_1 _4092_ (.A(net249),
    .B(net252),
    .C(net187),
    .D(net186),
    .X(_0938_));
 sky130_fd_sc_hd__nand4_4 _4093_ (.A(net249),
    .B(net252),
    .C(net188),
    .D(net185),
    .Y(_0939_));
 sky130_fd_sc_hd__and4_1 _4094_ (.A(net245),
    .B(net190),
    .C(_0937_),
    .D(_0939_),
    .X(_0940_));
 sky130_fd_sc_hd__nand4_4 _4095_ (.A(net245),
    .B(net190),
    .C(_0937_),
    .D(_0939_),
    .Y(_0941_));
 sky130_fd_sc_hd__a22o_2 _4096_ (.A1(\as2650.r0[4] ),
    .A2(net190),
    .B1(_0937_),
    .B2(_0939_),
    .X(_0942_));
 sky130_fd_sc_hd__nand3_4 _4097_ (.A(_0935_),
    .B(_0941_),
    .C(_0942_),
    .Y(_0943_));
 sky130_fd_sc_hd__a21o_1 _4098_ (.A1(_0941_),
    .A2(_0942_),
    .B1(_0935_),
    .X(_0944_));
 sky130_fd_sc_hd__and3b_1 _4099_ (.A_N(_0916_),
    .B(_0943_),
    .C(_0944_),
    .X(_0945_));
 sky130_fd_sc_hd__a21bo_2 _4100_ (.A1(_0943_),
    .A2(_0944_),
    .B1_N(_0916_),
    .X(_0946_));
 sky130_fd_sc_hd__nand2b_4 _4101_ (.A_N(_0945_),
    .B(_0946_),
    .Y(_0947_));
 sky130_fd_sc_hd__o211a_2 _4102_ (.A1(_0911_),
    .A2(_0913_),
    .B1(net242),
    .C1(net191),
    .X(_0948_));
 sky130_fd_sc_hd__a211oi_4 _4103_ (.A1(net242),
    .A2(net191),
    .B1(_0911_),
    .C1(_0913_),
    .Y(_0949_));
 sky130_fd_sc_hd__nor2_4 _4104_ (.A(_0948_),
    .B(_0949_),
    .Y(_0950_));
 sky130_fd_sc_hd__xnor2_4 _4105_ (.A(_0947_),
    .B(_0950_),
    .Y(_0951_));
 sky130_fd_sc_hd__a31o_2 _4106_ (.A1(net245),
    .A2(net191),
    .A3(_0918_),
    .B1(_0921_),
    .X(_0952_));
 sky130_fd_sc_hd__and2_1 _4107_ (.A(_0951_),
    .B(_0952_),
    .X(_0953_));
 sky130_fd_sc_hd__xor2_2 _4108_ (.A(_0951_),
    .B(_0952_),
    .X(_0954_));
 sky130_fd_sc_hd__and2_1 _4109_ (.A(_0925_),
    .B(_0954_),
    .X(_0955_));
 sky130_fd_sc_hd__xor2_1 _4110_ (.A(_0925_),
    .B(_0954_),
    .X(_0956_));
 sky130_fd_sc_hd__o21a_1 _4111_ (.A1(_0927_),
    .A2(_0929_),
    .B1(_0956_),
    .X(_0957_));
 sky130_fd_sc_hd__nor3_1 _4112_ (.A(_0927_),
    .B(_0929_),
    .C(_0956_),
    .Y(_0958_));
 sky130_fd_sc_hd__or2_2 _4113_ (.A(_0957_),
    .B(_0958_),
    .X(_0959_));
 sky130_fd_sc_hd__nor2_1 _4114_ (.A(net43),
    .B(_0959_),
    .Y(_0960_));
 sky130_fd_sc_hd__a221o_1 _4115_ (.A1(_0611_),
    .A2(_0873_),
    .B1(_0874_),
    .B2(\as2650.r123_2[1][5] ),
    .C1(_0960_),
    .X(_0095_));
 sky130_fd_sc_hd__a21o_1 _4116_ (.A1(_0946_),
    .A2(_0950_),
    .B1(_0945_),
    .X(_0961_));
 sky130_fd_sc_hd__o211a_1 _4117_ (.A1(_0938_),
    .A2(_0940_),
    .B1(net238),
    .C1(net191),
    .X(_0962_));
 sky130_fd_sc_hd__inv_2 _4118_ (.A(_0962_),
    .Y(_0963_));
 sky130_fd_sc_hd__a211o_1 _4119_ (.A1(net238),
    .A2(net191),
    .B1(_0938_),
    .C1(_0940_),
    .X(_0964_));
 sky130_fd_sc_hd__and2_2 _4120_ (.A(_0963_),
    .B(_0964_),
    .X(_0965_));
 sky130_fd_sc_hd__a22o_2 _4121_ (.A1(net255),
    .A2(net182),
    .B1(net180),
    .B2(net263),
    .X(_0966_));
 sky130_fd_sc_hd__nand4_4 _4122_ (.A(net255),
    .B(net263),
    .C(net182),
    .D(net180),
    .Y(_0967_));
 sky130_fd_sc_hd__a22o_2 _4123_ (.A1(net252),
    .A2(net184),
    .B1(_0966_),
    .B2(_0967_),
    .X(_0968_));
 sky130_fd_sc_hd__nand4_4 _4124_ (.A(net252),
    .B(net184),
    .C(_0966_),
    .D(_0967_),
    .Y(_0969_));
 sky130_fd_sc_hd__nand3_4 _4125_ (.A(_0934_),
    .B(_0968_),
    .C(_0969_),
    .Y(_0970_));
 sky130_fd_sc_hd__a21o_2 _4126_ (.A1(_0968_),
    .A2(_0969_),
    .B1(_0934_),
    .X(_0971_));
 sky130_fd_sc_hd__nand2_2 _4127_ (.A(net241),
    .B(net190),
    .Y(_0972_));
 sky130_fd_sc_hd__a22o_1 _4128_ (.A1(net244),
    .A2(net188),
    .B1(net185),
    .B2(net247),
    .X(_0973_));
 sky130_fd_sc_hd__nand2_2 _4129_ (.A(net244),
    .B(net185),
    .Y(_0974_));
 sky130_fd_sc_hd__nor2_1 _4130_ (.A(_0936_),
    .B(_0974_),
    .Y(_0975_));
 sky130_fd_sc_hd__o21a_2 _4131_ (.A1(_0936_),
    .A2(_0974_),
    .B1(_0973_),
    .X(_0976_));
 sky130_fd_sc_hd__xnor2_4 _4132_ (.A(_0972_),
    .B(_0976_),
    .Y(_0977_));
 sky130_fd_sc_hd__a21oi_4 _4133_ (.A1(_0970_),
    .A2(_0971_),
    .B1(_0977_),
    .Y(_0978_));
 sky130_fd_sc_hd__and3_2 _4134_ (.A(_0970_),
    .B(_0971_),
    .C(_0977_),
    .X(_0979_));
 sky130_fd_sc_hd__or3_4 _4135_ (.A(_0943_),
    .B(_0978_),
    .C(_0979_),
    .X(_0980_));
 sky130_fd_sc_hd__o21ai_4 _4136_ (.A1(_0978_),
    .A2(_0979_),
    .B1(_0943_),
    .Y(_0981_));
 sky130_fd_sc_hd__nand3_4 _4137_ (.A(_0965_),
    .B(_0980_),
    .C(_0981_),
    .Y(_0982_));
 sky130_fd_sc_hd__a21o_1 _4138_ (.A1(_0980_),
    .A2(_0981_),
    .B1(_0965_),
    .X(_0983_));
 sky130_fd_sc_hd__a21o_1 _4139_ (.A1(_0982_),
    .A2(_0983_),
    .B1(_0961_),
    .X(_0984_));
 sky130_fd_sc_hd__nand3_2 _4140_ (.A(_0961_),
    .B(_0982_),
    .C(_0983_),
    .Y(_0985_));
 sky130_fd_sc_hd__a21o_1 _4141_ (.A1(_0984_),
    .A2(_0985_),
    .B1(_0948_),
    .X(_0986_));
 sky130_fd_sc_hd__nand3_2 _4142_ (.A(_0948_),
    .B(_0984_),
    .C(_0985_),
    .Y(_0987_));
 sky130_fd_sc_hd__and3_2 _4143_ (.A(_0953_),
    .B(_0986_),
    .C(_0987_),
    .X(_0988_));
 sky130_fd_sc_hd__nand3_1 _4144_ (.A(_0953_),
    .B(_0986_),
    .C(_0987_),
    .Y(_0989_));
 sky130_fd_sc_hd__a21o_1 _4145_ (.A1(_0986_),
    .A2(_0987_),
    .B1(_0953_),
    .X(_0990_));
 sky130_fd_sc_hd__o211a_2 _4146_ (.A1(_0955_),
    .A2(_0957_),
    .B1(_0989_),
    .C1(_0990_),
    .X(_0991_));
 sky130_fd_sc_hd__a211o_1 _4147_ (.A1(_0989_),
    .A2(_0990_),
    .B1(_0955_),
    .C1(_0957_),
    .X(_0992_));
 sky130_fd_sc_hd__nand2b_1 _4148_ (.A_N(_0991_),
    .B(_0992_),
    .Y(_0993_));
 sky130_fd_sc_hd__nor2_1 _4149_ (.A(_0876_),
    .B(_0993_),
    .Y(_0994_));
 sky130_fd_sc_hd__a221o_1 _4150_ (.A1(_0620_),
    .A2(_0873_),
    .B1(_0874_),
    .B2(\as2650.r123_2[1][6] ),
    .C1(_0994_),
    .X(_0096_));
 sky130_fd_sc_hd__nand2_4 _4151_ (.A(_0980_),
    .B(_0982_),
    .Y(_0995_));
 sky130_fd_sc_hd__a21boi_4 _4152_ (.A1(_0971_),
    .A2(_0977_),
    .B1_N(_0970_),
    .Y(_0996_));
 sky130_fd_sc_hd__nand2_2 _4153_ (.A(net241),
    .B(net188),
    .Y(_0997_));
 sky130_fd_sc_hd__and2_1 _4154_ (.A(_0974_),
    .B(_0997_),
    .X(_0998_));
 sky130_fd_sc_hd__nor2_2 _4155_ (.A(_0974_),
    .B(_0997_),
    .Y(_0999_));
 sky130_fd_sc_hd__and4bb_2 _4156_ (.A_N(_0998_),
    .B_N(_0999_),
    .C(net239),
    .D(net190),
    .X(_1000_));
 sky130_fd_sc_hd__o2bb2a_1 _4157_ (.A1_N(net236),
    .A2_N(net190),
    .B1(_0998_),
    .B2(_0999_),
    .X(_1001_));
 sky130_fd_sc_hd__or2_4 _4158_ (.A(_1000_),
    .B(_1001_),
    .X(_1002_));
 sky130_fd_sc_hd__nand2_4 _4159_ (.A(_0967_),
    .B(_0969_),
    .Y(_1003_));
 sky130_fd_sc_hd__nand2_2 _4160_ (.A(net247),
    .B(net183),
    .Y(_1004_));
 sky130_fd_sc_hd__a22oi_4 _4161_ (.A1(net251),
    .A2(net181),
    .B1(net179),
    .B2(net255),
    .Y(_1005_));
 sky130_fd_sc_hd__and4_2 _4162_ (.A(net251),
    .B(net255),
    .C(net181),
    .D(net179),
    .X(_1006_));
 sky130_fd_sc_hd__nor2_4 _4163_ (.A(_1005_),
    .B(_1006_),
    .Y(_1007_));
 sky130_fd_sc_hd__and3_1 _4164_ (.A(net247),
    .B(net183),
    .C(_1007_),
    .X(_1008_));
 sky130_fd_sc_hd__xnor2_4 _4165_ (.A(_1004_),
    .B(_1007_),
    .Y(_1009_));
 sky130_fd_sc_hd__and2_1 _4166_ (.A(_1003_),
    .B(_1009_),
    .X(_1010_));
 sky130_fd_sc_hd__xnor2_4 _4167_ (.A(_1003_),
    .B(_1009_),
    .Y(_1011_));
 sky130_fd_sc_hd__nor2_1 _4168_ (.A(_1002_),
    .B(_1011_),
    .Y(_1012_));
 sky130_fd_sc_hd__xor2_4 _4169_ (.A(_1002_),
    .B(_1011_),
    .X(_1013_));
 sky130_fd_sc_hd__nand2b_2 _4170_ (.A_N(_0996_),
    .B(_1013_),
    .Y(_1014_));
 sky130_fd_sc_hd__xor2_4 _4171_ (.A(_0996_),
    .B(_1013_),
    .X(_1015_));
 sky130_fd_sc_hd__a31o_2 _4172_ (.A1(net241),
    .A2(net190),
    .A3(_0973_),
    .B1(_0975_),
    .X(_1016_));
 sky130_fd_sc_hd__nand2_1 _4173_ (.A(net234),
    .B(net191),
    .Y(_1017_));
 sky130_fd_sc_hd__and3_2 _4174_ (.A(net234),
    .B(net191),
    .C(_1016_),
    .X(_1018_));
 sky130_fd_sc_hd__xnor2_2 _4175_ (.A(_1016_),
    .B(_1017_),
    .Y(_1019_));
 sky130_fd_sc_hd__and3_4 _4176_ (.A(net259),
    .B(net175),
    .C(_1019_),
    .X(_1020_));
 sky130_fd_sc_hd__a21oi_2 _4177_ (.A1(net259),
    .A2(net175),
    .B1(_1019_),
    .Y(_1021_));
 sky130_fd_sc_hd__nor2_4 _4178_ (.A(_1020_),
    .B(_1021_),
    .Y(_1022_));
 sky130_fd_sc_hd__nand2b_2 _4179_ (.A_N(_1015_),
    .B(_1022_),
    .Y(_1023_));
 sky130_fd_sc_hd__xnor2_4 _4180_ (.A(_1015_),
    .B(_1022_),
    .Y(_1024_));
 sky130_fd_sc_hd__and2_2 _4181_ (.A(_0995_),
    .B(_1024_),
    .X(_1025_));
 sky130_fd_sc_hd__xnor2_4 _4182_ (.A(_0995_),
    .B(_1024_),
    .Y(_1026_));
 sky130_fd_sc_hd__nor2_2 _4183_ (.A(_0963_),
    .B(_1026_),
    .Y(_1027_));
 sky130_fd_sc_hd__xnor2_4 _4184_ (.A(_0963_),
    .B(_1026_),
    .Y(_1028_));
 sky130_fd_sc_hd__and2_2 _4185_ (.A(_0985_),
    .B(_0987_),
    .X(_1029_));
 sky130_fd_sc_hd__or2_2 _4186_ (.A(_1028_),
    .B(_1029_),
    .X(_1030_));
 sky130_fd_sc_hd__xor2_4 _4187_ (.A(_1028_),
    .B(_1029_),
    .X(_1031_));
 sky130_fd_sc_hd__or3_1 _4188_ (.A(_0988_),
    .B(_0991_),
    .C(_1031_),
    .X(_1032_));
 sky130_fd_sc_hd__o21ai_4 _4189_ (.A1(_0988_),
    .A2(_0991_),
    .B1(_1031_),
    .Y(_1033_));
 sky130_fd_sc_hd__nand2_1 _4190_ (.A(_1032_),
    .B(_1033_),
    .Y(_1034_));
 sky130_fd_sc_hd__nor2_1 _4191_ (.A(net43),
    .B(_1034_),
    .Y(_1035_));
 sky130_fd_sc_hd__a221o_1 _4192_ (.A1(_0628_),
    .A2(_0873_),
    .B1(_0874_),
    .B2(\as2650.r123_2[1][7] ),
    .C1(_1035_),
    .X(_0097_));
 sky130_fd_sc_hd__nor2_8 _4193_ (.A(net47),
    .B(_0679_),
    .Y(_1036_));
 sky130_fd_sc_hd__mux2_1 _4194_ (.A0(\as2650.stack[3][0] ),
    .A1(net287),
    .S(_1036_),
    .X(_1037_));
 sky130_fd_sc_hd__mux2_1 _4195_ (.A0(net259),
    .A1(_1037_),
    .S(_0510_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _4196_ (.A0(\as2650.stack[3][1] ),
    .A1(net284),
    .S(_1036_),
    .X(_1038_));
 sky130_fd_sc_hd__mux2_1 _4197_ (.A0(net254),
    .A1(_1038_),
    .S(_0510_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _4198_ (.A0(\as2650.stack[3][2] ),
    .A1(net281),
    .S(_1036_),
    .X(_1039_));
 sky130_fd_sc_hd__mux2_1 _4199_ (.A0(net250),
    .A1(_1039_),
    .S(_0510_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _4200_ (.A0(\as2650.stack[3][3] ),
    .A1(net278),
    .S(_1036_),
    .X(_1040_));
 sky130_fd_sc_hd__mux2_1 _4201_ (.A0(net246),
    .A1(_1040_),
    .S(_0510_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _4202_ (.A0(\as2650.stack[3][4] ),
    .A1(net275),
    .S(_1036_),
    .X(_1041_));
 sky130_fd_sc_hd__mux2_1 _4203_ (.A0(net243),
    .A1(_1041_),
    .S(_0510_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _4204_ (.A0(\as2650.stack[3][5] ),
    .A1(net274),
    .S(_1036_),
    .X(_1042_));
 sky130_fd_sc_hd__mux2_1 _4205_ (.A0(net240),
    .A1(_1042_),
    .S(_0510_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _4206_ (.A0(\as2650.stack[3][6] ),
    .A1(net272),
    .S(_1036_),
    .X(_1043_));
 sky130_fd_sc_hd__mux2_1 _4207_ (.A0(net237),
    .A1(_1043_),
    .S(_0510_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _4208_ (.A0(\as2650.stack[3][7] ),
    .A1(net270),
    .S(_1036_),
    .X(_1044_));
 sky130_fd_sc_hd__mux2_1 _4209_ (.A0(net232),
    .A1(_1044_),
    .S(_0510_),
    .X(_0113_));
 sky130_fd_sc_hd__nor2_4 _4210_ (.A(_0999_),
    .B(_1000_),
    .Y(_1045_));
 sky130_fd_sc_hd__nand2_4 _4211_ (.A(net255),
    .B(net175),
    .Y(_1046_));
 sky130_fd_sc_hd__nor2_4 _4212_ (.A(_1045_),
    .B(_1046_),
    .Y(_1047_));
 sky130_fd_sc_hd__xnor2_4 _4213_ (.A(_1045_),
    .B(_1046_),
    .Y(_1048_));
 sky130_fd_sc_hd__a22o_1 _4214_ (.A1(net239),
    .A2(net188),
    .B1(net185),
    .B2(net242),
    .X(_1049_));
 sky130_fd_sc_hd__nand2_2 _4215_ (.A(net236),
    .B(net185),
    .Y(_1050_));
 sky130_fd_sc_hd__nor2_1 _4216_ (.A(_0997_),
    .B(_1050_),
    .Y(_1051_));
 sky130_fd_sc_hd__o21ai_2 _4217_ (.A1(_0997_),
    .A2(_1050_),
    .B1(_1049_),
    .Y(_1052_));
 sky130_fd_sc_hd__nand2_1 _4218_ (.A(net233),
    .B(net190),
    .Y(_1053_));
 sky130_fd_sc_hd__xnor2_2 _4219_ (.A(_1052_),
    .B(_1053_),
    .Y(_1054_));
 sky130_fd_sc_hd__nand2_1 _4220_ (.A(net244),
    .B(net183),
    .Y(_1055_));
 sky130_fd_sc_hd__and4_1 _4221_ (.A(net248),
    .B(net251),
    .C(net181),
    .D(net179),
    .X(_1056_));
 sky130_fd_sc_hd__a22o_1 _4222_ (.A1(net248),
    .A2(net181),
    .B1(net179),
    .B2(net251),
    .X(_1057_));
 sky130_fd_sc_hd__and2b_1 _4223_ (.A_N(_1056_),
    .B(_1057_),
    .X(_1058_));
 sky130_fd_sc_hd__xnor2_1 _4224_ (.A(_1055_),
    .B(_1058_),
    .Y(_1059_));
 sky130_fd_sc_hd__o21a_2 _4225_ (.A1(_1006_),
    .A2(_1008_),
    .B1(_1059_),
    .X(_1060_));
 sky130_fd_sc_hd__nor3_1 _4226_ (.A(_1006_),
    .B(_1008_),
    .C(_1059_),
    .Y(_1061_));
 sky130_fd_sc_hd__nor2_2 _4227_ (.A(_1060_),
    .B(_1061_),
    .Y(_1062_));
 sky130_fd_sc_hd__and2b_2 _4228_ (.A_N(_1054_),
    .B(_1062_),
    .X(_1063_));
 sky130_fd_sc_hd__xnor2_2 _4229_ (.A(_1054_),
    .B(_1062_),
    .Y(_1064_));
 sky130_fd_sc_hd__o21a_4 _4230_ (.A1(_1010_),
    .A2(_1012_),
    .B1(_1064_),
    .X(_1065_));
 sky130_fd_sc_hd__nor3_2 _4231_ (.A(_1010_),
    .B(_1012_),
    .C(_1064_),
    .Y(_1066_));
 sky130_fd_sc_hd__nor3_4 _4232_ (.A(_1048_),
    .B(_1065_),
    .C(_1066_),
    .Y(_1067_));
 sky130_fd_sc_hd__o21a_2 _4233_ (.A1(_1065_),
    .A2(_1066_),
    .B1(_1048_),
    .X(_1068_));
 sky130_fd_sc_hd__a211o_4 _4234_ (.A1(_1014_),
    .A2(_1023_),
    .B1(_1067_),
    .C1(_1068_),
    .X(_1069_));
 sky130_fd_sc_hd__o211ai_4 _4235_ (.A1(_1067_),
    .A2(_1068_),
    .B1(_1014_),
    .C1(_1023_),
    .Y(_1070_));
 sky130_fd_sc_hd__o211ai_4 _4236_ (.A1(_1018_),
    .A2(_1020_),
    .B1(_1069_),
    .C1(_1070_),
    .Y(_1071_));
 sky130_fd_sc_hd__a211o_2 _4237_ (.A1(_1069_),
    .A2(_1070_),
    .B1(_1018_),
    .C1(_1020_),
    .X(_1072_));
 sky130_fd_sc_hd__o211a_4 _4238_ (.A1(_1025_),
    .A2(_1027_),
    .B1(_1071_),
    .C1(_1072_),
    .X(_1073_));
 sky130_fd_sc_hd__a211oi_4 _4239_ (.A1(_1071_),
    .A2(_1072_),
    .B1(_1025_),
    .C1(_1027_),
    .Y(_1074_));
 sky130_fd_sc_hd__a211oi_4 _4240_ (.A1(_1030_),
    .A2(_1033_),
    .B1(_1073_),
    .C1(_1074_),
    .Y(_1075_));
 sky130_fd_sc_hd__o211a_1 _4241_ (.A1(_1073_),
    .A2(_1074_),
    .B1(_1030_),
    .C1(_1033_),
    .X(_1076_));
 sky130_fd_sc_hd__or2_1 _4242_ (.A(_1075_),
    .B(_1076_),
    .X(_1077_));
 sky130_fd_sc_hd__nor2_1 _4243_ (.A(_0876_),
    .B(_1077_),
    .Y(_1078_));
 sky130_fd_sc_hd__nor2_8 _4244_ (.A(_2584_),
    .B(_0550_),
    .Y(_1079_));
 sky130_fd_sc_hd__nor2_8 _4245_ (.A(_0872_),
    .B(_1079_),
    .Y(_1080_));
 sky130_fd_sc_hd__a221o_1 _4246_ (.A1(_0547_),
    .A2(_1079_),
    .B1(_1080_),
    .B2(\as2650.r123_2[2][0] ),
    .C1(_1078_),
    .X(_0114_));
 sky130_fd_sc_hd__a31o_1 _4247_ (.A1(net233),
    .A2(net190),
    .A3(_1049_),
    .B1(_1051_),
    .X(_1081_));
 sky130_fd_sc_hd__and3_4 _4248_ (.A(net251),
    .B(net174),
    .C(_1081_),
    .X(_1082_));
 sky130_fd_sc_hd__a21oi_1 _4249_ (.A1(net251),
    .A2(net174),
    .B1(_1081_),
    .Y(_1083_));
 sky130_fd_sc_hd__or2_2 _4250_ (.A(_1082_),
    .B(_1083_),
    .X(_1084_));
 sky130_fd_sc_hd__nand2_1 _4251_ (.A(net233),
    .B(net188),
    .Y(_1085_));
 sky130_fd_sc_hd__nand2_2 _4252_ (.A(net233),
    .B(net185),
    .Y(_1086_));
 sky130_fd_sc_hd__and4_1 _4253_ (.A(net233),
    .B(net236),
    .C(net188),
    .D(net185),
    .X(_1087_));
 sky130_fd_sc_hd__a21o_2 _4254_ (.A1(_1050_),
    .A2(_1085_),
    .B1(_1087_),
    .X(_1088_));
 sky130_fd_sc_hd__and4_2 _4255_ (.A(net244),
    .B(net248),
    .C(net181),
    .D(net179),
    .X(_1089_));
 sky130_fd_sc_hd__a22oi_1 _4256_ (.A1(net244),
    .A2(net181),
    .B1(net180),
    .B2(net248),
    .Y(_1090_));
 sky130_fd_sc_hd__nor2_1 _4257_ (.A(_1089_),
    .B(_1090_),
    .Y(_1091_));
 sky130_fd_sc_hd__and3_2 _4258_ (.A(net241),
    .B(net183),
    .C(_1091_),
    .X(_1092_));
 sky130_fd_sc_hd__a21o_1 _4259_ (.A1(net241),
    .A2(net183),
    .B1(_1091_),
    .X(_1093_));
 sky130_fd_sc_hd__and2b_4 _4260_ (.A_N(_1092_),
    .B(_1093_),
    .X(_1094_));
 sky130_fd_sc_hd__a31o_2 _4261_ (.A1(net244),
    .A2(net183),
    .A3(_1057_),
    .B1(_1056_),
    .X(_1095_));
 sky130_fd_sc_hd__xnor2_4 _4262_ (.A(_1094_),
    .B(_1095_),
    .Y(_1096_));
 sky130_fd_sc_hd__xor2_4 _4263_ (.A(_1088_),
    .B(_1096_),
    .X(_1097_));
 sky130_fd_sc_hd__o21a_2 _4264_ (.A1(_1060_),
    .A2(_1063_),
    .B1(_1097_),
    .X(_1098_));
 sky130_fd_sc_hd__nor3_4 _4265_ (.A(_1060_),
    .B(_1063_),
    .C(_1097_),
    .Y(_1099_));
 sky130_fd_sc_hd__nor3_4 _4266_ (.A(_1084_),
    .B(_1098_),
    .C(_1099_),
    .Y(_1100_));
 sky130_fd_sc_hd__o21a_1 _4267_ (.A1(_1098_),
    .A2(_1099_),
    .B1(_1084_),
    .X(_1101_));
 sky130_fd_sc_hd__nor2_2 _4268_ (.A(_1100_),
    .B(_1101_),
    .Y(_1102_));
 sky130_fd_sc_hd__nor2_4 _4269_ (.A(_1065_),
    .B(_1067_),
    .Y(_1103_));
 sky130_fd_sc_hd__or3_1 _4270_ (.A(_1100_),
    .B(_1101_),
    .C(_1103_),
    .X(_1104_));
 sky130_fd_sc_hd__xnor2_4 _4271_ (.A(_1102_),
    .B(_1103_),
    .Y(_1105_));
 sky130_fd_sc_hd__xnor2_4 _4272_ (.A(_1047_),
    .B(_1105_),
    .Y(_1106_));
 sky130_fd_sc_hd__nand2_2 _4273_ (.A(_1069_),
    .B(_1071_),
    .Y(_1107_));
 sky130_fd_sc_hd__nand2b_1 _4274_ (.A_N(_1106_),
    .B(_1107_),
    .Y(_1108_));
 sky130_fd_sc_hd__xnor2_2 _4275_ (.A(_1106_),
    .B(_1107_),
    .Y(_1109_));
 sky130_fd_sc_hd__o21ai_2 _4276_ (.A1(_1073_),
    .A2(_1075_),
    .B1(_1109_),
    .Y(_1110_));
 sky130_fd_sc_hd__or3_1 _4277_ (.A(_1073_),
    .B(_1075_),
    .C(_1109_),
    .X(_1111_));
 sky130_fd_sc_hd__nand2_1 _4278_ (.A(_1110_),
    .B(_1111_),
    .Y(_1112_));
 sky130_fd_sc_hd__nor2_1 _4279_ (.A(net43),
    .B(_1112_),
    .Y(_1113_));
 sky130_fd_sc_hd__a221o_1 _4280_ (.A1(_0570_),
    .A2(_1079_),
    .B1(_1080_),
    .B2(\as2650.r123_2[2][1] ),
    .C1(_1113_),
    .X(_0115_));
 sky130_fd_sc_hd__and3_1 _4281_ (.A(net247),
    .B(net174),
    .C(_1087_),
    .X(_1114_));
 sky130_fd_sc_hd__a21oi_1 _4282_ (.A1(net247),
    .A2(net174),
    .B1(_1087_),
    .Y(_1115_));
 sky130_fd_sc_hd__or2_1 _4283_ (.A(_1114_),
    .B(_1115_),
    .X(_1116_));
 sky130_fd_sc_hd__nand2_1 _4284_ (.A(net241),
    .B(net179),
    .Y(_1117_));
 sky130_fd_sc_hd__and4_2 _4285_ (.A(net241),
    .B(net244),
    .C(net181),
    .D(net179),
    .X(_1118_));
 sky130_fd_sc_hd__a22oi_2 _4286_ (.A1(net241),
    .A2(net181),
    .B1(net179),
    .B2(net244),
    .Y(_1119_));
 sky130_fd_sc_hd__nor2_2 _4287_ (.A(_1118_),
    .B(_1119_),
    .Y(_1120_));
 sky130_fd_sc_hd__nand2_1 _4288_ (.A(net236),
    .B(net183),
    .Y(_1121_));
 sky130_fd_sc_hd__and3_2 _4289_ (.A(net236),
    .B(net183),
    .C(_1120_),
    .X(_1122_));
 sky130_fd_sc_hd__xnor2_2 _4290_ (.A(_1120_),
    .B(_1121_),
    .Y(_1123_));
 sky130_fd_sc_hd__o21ai_4 _4291_ (.A1(_1089_),
    .A2(_1092_),
    .B1(_1123_),
    .Y(_1124_));
 sky130_fd_sc_hd__or3_1 _4292_ (.A(_1089_),
    .B(_1092_),
    .C(_1123_),
    .X(_1125_));
 sky130_fd_sc_hd__nand2_2 _4293_ (.A(_1124_),
    .B(_1125_),
    .Y(_1126_));
 sky130_fd_sc_hd__or2_1 _4294_ (.A(_1086_),
    .B(_1126_),
    .X(_1127_));
 sky130_fd_sc_hd__xor2_2 _4295_ (.A(_1086_),
    .B(_1126_),
    .X(_1128_));
 sky130_fd_sc_hd__a2bb2o_1 _4296_ (.A1_N(_1088_),
    .A2_N(_1096_),
    .B1(_1095_),
    .B2(_1094_),
    .X(_1129_));
 sky130_fd_sc_hd__xnor2_1 _4297_ (.A(_1128_),
    .B(_1129_),
    .Y(_1130_));
 sky130_fd_sc_hd__nor2_1 _4298_ (.A(_1116_),
    .B(_1130_),
    .Y(_1131_));
 sky130_fd_sc_hd__and2_1 _4299_ (.A(_1116_),
    .B(_1130_),
    .X(_1132_));
 sky130_fd_sc_hd__nor2_1 _4300_ (.A(_1131_),
    .B(_1132_),
    .Y(_1133_));
 sky130_fd_sc_hd__o21a_2 _4301_ (.A1(_1098_),
    .A2(_1100_),
    .B1(_1133_),
    .X(_1134_));
 sky130_fd_sc_hd__nor3_2 _4302_ (.A(_1098_),
    .B(_1100_),
    .C(_1133_),
    .Y(_1135_));
 sky130_fd_sc_hd__nor2_4 _4303_ (.A(_1134_),
    .B(_1135_),
    .Y(_1136_));
 sky130_fd_sc_hd__xnor2_4 _4304_ (.A(_1082_),
    .B(_1136_),
    .Y(_1137_));
 sky130_fd_sc_hd__a21bo_1 _4305_ (.A1(_1047_),
    .A2(_1105_),
    .B1_N(_1104_),
    .X(_1138_));
 sky130_fd_sc_hd__nand2b_1 _4306_ (.A_N(_1137_),
    .B(_1138_),
    .Y(_1139_));
 sky130_fd_sc_hd__xor2_2 _4307_ (.A(_1137_),
    .B(_1138_),
    .X(_1140_));
 sky130_fd_sc_hd__a21oi_1 _4308_ (.A1(_1108_),
    .A2(_1110_),
    .B1(_1140_),
    .Y(_1141_));
 sky130_fd_sc_hd__a21o_1 _4309_ (.A1(_1108_),
    .A2(_1110_),
    .B1(_1140_),
    .X(_1142_));
 sky130_fd_sc_hd__and3_1 _4310_ (.A(_1108_),
    .B(_1110_),
    .C(_1140_),
    .X(_1143_));
 sky130_fd_sc_hd__or2_1 _4311_ (.A(_1141_),
    .B(_1143_),
    .X(_1144_));
 sky130_fd_sc_hd__nor2_1 _4312_ (.A(net43),
    .B(_1144_),
    .Y(_1145_));
 sky130_fd_sc_hd__a221o_1 _4313_ (.A1(_0582_),
    .A2(_1079_),
    .B1(_1080_),
    .B2(\as2650.r123_2[2][2] ),
    .C1(_1145_),
    .X(_0116_));
 sky130_fd_sc_hd__nand2_1 _4314_ (.A(net236),
    .B(net181),
    .Y(_1146_));
 sky130_fd_sc_hd__and2_1 _4315_ (.A(_1117_),
    .B(_1146_),
    .X(_1147_));
 sky130_fd_sc_hd__nor2_1 _4316_ (.A(_1117_),
    .B(_1146_),
    .Y(_1148_));
 sky130_fd_sc_hd__nor2_2 _4317_ (.A(_1147_),
    .B(_1148_),
    .Y(_1149_));
 sky130_fd_sc_hd__nand2_1 _4318_ (.A(net233),
    .B(net183),
    .Y(_1150_));
 sky130_fd_sc_hd__xnor2_2 _4319_ (.A(_1149_),
    .B(_1150_),
    .Y(_1151_));
 sky130_fd_sc_hd__o21ai_4 _4320_ (.A1(_1118_),
    .A2(_1122_),
    .B1(_1151_),
    .Y(_1152_));
 sky130_fd_sc_hd__or3_1 _4321_ (.A(_1118_),
    .B(_1122_),
    .C(_1151_),
    .X(_1153_));
 sky130_fd_sc_hd__nand2_1 _4322_ (.A(_1152_),
    .B(_1153_),
    .Y(_1154_));
 sky130_fd_sc_hd__a21oi_2 _4323_ (.A1(_1124_),
    .A2(_1127_),
    .B1(_1154_),
    .Y(_1155_));
 sky130_fd_sc_hd__and3_1 _4324_ (.A(_1124_),
    .B(_1127_),
    .C(_1154_),
    .X(_1156_));
 sky130_fd_sc_hd__or2_1 _4325_ (.A(_1155_),
    .B(_1156_),
    .X(_1157_));
 sky130_fd_sc_hd__nand2_1 _4326_ (.A(net244),
    .B(net174),
    .Y(_1158_));
 sky130_fd_sc_hd__nor2_1 _4327_ (.A(_1157_),
    .B(_1158_),
    .Y(_1159_));
 sky130_fd_sc_hd__xnor2_1 _4328_ (.A(_1157_),
    .B(_1158_),
    .Y(_1160_));
 sky130_fd_sc_hd__a21o_1 _4329_ (.A1(_1128_),
    .A2(_1129_),
    .B1(_1131_),
    .X(_1161_));
 sky130_fd_sc_hd__nand2b_1 _4330_ (.A_N(_1160_),
    .B(_1161_),
    .Y(_1162_));
 sky130_fd_sc_hd__xnor2_1 _4331_ (.A(_1160_),
    .B(_1161_),
    .Y(_1163_));
 sky130_fd_sc_hd__nand2_1 _4332_ (.A(_1114_),
    .B(_1163_),
    .Y(_1164_));
 sky130_fd_sc_hd__or2_1 _4333_ (.A(_1114_),
    .B(_1163_),
    .X(_1165_));
 sky130_fd_sc_hd__and2_1 _4334_ (.A(_1164_),
    .B(_1165_),
    .X(_1166_));
 sky130_fd_sc_hd__a21oi_1 _4335_ (.A1(_1082_),
    .A2(_1136_),
    .B1(_1134_),
    .Y(_1167_));
 sky130_fd_sc_hd__nand2b_1 _4336_ (.A_N(_1167_),
    .B(_1166_),
    .Y(_1168_));
 sky130_fd_sc_hd__nand2b_1 _4337_ (.A_N(_1166_),
    .B(_1167_),
    .Y(_1169_));
 sky130_fd_sc_hd__nand2_1 _4338_ (.A(_1168_),
    .B(_1169_),
    .Y(_1170_));
 sky130_fd_sc_hd__a21o_1 _4339_ (.A1(_1139_),
    .A2(_1142_),
    .B1(_1170_),
    .X(_1171_));
 sky130_fd_sc_hd__nand3_1 _4340_ (.A(_1139_),
    .B(_1142_),
    .C(_1170_),
    .Y(_1172_));
 sky130_fd_sc_hd__nand2_1 _4341_ (.A(_1171_),
    .B(_1172_),
    .Y(_1173_));
 sky130_fd_sc_hd__nor2_1 _4342_ (.A(net43),
    .B(_1173_),
    .Y(_1174_));
 sky130_fd_sc_hd__a221o_1 _4343_ (.A1(_0592_),
    .A2(_1079_),
    .B1(_1080_),
    .B2(\as2650.r123_2[2][3] ),
    .C1(_1174_),
    .X(_0117_));
 sky130_fd_sc_hd__a22o_1 _4344_ (.A1(net234),
    .A2(net182),
    .B1(net179),
    .B2(net236),
    .X(_1175_));
 sky130_fd_sc_hd__nand4_4 _4345_ (.A(net233),
    .B(net236),
    .C(net182),
    .D(net180),
    .Y(_1176_));
 sky130_fd_sc_hd__inv_2 _4346_ (.A(_1176_),
    .Y(_1177_));
 sky130_fd_sc_hd__nand2_1 _4347_ (.A(_1175_),
    .B(_1176_),
    .Y(_1178_));
 sky130_fd_sc_hd__a31o_2 _4348_ (.A1(net233),
    .A2(net183),
    .A3(_1149_),
    .B1(_1148_),
    .X(_1179_));
 sky130_fd_sc_hd__and3_1 _4349_ (.A(_1175_),
    .B(_1176_),
    .C(_1179_),
    .X(_1180_));
 sky130_fd_sc_hd__xnor2_2 _4350_ (.A(_1178_),
    .B(_1179_),
    .Y(_1181_));
 sky130_fd_sc_hd__nand2b_1 _4351_ (.A_N(_1152_),
    .B(_1181_),
    .Y(_1182_));
 sky130_fd_sc_hd__xnor2_2 _4352_ (.A(_1152_),
    .B(_1181_),
    .Y(_1183_));
 sky130_fd_sc_hd__nand3_2 _4353_ (.A(net241),
    .B(net175),
    .C(_1183_),
    .Y(_1184_));
 sky130_fd_sc_hd__a21o_1 _4354_ (.A1(net241),
    .A2(net175),
    .B1(_1183_),
    .X(_1185_));
 sky130_fd_sc_hd__and2_1 _4355_ (.A(_1184_),
    .B(_1185_),
    .X(_1186_));
 sky130_fd_sc_hd__o21ai_2 _4356_ (.A1(_1155_),
    .A2(_1159_),
    .B1(_1186_),
    .Y(_1187_));
 sky130_fd_sc_hd__or3_1 _4357_ (.A(_1155_),
    .B(_1159_),
    .C(_1186_),
    .X(_1188_));
 sky130_fd_sc_hd__nand2_1 _4358_ (.A(_1187_),
    .B(_1188_),
    .Y(_1189_));
 sky130_fd_sc_hd__a21o_1 _4359_ (.A1(_1162_),
    .A2(_1164_),
    .B1(_1189_),
    .X(_1190_));
 sky130_fd_sc_hd__nand3_1 _4360_ (.A(_1162_),
    .B(_1164_),
    .C(_1189_),
    .Y(_1191_));
 sky130_fd_sc_hd__nand2_1 _4361_ (.A(_1190_),
    .B(_1191_),
    .Y(_1192_));
 sky130_fd_sc_hd__a21o_1 _4362_ (.A1(_1168_),
    .A2(_1171_),
    .B1(_1192_),
    .X(_1193_));
 sky130_fd_sc_hd__nand3_1 _4363_ (.A(_1168_),
    .B(_1171_),
    .C(_1192_),
    .Y(_1194_));
 sky130_fd_sc_hd__nand2_1 _4364_ (.A(_1193_),
    .B(_1194_),
    .Y(_1195_));
 sky130_fd_sc_hd__nor2_1 _4365_ (.A(net43),
    .B(_1195_),
    .Y(_1196_));
 sky130_fd_sc_hd__a221o_1 _4366_ (.A1(_0603_),
    .A2(_1079_),
    .B1(_1080_),
    .B2(\as2650.r123_2[2][4] ),
    .C1(_1196_),
    .X(_0118_));
 sky130_fd_sc_hd__and3_1 _4367_ (.A(net233),
    .B(net179),
    .C(_1146_),
    .X(_1197_));
 sky130_fd_sc_hd__xor2_1 _4368_ (.A(_1180_),
    .B(_1197_),
    .X(_1198_));
 sky130_fd_sc_hd__and3_1 _4369_ (.A(net236),
    .B(net174),
    .C(_1198_),
    .X(_1199_));
 sky130_fd_sc_hd__a21oi_1 _4370_ (.A1(net236),
    .A2(net174),
    .B1(_1198_),
    .Y(_1200_));
 sky130_fd_sc_hd__or2_1 _4371_ (.A(_1199_),
    .B(_1200_),
    .X(_1201_));
 sky130_fd_sc_hd__a21oi_2 _4372_ (.A1(_1182_),
    .A2(_1184_),
    .B1(_1201_),
    .Y(_1202_));
 sky130_fd_sc_hd__and3_1 _4373_ (.A(_1182_),
    .B(_1184_),
    .C(_1201_),
    .X(_1203_));
 sky130_fd_sc_hd__or2_1 _4374_ (.A(_1202_),
    .B(_1203_),
    .X(_1204_));
 sky130_fd_sc_hd__or2_1 _4375_ (.A(_1187_),
    .B(_1204_),
    .X(_1205_));
 sky130_fd_sc_hd__nand2_1 _4376_ (.A(_1187_),
    .B(_1204_),
    .Y(_1206_));
 sky130_fd_sc_hd__nand2_1 _4377_ (.A(_1205_),
    .B(_1206_),
    .Y(_1207_));
 sky130_fd_sc_hd__a21o_1 _4378_ (.A1(_1190_),
    .A2(_1193_),
    .B1(_1207_),
    .X(_1208_));
 sky130_fd_sc_hd__nand3_1 _4379_ (.A(_1190_),
    .B(_1193_),
    .C(_1207_),
    .Y(_1209_));
 sky130_fd_sc_hd__nand2_1 _4380_ (.A(_1208_),
    .B(_1209_),
    .Y(_1210_));
 sky130_fd_sc_hd__o2bb2a_1 _4381_ (.A1_N(\as2650.r123_2[2][5] ),
    .A2_N(_1080_),
    .B1(_1210_),
    .B2(net43),
    .X(_1211_));
 sky130_fd_sc_hd__a21bo_1 _4382_ (.A1(_0611_),
    .A2(_1079_),
    .B1_N(_1211_),
    .X(_0119_));
 sky130_fd_sc_hd__a21o_1 _4383_ (.A1(_1180_),
    .A2(_1197_),
    .B1(_1199_),
    .X(_1212_));
 sky130_fd_sc_hd__nand2_1 _4384_ (.A(net233),
    .B(net174),
    .Y(_1213_));
 sky130_fd_sc_hd__mux2_2 _4385_ (.A0(net174),
    .A1(_1213_),
    .S(_1176_),
    .X(_1214_));
 sky130_fd_sc_hd__and2b_1 _4386_ (.A_N(_1214_),
    .B(_1212_),
    .X(_1215_));
 sky130_fd_sc_hd__xnor2_2 _4387_ (.A(_1212_),
    .B(_1214_),
    .Y(_1216_));
 sky130_fd_sc_hd__xnor2_1 _4388_ (.A(_1202_),
    .B(_1216_),
    .Y(_1217_));
 sky130_fd_sc_hd__a21oi_1 _4389_ (.A1(_1205_),
    .A2(_1208_),
    .B1(_1217_),
    .Y(_1218_));
 sky130_fd_sc_hd__and3_1 _4390_ (.A(_1205_),
    .B(_1208_),
    .C(_1217_),
    .X(_1219_));
 sky130_fd_sc_hd__nor2_1 _4391_ (.A(_1218_),
    .B(_1219_),
    .Y(_1220_));
 sky130_fd_sc_hd__a22o_1 _4392_ (.A1(_0620_),
    .A2(_1079_),
    .B1(_1080_),
    .B2(\as2650.r123_2[2][6] ),
    .X(_1221_));
 sky130_fd_sc_hd__a21o_1 _4393_ (.A1(_0875_),
    .A2(_1220_),
    .B1(_1221_),
    .X(_0120_));
 sky130_fd_sc_hd__a21o_1 _4394_ (.A1(_1202_),
    .A2(_1216_),
    .B1(_1215_),
    .X(_1222_));
 sky130_fd_sc_hd__a211o_1 _4395_ (.A1(net174),
    .A2(_1177_),
    .B1(_1218_),
    .C1(_1222_),
    .X(_1223_));
 sky130_fd_sc_hd__a22o_1 _4396_ (.A1(_0628_),
    .A2(_1079_),
    .B1(_1080_),
    .B2(\as2650.r123_2[2][7] ),
    .X(_1224_));
 sky130_fd_sc_hd__a21o_1 _4397_ (.A1(_0875_),
    .A2(_1223_),
    .B1(_1224_),
    .X(_0121_));
 sky130_fd_sc_hd__nor2_8 _4398_ (.A(_2623_),
    .B(_2793_),
    .Y(_1225_));
 sky130_fd_sc_hd__mux2_1 _4399_ (.A0(net286),
    .A1(\as2650.stack[4][0] ),
    .S(_0511_),
    .X(_1226_));
 sky130_fd_sc_hd__mux2_1 _4400_ (.A0(net259),
    .A1(_1226_),
    .S(_0498_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _4401_ (.A0(\as2650.stack[4][1] ),
    .A1(net282),
    .S(_1225_),
    .X(_1227_));
 sky130_fd_sc_hd__mux2_1 _4402_ (.A0(net254),
    .A1(_1227_),
    .S(_0498_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _4403_ (.A0(\as2650.stack[4][2] ),
    .A1(net280),
    .S(_1225_),
    .X(_1228_));
 sky130_fd_sc_hd__mux2_1 _4404_ (.A0(net250),
    .A1(_1228_),
    .S(_0498_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _4405_ (.A0(\as2650.stack[4][3] ),
    .A1(net277),
    .S(_1225_),
    .X(_1229_));
 sky130_fd_sc_hd__mux2_1 _4406_ (.A0(net246),
    .A1(_1229_),
    .S(_0498_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _4407_ (.A0(\as2650.stack[4][4] ),
    .A1(net276),
    .S(_1225_),
    .X(_1230_));
 sky130_fd_sc_hd__mux2_1 _4408_ (.A0(net243),
    .A1(_1230_),
    .S(_0498_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _4409_ (.A0(\as2650.stack[4][5] ),
    .A1(net273),
    .S(_1225_),
    .X(_1231_));
 sky130_fd_sc_hd__mux2_1 _4410_ (.A0(net240),
    .A1(_1231_),
    .S(_0498_),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _4411_ (.A0(\as2650.stack[4][6] ),
    .A1(net271),
    .S(_1225_),
    .X(_1232_));
 sky130_fd_sc_hd__mux2_1 _4412_ (.A0(net237),
    .A1(_1232_),
    .S(_0498_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _4413_ (.A0(\as2650.stack[4][7] ),
    .A1(net269),
    .S(_1225_),
    .X(_1233_));
 sky130_fd_sc_hd__mux2_1 _4414_ (.A0(net232),
    .A1(_1233_),
    .S(_0498_),
    .X(_0129_));
 sky130_fd_sc_hd__nor3_4 _4415_ (.A(net220),
    .B(net168),
    .C(net47),
    .Y(_1234_));
 sky130_fd_sc_hd__mux2_1 _4416_ (.A0(net287),
    .A1(\as2650.stack[2][0] ),
    .S(_0753_),
    .X(_1235_));
 sky130_fd_sc_hd__mux2_1 _4417_ (.A0(net259),
    .A1(_1235_),
    .S(_0680_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _4418_ (.A0(\as2650.stack[2][1] ),
    .A1(net284),
    .S(_1234_),
    .X(_1236_));
 sky130_fd_sc_hd__mux2_1 _4419_ (.A0(net254),
    .A1(_1236_),
    .S(_0680_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _4420_ (.A0(\as2650.stack[2][2] ),
    .A1(net281),
    .S(_1234_),
    .X(_1237_));
 sky130_fd_sc_hd__mux2_1 _4421_ (.A0(net250),
    .A1(_1237_),
    .S(_0680_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _4422_ (.A0(\as2650.stack[2][3] ),
    .A1(net278),
    .S(_1234_),
    .X(_1238_));
 sky130_fd_sc_hd__mux2_1 _4423_ (.A0(net246),
    .A1(_1238_),
    .S(_0680_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _4424_ (.A0(\as2650.stack[2][4] ),
    .A1(net275),
    .S(_1234_),
    .X(_1239_));
 sky130_fd_sc_hd__mux2_1 _4425_ (.A0(net243),
    .A1(_1239_),
    .S(_0680_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _4426_ (.A0(\as2650.stack[2][5] ),
    .A1(net274),
    .S(_1234_),
    .X(_1240_));
 sky130_fd_sc_hd__mux2_1 _4427_ (.A0(net240),
    .A1(_1240_),
    .S(_0680_),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _4428_ (.A0(\as2650.stack[2][6] ),
    .A1(net272),
    .S(_1234_),
    .X(_1241_));
 sky130_fd_sc_hd__mux2_1 _4429_ (.A0(net237),
    .A1(_1241_),
    .S(_0680_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _4430_ (.A0(\as2650.stack[2][7] ),
    .A1(net270),
    .S(_1234_),
    .X(_1242_));
 sky130_fd_sc_hd__mux2_1 _4431_ (.A0(net232),
    .A1(_1242_),
    .S(_0680_),
    .X(_0137_));
 sky130_fd_sc_hd__nor3_4 _4432_ (.A(net220),
    .B(net47),
    .C(net157),
    .Y(_1243_));
 sky130_fd_sc_hd__mux2_1 _4433_ (.A0(\as2650.stack[1][0] ),
    .A1(net287),
    .S(_1243_),
    .X(_1244_));
 sky130_fd_sc_hd__mux2_1 _4434_ (.A0(net259),
    .A1(_1244_),
    .S(_0752_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _4435_ (.A0(\as2650.stack[1][1] ),
    .A1(net284),
    .S(_1243_),
    .X(_1245_));
 sky130_fd_sc_hd__mux2_1 _4436_ (.A0(net254),
    .A1(_1245_),
    .S(_0752_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _4437_ (.A0(\as2650.stack[1][2] ),
    .A1(net281),
    .S(_1243_),
    .X(_1246_));
 sky130_fd_sc_hd__mux2_1 _4438_ (.A0(net250),
    .A1(_1246_),
    .S(_0752_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _4439_ (.A0(\as2650.stack[1][3] ),
    .A1(net278),
    .S(_1243_),
    .X(_1247_));
 sky130_fd_sc_hd__mux2_1 _4440_ (.A0(net247),
    .A1(_1247_),
    .S(_0752_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _4441_ (.A0(\as2650.stack[1][4] ),
    .A1(net275),
    .S(_1243_),
    .X(_1248_));
 sky130_fd_sc_hd__mux2_1 _4442_ (.A0(net243),
    .A1(_1248_),
    .S(_0752_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _4443_ (.A0(\as2650.stack[1][5] ),
    .A1(net274),
    .S(_1243_),
    .X(_1249_));
 sky130_fd_sc_hd__mux2_1 _4444_ (.A0(net240),
    .A1(_1249_),
    .S(_0752_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _4445_ (.A0(\as2650.stack[1][6] ),
    .A1(net272),
    .S(_1243_),
    .X(_1250_));
 sky130_fd_sc_hd__mux2_1 _4446_ (.A0(net237),
    .A1(_1250_),
    .S(_0752_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _4447_ (.A0(\as2650.stack[1][7] ),
    .A1(net270),
    .S(_1243_),
    .X(_1251_));
 sky130_fd_sc_hd__mux2_1 _4448_ (.A0(net232),
    .A1(_1251_),
    .S(_0752_),
    .X(_0145_));
 sky130_fd_sc_hd__o21ai_1 _4449_ (.A1(_0687_),
    .A2(_0690_),
    .B1(_2607_),
    .Y(_1252_));
 sky130_fd_sc_hd__a31o_1 _4450_ (.A1(net139),
    .A2(net162),
    .A3(_2627_),
    .B1(net137),
    .X(_1253_));
 sky130_fd_sc_hd__a21oi_1 _4451_ (.A1(net73),
    .A2(net54),
    .B1(_1253_),
    .Y(_1254_));
 sky130_fd_sc_hd__nor2_4 _4452_ (.A(net134),
    .B(net161),
    .Y(_1255_));
 sky130_fd_sc_hd__nand2_1 _4453_ (.A(_2537_),
    .B(_2594_),
    .Y(_1256_));
 sky130_fd_sc_hd__nor2_1 _4454_ (.A(net135),
    .B(net161),
    .Y(_1257_));
 sky130_fd_sc_hd__a32o_1 _4455_ (.A1(net124),
    .A2(_0709_),
    .A3(_1257_),
    .B1(_1256_),
    .B2(_1255_),
    .X(_1258_));
 sky130_fd_sc_hd__and4_1 _4456_ (.A(net225),
    .B(net141),
    .C(_2603_),
    .D(_1258_),
    .X(_1259_));
 sky130_fd_sc_hd__a211oi_4 _4457_ (.A1(net203),
    .A2(net87),
    .B1(_0713_),
    .C1(net90),
    .Y(_1260_));
 sky130_fd_sc_hd__a21oi_4 _4458_ (.A1(net303),
    .A2(net141),
    .B1(_2590_),
    .Y(_1261_));
 sky130_fd_sc_hd__or3b_1 _4459_ (.A(_2561_),
    .B(_0731_),
    .C_N(_1260_),
    .X(_1262_));
 sky130_fd_sc_hd__or4b_1 _4460_ (.A(_1254_),
    .B(_1262_),
    .C(_1259_),
    .D_N(_2595_),
    .X(_1263_));
 sky130_fd_sc_hd__a211o_4 _4461_ (.A1(net54),
    .A2(_1252_),
    .B1(_1261_),
    .C1(_1263_),
    .X(_1264_));
 sky130_fd_sc_hd__mux2_1 _4462_ (.A0(net349),
    .A1(net296),
    .S(_1264_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _4463_ (.A0(net344),
    .A1(net295),
    .S(_1264_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _4464_ (.A0(net341),
    .A1(\as2650.addr_buff[2] ),
    .S(_1264_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _4465_ (.A0(net338),
    .A1(\as2650.addr_buff[3] ),
    .S(_1264_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _4466_ (.A0(net335),
    .A1(\as2650.addr_buff[4] ),
    .S(_1264_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _4467_ (.A0(net332),
    .A1(\as2650.addr_buff[5] ),
    .S(_1264_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _4468_ (.A0(net331),
    .A1(\as2650.addr_buff[6] ),
    .S(_1264_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _4469_ (.A0(net326),
    .A1(\as2650.addr_buff[7] ),
    .S(_1264_),
    .X(_0161_));
 sky130_fd_sc_hd__and3b_4 _4470_ (.A_N(net47),
    .B(net172),
    .C(_2529_),
    .X(_1265_));
 sky130_fd_sc_hd__mux2_1 _4471_ (.A0(\as2650.stack[0][0] ),
    .A1(net287),
    .S(_1265_),
    .X(_1266_));
 sky130_fd_sc_hd__mux2_1 _4472_ (.A0(net259),
    .A1(_1266_),
    .S(_0859_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _4473_ (.A0(\as2650.stack[0][1] ),
    .A1(net284),
    .S(_1265_),
    .X(_1267_));
 sky130_fd_sc_hd__mux2_1 _4474_ (.A0(net254),
    .A1(_1267_),
    .S(_0859_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _4475_ (.A0(\as2650.stack[0][2] ),
    .A1(net281),
    .S(_1265_),
    .X(_1268_));
 sky130_fd_sc_hd__mux2_1 _4476_ (.A0(net250),
    .A1(_1268_),
    .S(_0859_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _4477_ (.A0(\as2650.stack[0][3] ),
    .A1(net278),
    .S(_1265_),
    .X(_1269_));
 sky130_fd_sc_hd__mux2_1 _4478_ (.A0(net247),
    .A1(_1269_),
    .S(_0859_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _4479_ (.A0(\as2650.stack[0][4] ),
    .A1(net275),
    .S(_1265_),
    .X(_1270_));
 sky130_fd_sc_hd__mux2_1 _4480_ (.A0(net243),
    .A1(_1270_),
    .S(_0859_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _4481_ (.A0(\as2650.stack[0][5] ),
    .A1(net274),
    .S(_1265_),
    .X(_1271_));
 sky130_fd_sc_hd__mux2_1 _4482_ (.A0(net240),
    .A1(_1271_),
    .S(_0859_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _4483_ (.A0(\as2650.stack[0][6] ),
    .A1(net272),
    .S(_1265_),
    .X(_1272_));
 sky130_fd_sc_hd__mux2_1 _4484_ (.A0(net237),
    .A1(_1272_),
    .S(_0859_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _4485_ (.A0(\as2650.stack[0][7] ),
    .A1(net270),
    .S(_1265_),
    .X(_1273_));
 sky130_fd_sc_hd__mux2_1 _4486_ (.A0(net232),
    .A1(_1273_),
    .S(_0859_),
    .X(_0169_));
 sky130_fd_sc_hd__o31a_1 _4487_ (.A1(net150),
    .A2(net131),
    .A3(net61),
    .B1(net141),
    .X(_1274_));
 sky130_fd_sc_hd__nor2_2 _4488_ (.A(net293),
    .B(net162),
    .Y(_1275_));
 sky130_fd_sc_hd__and4_1 _4489_ (.A(_2682_),
    .B(net92),
    .C(_0714_),
    .D(_1275_),
    .X(_1276_));
 sky130_fd_sc_hd__or4_2 _4490_ (.A(net208),
    .B(net230),
    .C(_2652_),
    .D(_0710_),
    .X(_1277_));
 sky130_fd_sc_hd__and3_1 _4491_ (.A(_0729_),
    .B(_1276_),
    .C(_1277_),
    .X(_1278_));
 sky130_fd_sc_hd__o221a_4 _4492_ (.A1(_2606_),
    .A2(_0799_),
    .B1(_1274_),
    .B2(_0715_),
    .C1(_1278_),
    .X(_1279_));
 sky130_fd_sc_hd__o211ai_4 _4493_ (.A1(net203),
    .A2(_2610_),
    .B1(_0710_),
    .C1(_1279_),
    .Y(_1280_));
 sky130_fd_sc_hd__o211a_1 _4494_ (.A1(net27),
    .A2(_1279_),
    .B1(_1280_),
    .C1(net316),
    .X(_0170_));
 sky130_fd_sc_hd__and3_1 _4495_ (.A(net79),
    .B(net92),
    .C(_0790_),
    .X(_1281_));
 sky130_fd_sc_hd__and3_1 _4496_ (.A(_2535_),
    .B(_0712_),
    .C(_1281_),
    .X(_1282_));
 sky130_fd_sc_hd__mux2_1 _4497_ (.A0(net29),
    .A1(net299),
    .S(_1282_),
    .X(_1283_));
 sky130_fd_sc_hd__and2_1 _4498_ (.A(net316),
    .B(_1283_),
    .X(_0171_));
 sky130_fd_sc_hd__nor2_1 _4499_ (.A(_0696_),
    .B(_0718_),
    .Y(_1284_));
 sky130_fd_sc_hd__a31o_1 _4500_ (.A1(net164),
    .A2(net126),
    .A3(_0791_),
    .B1(_1284_),
    .X(_1285_));
 sky130_fd_sc_hd__a31o_1 _4501_ (.A1(net297),
    .A2(_2612_),
    .A3(_0790_),
    .B1(_1285_),
    .X(_1286_));
 sky130_fd_sc_hd__a211o_1 _4502_ (.A1(net148),
    .A2(net115),
    .B1(net151),
    .C1(_0727_),
    .X(_1287_));
 sky130_fd_sc_hd__a2111o_2 _4503_ (.A1(_0697_),
    .A2(_1287_),
    .B1(_0711_),
    .C1(net292),
    .D1(_1286_),
    .X(_1288_));
 sky130_fd_sc_hd__nor2_1 _4504_ (.A(net163),
    .B(_1288_),
    .Y(_1289_));
 sky130_fd_sc_hd__a211o_1 _4505_ (.A1(net28),
    .A2(_1288_),
    .B1(_1289_),
    .C1(net347),
    .X(_0172_));
 sky130_fd_sc_hd__o31a_1 _4506_ (.A1(net65),
    .A2(_0782_),
    .A3(_0796_),
    .B1(net79),
    .X(_1290_));
 sky130_fd_sc_hd__nand2_1 _4507_ (.A(net81),
    .B(_0802_),
    .Y(_1291_));
 sky130_fd_sc_hd__or2_2 _4508_ (.A(_0797_),
    .B(_1291_),
    .X(_1292_));
 sky130_fd_sc_hd__o22a_1 _4509_ (.A1(net146),
    .A2(_0654_),
    .B1(_0696_),
    .B2(_2655_),
    .X(_1293_));
 sky130_fd_sc_hd__o31ai_4 _4510_ (.A1(net226),
    .A2(_0696_),
    .A3(_1292_),
    .B1(_1293_),
    .Y(_1294_));
 sky130_fd_sc_hd__a21oi_4 _4511_ (.A1(_2774_),
    .A2(_0660_),
    .B1(_2810_),
    .Y(_1295_));
 sky130_fd_sc_hd__inv_2 _4512_ (.A(_1295_),
    .Y(_1296_));
 sky130_fd_sc_hd__and3_1 _4513_ (.A(_2662_),
    .B(net153),
    .C(_0697_),
    .X(_1297_));
 sky130_fd_sc_hd__nor2_1 _4514_ (.A(_2805_),
    .B(_0805_),
    .Y(_1298_));
 sky130_fd_sc_hd__or2_1 _4515_ (.A(_2805_),
    .B(_0805_),
    .X(_1299_));
 sky130_fd_sc_hd__or4_1 _4516_ (.A(_0711_),
    .B(_1284_),
    .C(_1297_),
    .D(_1298_),
    .X(_1300_));
 sky130_fd_sc_hd__or4_1 _4517_ (.A(_1290_),
    .B(_1294_),
    .C(_1296_),
    .D(_1300_),
    .X(_1301_));
 sky130_fd_sc_hd__o21ai_1 _4518_ (.A1(net230),
    .A2(_2679_),
    .B1(_0710_),
    .Y(_1302_));
 sky130_fd_sc_hd__a21o_1 _4519_ (.A1(_0697_),
    .A2(_1302_),
    .B1(_0716_),
    .X(_1303_));
 sky130_fd_sc_hd__a21o_1 _4520_ (.A1(_0697_),
    .A2(_1259_),
    .B1(_1303_),
    .X(_1304_));
 sky130_fd_sc_hd__nor2_1 _4521_ (.A(net163),
    .B(_2668_),
    .Y(_1305_));
 sky130_fd_sc_hd__or3_4 _4522_ (.A(net80),
    .B(_0690_),
    .C(_0711_),
    .X(_1306_));
 sky130_fd_sc_hd__nor2_1 _4523_ (.A(_0701_),
    .B(_1306_),
    .Y(_1307_));
 sky130_fd_sc_hd__or3_1 _4524_ (.A(_0691_),
    .B(_0701_),
    .C(_1306_),
    .X(_1308_));
 sky130_fd_sc_hd__nor2_1 _4525_ (.A(net202),
    .B(net89),
    .Y(_1309_));
 sky130_fd_sc_hd__nand2_4 _4526_ (.A(net225),
    .B(net88),
    .Y(_1310_));
 sky130_fd_sc_hd__a311o_1 _4527_ (.A1(net222),
    .A2(net164),
    .A3(net121),
    .B1(_0713_),
    .C1(net292),
    .X(_1311_));
 sky130_fd_sc_hd__o32a_2 _4528_ (.A1(net205),
    .A2(_2586_),
    .A3(_0666_),
    .B1(_0667_),
    .B2(_2572_),
    .X(_1312_));
 sky130_fd_sc_hd__nand2_2 _4529_ (.A(net230),
    .B(_2590_),
    .Y(_1313_));
 sky130_fd_sc_hd__or3_2 _4530_ (.A(net141),
    .B(_1312_),
    .C(_1313_),
    .X(_1314_));
 sky130_fd_sc_hd__and3b_1 _4531_ (.A_N(_1311_),
    .B(_1314_),
    .C(_2696_),
    .X(_1315_));
 sky130_fd_sc_hd__nand2_2 _4532_ (.A(_1308_),
    .B(_1315_),
    .Y(_1316_));
 sky130_fd_sc_hd__or3_1 _4533_ (.A(net204),
    .B(_0635_),
    .C(_0793_),
    .X(_1317_));
 sky130_fd_sc_hd__a41o_2 _4534_ (.A1(net225),
    .A2(_0634_),
    .A3(_0697_),
    .A4(_0794_),
    .B1(_2580_),
    .X(_1318_));
 sky130_fd_sc_hd__or4_4 _4535_ (.A(_1301_),
    .B(_1304_),
    .C(_1316_),
    .D(_1318_),
    .X(_1319_));
 sky130_fd_sc_hd__or4_1 _4536_ (.A(_2709_),
    .B(_2822_),
    .C(_2870_),
    .D(_2914_),
    .X(_1320_));
 sky130_fd_sc_hd__or4b_2 _4537_ (.A(_0321_),
    .B(_0426_),
    .C(_1320_),
    .D_N(_0381_),
    .X(_1321_));
 sky130_fd_sc_hd__nor2_2 _4538_ (.A(_0463_),
    .B(_1321_),
    .Y(_1322_));
 sky130_fd_sc_hd__or3_4 _4539_ (.A(_2649_),
    .B(_0463_),
    .C(_1321_),
    .X(_1323_));
 sky130_fd_sc_hd__or3_4 _4540_ (.A(net137),
    .B(_2690_),
    .C(_1323_),
    .X(_1324_));
 sky130_fd_sc_hd__nand2b_2 _4541_ (.A_N(_0803_),
    .B(_1324_),
    .Y(_1325_));
 sky130_fd_sc_hd__nor2_1 _4542_ (.A(_1319_),
    .B(net42),
    .Y(_1326_));
 sky130_fd_sc_hd__nand2_2 _4543_ (.A(net286),
    .B(net349),
    .Y(_1327_));
 sky130_fd_sc_hd__or2_1 _4544_ (.A(net286),
    .B(net349),
    .X(_1328_));
 sky130_fd_sc_hd__nand2_2 _4545_ (.A(_1327_),
    .B(_1328_),
    .Y(_1329_));
 sky130_fd_sc_hd__mux2_1 _4546_ (.A0(_2542_),
    .A1(_1329_),
    .S(net323),
    .X(_1330_));
 sky130_fd_sc_hd__o211a_1 _4547_ (.A1(net137),
    .A2(net161),
    .B1(net208),
    .C1(net140),
    .X(_1331_));
 sky130_fd_sc_hd__nand2_1 _4548_ (.A(net349),
    .B(net127),
    .Y(_1332_));
 sky130_fd_sc_hd__nor2_4 _4549_ (.A(net206),
    .B(net76),
    .Y(_1333_));
 sky130_fd_sc_hd__nor2_4 _4550_ (.A(net120),
    .B(net161),
    .Y(_1334_));
 sky130_fd_sc_hd__nor2_4 _4551_ (.A(net208),
    .B(_2610_),
    .Y(_1335_));
 sky130_fd_sc_hd__nand2_1 _4552_ (.A(net302),
    .B(net161),
    .Y(_1336_));
 sky130_fd_sc_hd__nor2_1 _4553_ (.A(net76),
    .B(_1335_),
    .Y(_1337_));
 sky130_fd_sc_hd__nand2_2 _4554_ (.A(net140),
    .B(net84),
    .Y(_1338_));
 sky130_fd_sc_hd__nor2_1 _4555_ (.A(net206),
    .B(_1338_),
    .Y(_1339_));
 sky130_fd_sc_hd__mux2_1 _4556_ (.A0(net127),
    .A1(_2616_),
    .S(net37),
    .X(_1340_));
 sky130_fd_sc_hd__o211a_1 _4557_ (.A1(_2615_),
    .A2(_1332_),
    .B1(_1334_),
    .C1(_1340_),
    .X(_1341_));
 sky130_fd_sc_hd__or2_4 _4558_ (.A(net120),
    .B(net116),
    .X(_1342_));
 sky130_fd_sc_hd__a21o_1 _4559_ (.A1(_1330_),
    .A2(_1342_),
    .B1(_1341_),
    .X(_1343_));
 sky130_fd_sc_hd__o2bb2a_1 _4560_ (.A1_N(net50),
    .A2_N(_1343_),
    .B1(_1339_),
    .B2(net285),
    .X(_1344_));
 sky130_fd_sc_hd__nand2_1 _4561_ (.A(_2687_),
    .B(_2746_),
    .Y(_1345_));
 sky130_fd_sc_hd__xor2_1 _4562_ (.A(net350),
    .B(_1345_),
    .X(_1346_));
 sky130_fd_sc_hd__nor2_8 _4563_ (.A(\as2650.addr_buff[7] ),
    .B(_2675_),
    .Y(_1347_));
 sky130_fd_sc_hd__nand2_1 _4564_ (.A(_2736_),
    .B(_1347_),
    .Y(_1348_));
 sky130_fd_sc_hd__xor2_1 _4565_ (.A(net350),
    .B(_1348_),
    .X(_1349_));
 sky130_fd_sc_hd__a22o_2 _4566_ (.A1(_0686_),
    .A2(_1346_),
    .B1(_1349_),
    .B2(net74),
    .X(_1350_));
 sky130_fd_sc_hd__nor2_1 _4567_ (.A(net85),
    .B(_1329_),
    .Y(_1351_));
 sky130_fd_sc_hd__a221o_1 _4568_ (.A1(net37),
    .A2(net91),
    .B1(_0688_),
    .B2(_1350_),
    .C1(_1351_),
    .X(_1352_));
 sky130_fd_sc_hd__o2bb2a_2 _4569_ (.A1_N(net225),
    .A2_N(_1344_),
    .B1(_1352_),
    .B2(_0694_),
    .X(_1353_));
 sky130_fd_sc_hd__o221ai_4 _4570_ (.A1(_2534_),
    .A2(net51),
    .B1(_1353_),
    .B2(net89),
    .C1(net39),
    .Y(_1354_));
 sky130_fd_sc_hd__o211a_1 _4571_ (.A1(net37),
    .A2(net39),
    .B1(_1354_),
    .C1(net314),
    .X(_0173_));
 sky130_fd_sc_hd__and2_1 _4572_ (.A(net345),
    .B(_2838_),
    .X(_1355_));
 sky130_fd_sc_hd__or2_1 _4573_ (.A(net345),
    .B(_2838_),
    .X(_1356_));
 sky130_fd_sc_hd__and2b_1 _4574_ (.A_N(_1355_),
    .B(_1356_),
    .X(_1357_));
 sky130_fd_sc_hd__and2_1 _4575_ (.A(net350),
    .B(_2746_),
    .X(_1358_));
 sky130_fd_sc_hd__xor2_1 _4576_ (.A(_1357_),
    .B(_1358_),
    .X(_1359_));
 sky130_fd_sc_hd__nand2_1 _4577_ (.A(_2550_),
    .B(net176),
    .Y(_1360_));
 sky130_fd_sc_hd__o211a_1 _4578_ (.A1(net176),
    .A2(_1359_),
    .B1(_1360_),
    .C1(_0686_),
    .X(_1361_));
 sky130_fd_sc_hd__nor2_4 _4579_ (.A(net72),
    .B(_1347_),
    .Y(_1362_));
 sky130_fd_sc_hd__and2_1 _4580_ (.A(net345),
    .B(_2834_),
    .X(_1363_));
 sky130_fd_sc_hd__nand2_1 _4581_ (.A(net345),
    .B(_2834_),
    .Y(_1364_));
 sky130_fd_sc_hd__or2_1 _4582_ (.A(net345),
    .B(_2834_),
    .X(_1365_));
 sky130_fd_sc_hd__and2_1 _4583_ (.A(net350),
    .B(_2736_),
    .X(_1366_));
 sky130_fd_sc_hd__and3_1 _4584_ (.A(_1364_),
    .B(_1365_),
    .C(_1366_),
    .X(_1367_));
 sky130_fd_sc_hd__a21oi_1 _4585_ (.A1(_1364_),
    .A2(_1365_),
    .B1(_1366_),
    .Y(_1368_));
 sky130_fd_sc_hd__nor2_4 _4586_ (.A(_2673_),
    .B(_2675_),
    .Y(_1369_));
 sky130_fd_sc_hd__nor2_1 _4587_ (.A(_1367_),
    .B(_1368_),
    .Y(_1370_));
 sky130_fd_sc_hd__a221o_4 _4588_ (.A1(net345),
    .A2(_1362_),
    .B1(_1369_),
    .B2(_1370_),
    .C1(_1361_),
    .X(_1371_));
 sky130_fd_sc_hd__and2_1 _4589_ (.A(net282),
    .B(net344),
    .X(_1372_));
 sky130_fd_sc_hd__nand2_1 _4590_ (.A(net282),
    .B(net344),
    .Y(_1373_));
 sky130_fd_sc_hd__nor2_1 _4591_ (.A(net282),
    .B(net344),
    .Y(_1374_));
 sky130_fd_sc_hd__nor2_2 _4592_ (.A(_1372_),
    .B(_1374_),
    .Y(_1375_));
 sky130_fd_sc_hd__nand2_1 _4593_ (.A(_1328_),
    .B(_1375_),
    .Y(_1376_));
 sky130_fd_sc_hd__or2_1 _4594_ (.A(_1328_),
    .B(_1375_),
    .X(_1377_));
 sky130_fd_sc_hd__xor2_1 _4595_ (.A(net38),
    .B(net37),
    .X(_1378_));
 sky130_fd_sc_hd__a31o_1 _4596_ (.A1(net86),
    .A2(_1376_),
    .A3(_1377_),
    .B1(_0694_),
    .X(_1379_));
 sky130_fd_sc_hd__a22o_1 _4597_ (.A1(_0688_),
    .A2(_1371_),
    .B1(_1378_),
    .B2(net91),
    .X(_1380_));
 sky130_fd_sc_hd__or2_1 _4598_ (.A(_1379_),
    .B(_1380_),
    .X(_1381_));
 sky130_fd_sc_hd__and2_4 _4599_ (.A(net294),
    .B(net128),
    .X(_1382_));
 sky130_fd_sc_hd__nand2_8 _4600_ (.A(net294),
    .B(net128),
    .Y(_1383_));
 sky130_fd_sc_hd__nor2_1 _4601_ (.A(net149),
    .B(net120),
    .Y(_1384_));
 sky130_fd_sc_hd__o221a_1 _4602_ (.A1(net38),
    .A2(_2616_),
    .B1(_1378_),
    .B2(net127),
    .C1(_1384_),
    .X(_1385_));
 sky130_fd_sc_hd__o21a_1 _4603_ (.A1(net344),
    .A2(_1383_),
    .B1(_1385_),
    .X(_1386_));
 sky130_fd_sc_hd__xnor2_2 _4604_ (.A(_1327_),
    .B(_1375_),
    .Y(_1387_));
 sky130_fd_sc_hd__mux2_1 _4605_ (.A0(net38),
    .A1(_1387_),
    .S(net322),
    .X(_1388_));
 sky130_fd_sc_hd__a221o_1 _4606_ (.A1(net283),
    .A2(_1338_),
    .B1(_1388_),
    .B2(_1331_),
    .C1(net193),
    .X(_1389_));
 sky130_fd_sc_hd__and2_2 _4607_ (.A(net140),
    .B(_1342_),
    .X(_1390_));
 sky130_fd_sc_hd__or2_1 _4608_ (.A(_1386_),
    .B(_1389_),
    .X(_1391_));
 sky130_fd_sc_hd__o211a_1 _4609_ (.A1(net283),
    .A2(net151),
    .B1(_1381_),
    .C1(_1391_),
    .X(_1392_));
 sky130_fd_sc_hd__o22a_1 _4610_ (.A1(net283),
    .A2(net51),
    .B1(_1392_),
    .B2(net89),
    .X(_1393_));
 sky130_fd_sc_hd__or2_1 _4611_ (.A(net38),
    .B(net39),
    .X(_1394_));
 sky130_fd_sc_hd__o311a_1 _4612_ (.A1(_1319_),
    .A2(net42),
    .A3(_1393_),
    .B1(_1394_),
    .C1(net314),
    .X(_0174_));
 sky130_fd_sc_hd__a21oi_1 _4613_ (.A1(_1356_),
    .A2(_1358_),
    .B1(_1355_),
    .Y(_1395_));
 sky130_fd_sc_hd__or2_4 _4614_ (.A(net342),
    .B(_2886_),
    .X(_1396_));
 sky130_fd_sc_hd__nand2_1 _4615_ (.A(net342),
    .B(_2886_),
    .Y(_1397_));
 sky130_fd_sc_hd__a21oi_1 _4616_ (.A1(_1396_),
    .A2(_1397_),
    .B1(_1395_),
    .Y(_1398_));
 sky130_fd_sc_hd__a31o_1 _4617_ (.A1(_1395_),
    .A2(_1396_),
    .A3(_1397_),
    .B1(net176),
    .X(_1399_));
 sky130_fd_sc_hd__o22a_1 _4618_ (.A1(net342),
    .A2(_2687_),
    .B1(_1398_),
    .B2(_1399_),
    .X(_1400_));
 sky130_fd_sc_hd__nor2_1 _4619_ (.A(_1363_),
    .B(_1367_),
    .Y(_1401_));
 sky130_fd_sc_hd__or2_2 _4620_ (.A(net342),
    .B(_2882_),
    .X(_1402_));
 sky130_fd_sc_hd__nand2_1 _4621_ (.A(net342),
    .B(_2882_),
    .Y(_1403_));
 sky130_fd_sc_hd__nand2_1 _4622_ (.A(_1402_),
    .B(_1403_),
    .Y(_1404_));
 sky130_fd_sc_hd__xor2_1 _4623_ (.A(_1401_),
    .B(_1404_),
    .X(_1405_));
 sky130_fd_sc_hd__mux2_1 _4624_ (.A0(net342),
    .A1(_1405_),
    .S(_1347_),
    .X(_1406_));
 sky130_fd_sc_hd__a22o_2 _4625_ (.A1(_0686_),
    .A2(_1400_),
    .B1(_1406_),
    .B2(net74),
    .X(_1407_));
 sky130_fd_sc_hd__and3_1 _4626_ (.A(net13),
    .B(net38),
    .C(net37),
    .X(_1408_));
 sky130_fd_sc_hd__a21oi_1 _4627_ (.A1(net38),
    .A2(net37),
    .B1(net13),
    .Y(_1409_));
 sky130_fd_sc_hd__or2_1 _4628_ (.A(_1408_),
    .B(_1409_),
    .X(_1410_));
 sky130_fd_sc_hd__nand2_2 _4629_ (.A(net279),
    .B(net341),
    .Y(_1411_));
 sky130_fd_sc_hd__or2_2 _4630_ (.A(net279),
    .B(net341),
    .X(_1412_));
 sky130_fd_sc_hd__nand2_4 _4631_ (.A(_1411_),
    .B(_1412_),
    .Y(_1413_));
 sky130_fd_sc_hd__and3_1 _4632_ (.A(_1373_),
    .B(_1376_),
    .C(_1413_),
    .X(_1414_));
 sky130_fd_sc_hd__a21oi_1 _4633_ (.A1(_1373_),
    .A2(_1376_),
    .B1(_1413_),
    .Y(_1415_));
 sky130_fd_sc_hd__o31a_1 _4634_ (.A1(net85),
    .A2(_1414_),
    .A3(_1415_),
    .B1(net53),
    .X(_1416_));
 sky130_fd_sc_hd__o21ai_1 _4635_ (.A1(_0683_),
    .A2(_1410_),
    .B1(_1416_),
    .Y(_1417_));
 sky130_fd_sc_hd__a21o_1 _4636_ (.A1(_0688_),
    .A2(_1407_),
    .B1(_1417_),
    .X(_1418_));
 sky130_fd_sc_hd__o2bb2a_1 _4637_ (.A1_N(net123),
    .A2_N(_1410_),
    .B1(_2616_),
    .B2(net13),
    .X(_1419_));
 sky130_fd_sc_hd__o211a_1 _4638_ (.A1(net341),
    .A2(_1383_),
    .B1(_1419_),
    .C1(_1334_),
    .X(_1420_));
 sky130_fd_sc_hd__a21o_1 _4639_ (.A1(net279),
    .A2(_1338_),
    .B1(net193),
    .X(_1421_));
 sky130_fd_sc_hd__o21a_2 _4640_ (.A1(_1327_),
    .A2(_1374_),
    .B1(_1373_),
    .X(_1422_));
 sky130_fd_sc_hd__xor2_4 _4641_ (.A(_1413_),
    .B(_1422_),
    .X(_1423_));
 sky130_fd_sc_hd__mux2_1 _4642_ (.A0(net13),
    .A1(_1423_),
    .S(net322),
    .X(_1424_));
 sky130_fd_sc_hd__a221o_1 _4643_ (.A1(net140),
    .A2(_1420_),
    .B1(_1424_),
    .B2(_1390_),
    .C1(_1421_),
    .X(_1425_));
 sky130_fd_sc_hd__o211a_1 _4644_ (.A1(net279),
    .A2(net151),
    .B1(_1418_),
    .C1(_1425_),
    .X(_1426_));
 sky130_fd_sc_hd__or2_1 _4645_ (.A(net13),
    .B(net39),
    .X(_1427_));
 sky130_fd_sc_hd__o22a_1 _4646_ (.A1(net279),
    .A2(net51),
    .B1(_1426_),
    .B2(net89),
    .X(_1428_));
 sky130_fd_sc_hd__o311a_1 _4647_ (.A1(_1319_),
    .A2(net42),
    .A3(_1428_),
    .B1(_1427_),
    .C1(net315),
    .X(_0175_));
 sky130_fd_sc_hd__and2_1 _4648_ (.A(net14),
    .B(_1408_),
    .X(_1429_));
 sky130_fd_sc_hd__nor2_1 _4649_ (.A(net14),
    .B(_1408_),
    .Y(_1430_));
 sky130_fd_sc_hd__or2_1 _4650_ (.A(_1429_),
    .B(_1430_),
    .X(_1431_));
 sky130_fd_sc_hd__nand2_1 _4651_ (.A(net91),
    .B(_1431_),
    .Y(_1432_));
 sky130_fd_sc_hd__and2_1 _4652_ (.A(net339),
    .B(_0288_),
    .X(_1433_));
 sky130_fd_sc_hd__or2_2 _4653_ (.A(net339),
    .B(_0288_),
    .X(_1434_));
 sky130_fd_sc_hd__and2b_1 _4654_ (.A_N(_1433_),
    .B(_1434_),
    .X(_1435_));
 sky130_fd_sc_hd__a221o_2 _4655_ (.A1(net342),
    .A2(_2886_),
    .B1(_1356_),
    .B2(_1358_),
    .C1(_1355_),
    .X(_1436_));
 sky130_fd_sc_hd__nand2_1 _4656_ (.A(_1396_),
    .B(_1436_),
    .Y(_1437_));
 sky130_fd_sc_hd__xor2_1 _4657_ (.A(_1435_),
    .B(_1437_),
    .X(_1438_));
 sky130_fd_sc_hd__nand2_1 _4658_ (.A(net339),
    .B(_2686_),
    .Y(_1439_));
 sky130_fd_sc_hd__o211a_1 _4659_ (.A1(net176),
    .A2(_1438_),
    .B1(_1439_),
    .C1(_0686_),
    .X(_1440_));
 sky130_fd_sc_hd__nor2_1 _4660_ (.A(_2552_),
    .B(_0284_),
    .Y(_1441_));
 sky130_fd_sc_hd__nor2_1 _4661_ (.A(net339),
    .B(_2932_),
    .Y(_1442_));
 sky130_fd_sc_hd__nand2_1 _4662_ (.A(_2552_),
    .B(_0284_),
    .Y(_1443_));
 sky130_fd_sc_hd__a221o_1 _4663_ (.A1(net342),
    .A2(_2882_),
    .B1(_1365_),
    .B2(_1366_),
    .C1(_1363_),
    .X(_1444_));
 sky130_fd_sc_hd__a211o_1 _4664_ (.A1(_1402_),
    .A2(_1444_),
    .B1(_1442_),
    .C1(_1441_),
    .X(_1445_));
 sky130_fd_sc_hd__o211ai_1 _4665_ (.A1(_1441_),
    .A2(_1442_),
    .B1(_1444_),
    .C1(_1402_),
    .Y(_1446_));
 sky130_fd_sc_hd__a32o_1 _4666_ (.A1(_1369_),
    .A2(_1445_),
    .A3(_1446_),
    .B1(_1362_),
    .B2(_2552_),
    .X(_1447_));
 sky130_fd_sc_hd__nor2_2 _4667_ (.A(_1440_),
    .B(_1447_),
    .Y(_1448_));
 sky130_fd_sc_hd__o211a_1 _4668_ (.A1(_0689_),
    .A2(_1448_),
    .B1(_1432_),
    .C1(net85),
    .X(_1449_));
 sky130_fd_sc_hd__or2_1 _4669_ (.A(net277),
    .B(net338),
    .X(_1450_));
 sky130_fd_sc_hd__nand2_2 _4670_ (.A(net277),
    .B(net338),
    .Y(_1451_));
 sky130_fd_sc_hd__nand2_2 _4671_ (.A(_1450_),
    .B(_1451_),
    .Y(_1452_));
 sky130_fd_sc_hd__a21o_1 _4672_ (.A1(net279),
    .A2(net341),
    .B1(_1415_),
    .X(_1453_));
 sky130_fd_sc_hd__xnor2_1 _4673_ (.A(_1452_),
    .B(_1453_),
    .Y(_1454_));
 sky130_fd_sc_hd__a211o_1 _4674_ (.A1(net86),
    .A2(_1454_),
    .B1(_1449_),
    .C1(_0694_),
    .X(_1455_));
 sky130_fd_sc_hd__o21ai_1 _4675_ (.A1(net127),
    .A2(_1431_),
    .B1(_1334_),
    .Y(_1456_));
 sky130_fd_sc_hd__a31o_1 _4676_ (.A1(net294),
    .A2(net338),
    .A3(net127),
    .B1(_1456_),
    .X(_1457_));
 sky130_fd_sc_hd__a21oi_1 _4677_ (.A1(net14),
    .A2(_2615_),
    .B1(_1457_),
    .Y(_1458_));
 sky130_fd_sc_hd__o21a_1 _4678_ (.A1(_1413_),
    .A2(_1422_),
    .B1(_1411_),
    .X(_1459_));
 sky130_fd_sc_hd__xor2_2 _4679_ (.A(_1452_),
    .B(_1459_),
    .X(_1460_));
 sky130_fd_sc_hd__nand2_1 _4680_ (.A(net322),
    .B(_1460_),
    .Y(_1461_));
 sky130_fd_sc_hd__o211a_1 _4681_ (.A1(_2541_),
    .A2(net322),
    .B1(_1342_),
    .C1(_1461_),
    .X(_1462_));
 sky130_fd_sc_hd__nor2_1 _4682_ (.A(_1458_),
    .B(_1462_),
    .Y(_1463_));
 sky130_fd_sc_hd__o22a_1 _4683_ (.A1(net277),
    .A2(_1337_),
    .B1(_1463_),
    .B2(net76),
    .X(_1464_));
 sky130_fd_sc_hd__o221a_1 _4684_ (.A1(net277),
    .A2(net151),
    .B1(_1464_),
    .B2(net193),
    .C1(_1455_),
    .X(_1465_));
 sky130_fd_sc_hd__o22a_1 _4685_ (.A1(net277),
    .A2(net51),
    .B1(_1465_),
    .B2(net89),
    .X(_1466_));
 sky130_fd_sc_hd__or2_1 _4686_ (.A(net14),
    .B(net39),
    .X(_1467_));
 sky130_fd_sc_hd__o311a_1 _4687_ (.A1(_1319_),
    .A2(net42),
    .A3(_1466_),
    .B1(_1467_),
    .C1(net314),
    .X(_0176_));
 sky130_fd_sc_hd__o22a_1 _4688_ (.A1(net15),
    .A2(_2616_),
    .B1(_1383_),
    .B2(net337),
    .X(_1468_));
 sky130_fd_sc_hd__xnor2_1 _4689_ (.A(net15),
    .B(_1429_),
    .Y(_1469_));
 sky130_fd_sc_hd__inv_2 _4690_ (.A(_1469_),
    .Y(_1470_));
 sky130_fd_sc_hd__o211a_1 _4691_ (.A1(net127),
    .A2(_1470_),
    .B1(_1468_),
    .C1(_1334_),
    .X(_1471_));
 sky130_fd_sc_hd__nand2_2 _4692_ (.A(net276),
    .B(net337),
    .Y(_1472_));
 sky130_fd_sc_hd__or2_1 _4693_ (.A(net276),
    .B(net337),
    .X(_1473_));
 sky130_fd_sc_hd__nand2_1 _4694_ (.A(_1472_),
    .B(_1473_),
    .Y(_1474_));
 sky130_fd_sc_hd__o21bai_1 _4695_ (.A1(net277),
    .A2(net338),
    .B1_N(_1459_),
    .Y(_1475_));
 sky130_fd_sc_hd__a21o_2 _4696_ (.A1(_1451_),
    .A2(_1475_),
    .B1(_1474_),
    .X(_1476_));
 sky130_fd_sc_hd__nand3_1 _4697_ (.A(_1451_),
    .B(_1474_),
    .C(_1475_),
    .Y(_1477_));
 sky130_fd_sc_hd__nand2_1 _4698_ (.A(_1476_),
    .B(_1477_),
    .Y(_1478_));
 sky130_fd_sc_hd__nand2_1 _4699_ (.A(net322),
    .B(_1478_),
    .Y(_1479_));
 sky130_fd_sc_hd__or2_1 _4700_ (.A(net15),
    .B(net322),
    .X(_1480_));
 sky130_fd_sc_hd__a31o_1 _4701_ (.A1(_1342_),
    .A2(_1479_),
    .A3(_1480_),
    .B1(_1471_),
    .X(_1481_));
 sky130_fd_sc_hd__a221o_1 _4702_ (.A1(net276),
    .A2(_1338_),
    .B1(_1481_),
    .B2(net140),
    .C1(net193),
    .X(_1482_));
 sky130_fd_sc_hd__nor2_1 _4703_ (.A(_2553_),
    .B(_0341_),
    .Y(_1483_));
 sky130_fd_sc_hd__xnor2_2 _4704_ (.A(net335),
    .B(_0340_),
    .Y(_1484_));
 sky130_fd_sc_hd__a31oi_4 _4705_ (.A1(_1396_),
    .A2(_1434_),
    .A3(_1436_),
    .B1(_1433_),
    .Y(_1485_));
 sky130_fd_sc_hd__or2_1 _4706_ (.A(_1484_),
    .B(_1485_),
    .X(_1486_));
 sky130_fd_sc_hd__nand2_1 _4707_ (.A(_1484_),
    .B(_1485_),
    .Y(_1487_));
 sky130_fd_sc_hd__a21o_1 _4708_ (.A1(_1486_),
    .A2(_1487_),
    .B1(net176),
    .X(_1488_));
 sky130_fd_sc_hd__o211a_1 _4709_ (.A1(net335),
    .A2(_2687_),
    .B1(_0686_),
    .C1(_1488_),
    .X(_1489_));
 sky130_fd_sc_hd__and2_1 _4710_ (.A(net335),
    .B(_0337_),
    .X(_1490_));
 sky130_fd_sc_hd__or2_1 _4711_ (.A(net335),
    .B(_0337_),
    .X(_1491_));
 sky130_fd_sc_hd__and2b_1 _4712_ (.A_N(_1490_),
    .B(_1491_),
    .X(_1492_));
 sky130_fd_sc_hd__a31o_1 _4713_ (.A1(_1402_),
    .A2(_1443_),
    .A3(_1444_),
    .B1(_1441_),
    .X(_1493_));
 sky130_fd_sc_hd__nand2_1 _4714_ (.A(_1492_),
    .B(_1493_),
    .Y(_1494_));
 sky130_fd_sc_hd__o211a_1 _4715_ (.A1(_1492_),
    .A2(_1493_),
    .B1(_1494_),
    .C1(_1369_),
    .X(_1495_));
 sky130_fd_sc_hd__a211o_4 _4716_ (.A1(net335),
    .A2(_1362_),
    .B1(_1489_),
    .C1(_1495_),
    .X(_1496_));
 sky130_fd_sc_hd__nand2_1 _4717_ (.A(_1450_),
    .B(_1453_),
    .Y(_1497_));
 sky130_fd_sc_hd__a21o_2 _4718_ (.A1(_1451_),
    .A2(_1497_),
    .B1(_1474_),
    .X(_1498_));
 sky130_fd_sc_hd__inv_2 _4719_ (.A(_1498_),
    .Y(_1499_));
 sky130_fd_sc_hd__nand3_1 _4720_ (.A(_1451_),
    .B(_1474_),
    .C(_1497_),
    .Y(_1500_));
 sky130_fd_sc_hd__a32o_1 _4721_ (.A1(net86),
    .A2(_1498_),
    .A3(_1500_),
    .B1(_1496_),
    .B2(_0688_),
    .X(_1501_));
 sky130_fd_sc_hd__a211o_1 _4722_ (.A1(net91),
    .A2(_1470_),
    .B1(_1501_),
    .C1(_0694_),
    .X(_1502_));
 sky130_fd_sc_hd__o211a_1 _4723_ (.A1(net276),
    .A2(net151),
    .B1(_1482_),
    .C1(_1502_),
    .X(_1503_));
 sky130_fd_sc_hd__o22a_1 _4724_ (.A1(net276),
    .A2(net51),
    .B1(_1503_),
    .B2(net89),
    .X(_1504_));
 sky130_fd_sc_hd__or2_1 _4725_ (.A(net15),
    .B(net39),
    .X(_1505_));
 sky130_fd_sc_hd__o311a_1 _4726_ (.A1(_1319_),
    .A2(net42),
    .A3(_1504_),
    .B1(_1505_),
    .C1(net314),
    .X(_0177_));
 sky130_fd_sc_hd__and3_1 _4727_ (.A(net16),
    .B(net15),
    .C(_1429_),
    .X(_1506_));
 sky130_fd_sc_hd__a21oi_1 _4728_ (.A1(net15),
    .A2(_1429_),
    .B1(net16),
    .Y(_1507_));
 sky130_fd_sc_hd__or2_1 _4729_ (.A(_1506_),
    .B(_1507_),
    .X(_1508_));
 sky130_fd_sc_hd__a21oi_1 _4730_ (.A1(net91),
    .A2(_1508_),
    .B1(net86),
    .Y(_1509_));
 sky130_fd_sc_hd__and2_1 _4731_ (.A(net332),
    .B(_0396_),
    .X(_1510_));
 sky130_fd_sc_hd__nor2_2 _4732_ (.A(net332),
    .B(_0396_),
    .Y(_1511_));
 sky130_fd_sc_hd__or2_1 _4733_ (.A(_1510_),
    .B(_1511_),
    .X(_1512_));
 sky130_fd_sc_hd__o21ba_2 _4734_ (.A1(_1484_),
    .A2(_1485_),
    .B1_N(_1483_),
    .X(_1513_));
 sky130_fd_sc_hd__or2_1 _4735_ (.A(_1512_),
    .B(_1513_),
    .X(_1514_));
 sky130_fd_sc_hd__a21oi_1 _4736_ (.A1(_1512_),
    .A2(_1513_),
    .B1(net176),
    .Y(_1515_));
 sky130_fd_sc_hd__a22o_1 _4737_ (.A1(net332),
    .A2(net176),
    .B1(_1514_),
    .B2(_1515_),
    .X(_1516_));
 sky130_fd_sc_hd__and2_1 _4738_ (.A(net332),
    .B(_0394_),
    .X(_1517_));
 sky130_fd_sc_hd__or2_1 _4739_ (.A(net332),
    .B(_0394_),
    .X(_1518_));
 sky130_fd_sc_hd__nand2b_1 _4740_ (.A_N(_1517_),
    .B(_1518_),
    .Y(_1519_));
 sky130_fd_sc_hd__o21a_1 _4741_ (.A1(_1490_),
    .A2(_1493_),
    .B1(_1491_),
    .X(_1520_));
 sky130_fd_sc_hd__xnor2_1 _4742_ (.A(_1519_),
    .B(_1520_),
    .Y(_1521_));
 sky130_fd_sc_hd__mux2_1 _4743_ (.A0(net332),
    .A1(_1521_),
    .S(_1347_),
    .X(_1522_));
 sky130_fd_sc_hd__o22a_2 _4744_ (.A1(_0687_),
    .A2(_1516_),
    .B1(_1522_),
    .B2(net72),
    .X(_1523_));
 sky130_fd_sc_hd__o21ai_1 _4745_ (.A1(_0689_),
    .A2(_1523_),
    .B1(_1509_),
    .Y(_1524_));
 sky130_fd_sc_hd__nand2_2 _4746_ (.A(net273),
    .B(net334),
    .Y(_1525_));
 sky130_fd_sc_hd__or2_4 _4747_ (.A(net273),
    .B(net334),
    .X(_1526_));
 sky130_fd_sc_hd__nand2_4 _4748_ (.A(_1525_),
    .B(_1526_),
    .Y(_1527_));
 sky130_fd_sc_hd__a21oi_1 _4749_ (.A1(_1472_),
    .A2(_1498_),
    .B1(_1527_),
    .Y(_1528_));
 sky130_fd_sc_hd__a31o_1 _4750_ (.A1(_1472_),
    .A2(_1498_),
    .A3(_1527_),
    .B1(net85),
    .X(_1529_));
 sky130_fd_sc_hd__o211ai_1 _4751_ (.A1(_1528_),
    .A2(_1529_),
    .B1(net53),
    .C1(_1524_),
    .Y(_1530_));
 sky130_fd_sc_hd__o221a_1 _4752_ (.A1(_2540_),
    .A2(_2616_),
    .B1(_1383_),
    .B2(_2554_),
    .C1(_1334_),
    .X(_1531_));
 sky130_fd_sc_hd__nand2_1 _4753_ (.A(net334),
    .B(net129),
    .Y(_1532_));
 sky130_fd_sc_hd__o21a_1 _4754_ (.A1(net127),
    .A2(_1508_),
    .B1(_1531_),
    .X(_1533_));
 sky130_fd_sc_hd__nand2_1 _4755_ (.A(_1472_),
    .B(_1476_),
    .Y(_1534_));
 sky130_fd_sc_hd__xnor2_2 _4756_ (.A(_1527_),
    .B(_1534_),
    .Y(_1535_));
 sky130_fd_sc_hd__nand2_1 _4757_ (.A(net322),
    .B(_1535_),
    .Y(_1536_));
 sky130_fd_sc_hd__o211a_1 _4758_ (.A1(_2540_),
    .A2(net323),
    .B1(_1342_),
    .C1(_1536_),
    .X(_1537_));
 sky130_fd_sc_hd__nor2_1 _4759_ (.A(_1533_),
    .B(_1537_),
    .Y(_1538_));
 sky130_fd_sc_hd__o22a_1 _4760_ (.A1(net273),
    .A2(_1337_),
    .B1(_1538_),
    .B2(net76),
    .X(_1539_));
 sky130_fd_sc_hd__o221a_1 _4761_ (.A1(net273),
    .A2(net151),
    .B1(_1539_),
    .B2(net193),
    .C1(_1530_),
    .X(_1540_));
 sky130_fd_sc_hd__o22a_1 _4762_ (.A1(net273),
    .A2(net51),
    .B1(_1540_),
    .B2(net89),
    .X(_1541_));
 sky130_fd_sc_hd__or2_1 _4763_ (.A(net16),
    .B(net39),
    .X(_1542_));
 sky130_fd_sc_hd__o311a_1 _4764_ (.A1(_1319_),
    .A2(net42),
    .A3(_1541_),
    .B1(_1542_),
    .C1(net314),
    .X(_0178_));
 sky130_fd_sc_hd__and2_2 _4765_ (.A(net17),
    .B(_1506_),
    .X(_1543_));
 sky130_fd_sc_hd__nor2_1 _4766_ (.A(net17),
    .B(_1506_),
    .Y(_1544_));
 sky130_fd_sc_hd__or2_1 _4767_ (.A(_1543_),
    .B(_1544_),
    .X(_1545_));
 sky130_fd_sc_hd__nand2_1 _4768_ (.A(net123),
    .B(_1545_),
    .Y(_1546_));
 sky130_fd_sc_hd__o221a_1 _4769_ (.A1(net17),
    .A2(_2616_),
    .B1(_1383_),
    .B2(net328),
    .C1(_1334_),
    .X(_1547_));
 sky130_fd_sc_hd__and2_2 _4770_ (.A(net271),
    .B(net328),
    .X(_1548_));
 sky130_fd_sc_hd__nor2_2 _4771_ (.A(net271),
    .B(net328),
    .Y(_1549_));
 sky130_fd_sc_hd__nor2_4 _4772_ (.A(_1548_),
    .B(_1549_),
    .Y(_1550_));
 sky130_fd_sc_hd__nand2_1 _4773_ (.A(_1472_),
    .B(_1525_),
    .Y(_1551_));
 sky130_fd_sc_hd__nand2_2 _4774_ (.A(_1526_),
    .B(_1551_),
    .Y(_1552_));
 sky130_fd_sc_hd__o21ai_4 _4775_ (.A1(_1476_),
    .A2(_1527_),
    .B1(_1552_),
    .Y(_1553_));
 sky130_fd_sc_hd__xnor2_4 _4776_ (.A(_1550_),
    .B(_1553_),
    .Y(_1554_));
 sky130_fd_sc_hd__nand2_1 _4777_ (.A(net322),
    .B(_1554_),
    .Y(_1555_));
 sky130_fd_sc_hd__o211a_1 _4778_ (.A1(net17),
    .A2(net322),
    .B1(_1342_),
    .C1(_1555_),
    .X(_1556_));
 sky130_fd_sc_hd__a21o_1 _4779_ (.A1(_1546_),
    .A2(_1547_),
    .B1(_1556_),
    .X(_1557_));
 sky130_fd_sc_hd__a221o_1 _4780_ (.A1(net271),
    .A2(_1338_),
    .B1(_1557_),
    .B2(net140),
    .C1(net193),
    .X(_1558_));
 sky130_fd_sc_hd__and2_1 _4781_ (.A(net331),
    .B(_0439_),
    .X(_1559_));
 sky130_fd_sc_hd__xnor2_1 _4782_ (.A(net331),
    .B(_0439_),
    .Y(_1560_));
 sky130_fd_sc_hd__inv_2 _4783_ (.A(_1560_),
    .Y(_1561_));
 sky130_fd_sc_hd__o21bai_4 _4784_ (.A1(_1511_),
    .A2(_1513_),
    .B1_N(_1510_),
    .Y(_1562_));
 sky130_fd_sc_hd__xnor2_1 _4785_ (.A(_1561_),
    .B(_1562_),
    .Y(_1563_));
 sky130_fd_sc_hd__mux2_2 _4786_ (.A0(_2556_),
    .A1(_1563_),
    .S(_2687_),
    .X(_1564_));
 sky130_fd_sc_hd__xnor2_1 _4787_ (.A(_2556_),
    .B(_0436_),
    .Y(_1565_));
 sky130_fd_sc_hd__o21a_1 _4788_ (.A1(_1517_),
    .A2(_1520_),
    .B1(_1518_),
    .X(_1566_));
 sky130_fd_sc_hd__o211a_2 _4789_ (.A1(_1517_),
    .A2(_1520_),
    .B1(_1565_),
    .C1(_1518_),
    .X(_1567_));
 sky130_fd_sc_hd__o21ai_1 _4790_ (.A1(_1565_),
    .A2(_1566_),
    .B1(_1369_),
    .Y(_1568_));
 sky130_fd_sc_hd__o2bb2a_1 _4791_ (.A1_N(net331),
    .A2_N(_1362_),
    .B1(_1567_),
    .B2(_1568_),
    .X(_1569_));
 sky130_fd_sc_hd__o21ai_4 _4792_ (.A1(_0687_),
    .A2(_1564_),
    .B1(_1569_),
    .Y(_1570_));
 sky130_fd_sc_hd__o211a_1 _4793_ (.A1(_1499_),
    .A2(_1551_),
    .B1(_1550_),
    .C1(_1526_),
    .X(_1571_));
 sky130_fd_sc_hd__o221a_1 _4794_ (.A1(_1498_),
    .A2(_1527_),
    .B1(_1548_),
    .B2(_1549_),
    .C1(_1552_),
    .X(_1572_));
 sky130_fd_sc_hd__or3_1 _4795_ (.A(net85),
    .B(_1571_),
    .C(_1572_),
    .X(_1573_));
 sky130_fd_sc_hd__o211a_1 _4796_ (.A1(_0683_),
    .A2(_1545_),
    .B1(_1573_),
    .C1(net53),
    .X(_1574_));
 sky130_fd_sc_hd__a21bo_1 _4797_ (.A1(_0688_),
    .A2(_1570_),
    .B1_N(_1574_),
    .X(_1575_));
 sky130_fd_sc_hd__o211a_1 _4798_ (.A1(net271),
    .A2(net151),
    .B1(_1558_),
    .C1(_1575_),
    .X(_1576_));
 sky130_fd_sc_hd__or2_1 _4799_ (.A(net17),
    .B(net39),
    .X(_1577_));
 sky130_fd_sc_hd__o22a_1 _4800_ (.A1(net271),
    .A2(net51),
    .B1(_1576_),
    .B2(net89),
    .X(_1578_));
 sky130_fd_sc_hd__o311a_1 _4801_ (.A1(_1319_),
    .A2(net42),
    .A3(_1578_),
    .B1(_1577_),
    .C1(net314),
    .X(_0179_));
 sky130_fd_sc_hd__xnor2_1 _4802_ (.A(net18),
    .B(_1543_),
    .Y(_1579_));
 sky130_fd_sc_hd__a21oi_2 _4803_ (.A1(_1561_),
    .A2(_1562_),
    .B1(_1559_),
    .Y(_1580_));
 sky130_fd_sc_hd__nand2_1 _4804_ (.A(net326),
    .B(_0477_),
    .Y(_1581_));
 sky130_fd_sc_hd__nor2_1 _4805_ (.A(net326),
    .B(_0477_),
    .Y(_1582_));
 sky130_fd_sc_hd__or2_1 _4806_ (.A(net326),
    .B(_0477_),
    .X(_1583_));
 sky130_fd_sc_hd__nand2_1 _4807_ (.A(_1581_),
    .B(_1583_),
    .Y(_1584_));
 sky130_fd_sc_hd__or2_1 _4808_ (.A(_1580_),
    .B(_1584_),
    .X(_1585_));
 sky130_fd_sc_hd__a21oi_1 _4809_ (.A1(_1580_),
    .A2(_1584_),
    .B1(net176),
    .Y(_1586_));
 sky130_fd_sc_hd__a22o_1 _4810_ (.A1(net326),
    .A2(net176),
    .B1(_1585_),
    .B2(_1586_),
    .X(_1587_));
 sky130_fd_sc_hd__a21oi_4 _4811_ (.A1(net331),
    .A2(_0436_),
    .B1(_1567_),
    .Y(_1588_));
 sky130_fd_sc_hd__nand2_2 _4812_ (.A(net326),
    .B(_0474_),
    .Y(_1589_));
 sky130_fd_sc_hd__or2_1 _4813_ (.A(net326),
    .B(_0474_),
    .X(_1590_));
 sky130_fd_sc_hd__nand2_1 _4814_ (.A(_1589_),
    .B(_1590_),
    .Y(_1591_));
 sky130_fd_sc_hd__nand2_1 _4815_ (.A(_1588_),
    .B(_1591_),
    .Y(_1592_));
 sky130_fd_sc_hd__o21a_1 _4816_ (.A1(_1588_),
    .A2(_1591_),
    .B1(_1347_),
    .X(_1593_));
 sky130_fd_sc_hd__a2bb2o_1 _4817_ (.A1_N(net312),
    .A2_N(_1347_),
    .B1(_1592_),
    .B2(_1593_),
    .X(_1594_));
 sky130_fd_sc_hd__o22ai_4 _4818_ (.A1(_0687_),
    .A2(_1587_),
    .B1(_1594_),
    .B2(net72),
    .Y(_1595_));
 sky130_fd_sc_hd__a22o_1 _4819_ (.A1(net91),
    .A2(_1579_),
    .B1(_1595_),
    .B2(_0720_),
    .X(_1596_));
 sky130_fd_sc_hd__xor2_4 _4820_ (.A(net269),
    .B(net328),
    .X(_1597_));
 sky130_fd_sc_hd__o21ai_1 _4821_ (.A1(_1548_),
    .A2(_1571_),
    .B1(_1597_),
    .Y(_1598_));
 sky130_fd_sc_hd__or3_1 _4822_ (.A(_1548_),
    .B(_1571_),
    .C(_1597_),
    .X(_1599_));
 sky130_fd_sc_hd__a31o_1 _4823_ (.A1(net86),
    .A2(_1598_),
    .A3(_1599_),
    .B1(_0694_),
    .X(_1600_));
 sky130_fd_sc_hd__o21ba_1 _4824_ (.A1(net86),
    .A2(_1596_),
    .B1_N(_1600_),
    .X(_1601_));
 sky130_fd_sc_hd__nor2_1 _4825_ (.A(net127),
    .B(_1579_),
    .Y(_1602_));
 sky130_fd_sc_hd__a221o_1 _4826_ (.A1(net18),
    .A2(_2615_),
    .B1(_1382_),
    .B2(net324),
    .C1(net149),
    .X(_1603_));
 sky130_fd_sc_hd__o22a_1 _4827_ (.A1(net269),
    .A2(net84),
    .B1(_1602_),
    .B2(_1603_),
    .X(_1604_));
 sky130_fd_sc_hd__o22a_1 _4828_ (.A1(net269),
    .A2(net50),
    .B1(_1604_),
    .B2(net75),
    .X(_1605_));
 sky130_fd_sc_hd__nor2_1 _4829_ (.A(net202),
    .B(_1605_),
    .Y(_1606_));
 sky130_fd_sc_hd__a21oi_2 _4830_ (.A1(_1550_),
    .A2(_1553_),
    .B1(_1548_),
    .Y(_1607_));
 sky130_fd_sc_hd__xnor2_2 _4831_ (.A(_1597_),
    .B(_1607_),
    .Y(_1608_));
 sky130_fd_sc_hd__a21bo_1 _4832_ (.A1(net322),
    .A2(_1608_),
    .B1_N(_1390_),
    .X(_1609_));
 sky130_fd_sc_hd__a211oi_1 _4833_ (.A1(net18),
    .A2(net309),
    .B1(net193),
    .C1(_1609_),
    .Y(_1610_));
 sky130_fd_sc_hd__o31a_1 _4834_ (.A1(_1601_),
    .A2(_1606_),
    .A3(_1610_),
    .B1(net88),
    .X(_1611_));
 sky130_fd_sc_hd__nor2_1 _4835_ (.A(net269),
    .B(net51),
    .Y(_1612_));
 sky130_fd_sc_hd__o21ai_1 _4836_ (.A1(_1611_),
    .A2(_1612_),
    .B1(net39),
    .Y(_1613_));
 sky130_fd_sc_hd__o211a_1 _4837_ (.A1(net18),
    .A2(net39),
    .B1(_1613_),
    .C1(net314),
    .X(_0180_));
 sky130_fd_sc_hd__and3_1 _4838_ (.A(net19),
    .B(net18),
    .C(_1543_),
    .X(_1614_));
 sky130_fd_sc_hd__a21oi_1 _4839_ (.A1(net18),
    .A2(_1543_),
    .B1(net19),
    .Y(_1615_));
 sky130_fd_sc_hd__or2_1 _4840_ (.A(_1614_),
    .B(_1615_),
    .X(_1616_));
 sky130_fd_sc_hd__a211o_4 _4841_ (.A1(_1580_),
    .A2(_1581_),
    .B1(_1582_),
    .C1(net176),
    .X(_1617_));
 sky130_fd_sc_hd__nor2_1 _4842_ (.A(_2557_),
    .B(_1617_),
    .Y(_1618_));
 sky130_fd_sc_hd__nand2_1 _4843_ (.A(_2557_),
    .B(_1617_),
    .Y(_1619_));
 sky130_fd_sc_hd__nand2b_1 _4844_ (.A_N(_1618_),
    .B(_1619_),
    .Y(_1620_));
 sky130_fd_sc_hd__o21ai_4 _4845_ (.A1(net326),
    .A2(_0474_),
    .B1(_1347_),
    .Y(_1621_));
 sky130_fd_sc_hd__a21oi_4 _4846_ (.A1(_1588_),
    .A2(_1589_),
    .B1(_1621_),
    .Y(_1622_));
 sky130_fd_sc_hd__nand2_1 _4847_ (.A(net296),
    .B(_1622_),
    .Y(_1623_));
 sky130_fd_sc_hd__or2_1 _4848_ (.A(net296),
    .B(_1622_),
    .X(_1624_));
 sky130_fd_sc_hd__nand2_1 _4849_ (.A(_1623_),
    .B(_1624_),
    .Y(_1625_));
 sky130_fd_sc_hd__a22o_1 _4850_ (.A1(_0686_),
    .A2(_1620_),
    .B1(_1625_),
    .B2(net74),
    .X(_1626_));
 sky130_fd_sc_hd__a22o_1 _4851_ (.A1(net91),
    .A2(_1616_),
    .B1(_1626_),
    .B2(_0720_),
    .X(_1627_));
 sky130_fd_sc_hd__nand2_1 _4852_ (.A(net268),
    .B(net328),
    .Y(_1628_));
 sky130_fd_sc_hd__or2_1 _4853_ (.A(net268),
    .B(net328),
    .X(_1629_));
 sky130_fd_sc_hd__nand2_1 _4854_ (.A(_1628_),
    .B(_1629_),
    .Y(_1630_));
 sky130_fd_sc_hd__nand2_1 _4855_ (.A(_1550_),
    .B(_1597_),
    .Y(_1631_));
 sky130_fd_sc_hd__o21ai_1 _4856_ (.A1(net269),
    .A2(net271),
    .B1(net328),
    .Y(_1632_));
 sky130_fd_sc_hd__o21a_1 _4857_ (.A1(_1552_),
    .A2(_1631_),
    .B1(_1632_),
    .X(_1633_));
 sky130_fd_sc_hd__or2_1 _4858_ (.A(_1527_),
    .B(_1631_),
    .X(_1634_));
 sky130_fd_sc_hd__o21a_1 _4859_ (.A1(_1498_),
    .A2(_1634_),
    .B1(_1633_),
    .X(_1635_));
 sky130_fd_sc_hd__or2_2 _4860_ (.A(_1630_),
    .B(_1635_),
    .X(_1636_));
 sky130_fd_sc_hd__nand2_1 _4861_ (.A(_1630_),
    .B(_1635_),
    .Y(_1637_));
 sky130_fd_sc_hd__a31o_1 _4862_ (.A1(net86),
    .A2(_1636_),
    .A3(_1637_),
    .B1(_0694_),
    .X(_1638_));
 sky130_fd_sc_hd__o21ba_1 _4863_ (.A1(net86),
    .A2(_1627_),
    .B1_N(_1638_),
    .X(_1639_));
 sky130_fd_sc_hd__o221a_1 _4864_ (.A1(net19),
    .A2(_2616_),
    .B1(_1383_),
    .B2(net296),
    .C1(_1334_),
    .X(_1640_));
 sky130_fd_sc_hd__a21boi_1 _4865_ (.A1(net123),
    .A2(_1616_),
    .B1_N(_1640_),
    .Y(_1641_));
 sky130_fd_sc_hd__o21a_1 _4866_ (.A1(_1476_),
    .A2(_1634_),
    .B1(_1633_),
    .X(_1642_));
 sky130_fd_sc_hd__or2_1 _4867_ (.A(_1630_),
    .B(_1642_),
    .X(_1643_));
 sky130_fd_sc_hd__nand2_1 _4868_ (.A(_1630_),
    .B(_1642_),
    .Y(_1644_));
 sky130_fd_sc_hd__nand2_1 _4869_ (.A(_1643_),
    .B(_1644_),
    .Y(_1645_));
 sky130_fd_sc_hd__nand2_1 _4870_ (.A(net323),
    .B(_1645_),
    .Y(_1646_));
 sky130_fd_sc_hd__o211a_1 _4871_ (.A1(net19),
    .A2(net323),
    .B1(_1342_),
    .C1(_1646_),
    .X(_1647_));
 sky130_fd_sc_hd__o21ai_1 _4872_ (.A1(_1641_),
    .A2(_1647_),
    .B1(net50),
    .Y(_1648_));
 sky130_fd_sc_hd__or2_1 _4873_ (.A(_2532_),
    .B(_1339_),
    .X(_1649_));
 sky130_fd_sc_hd__a31o_1 _4874_ (.A1(net225),
    .A2(_1648_),
    .A3(_1649_),
    .B1(_1639_),
    .X(_1650_));
 sky130_fd_sc_hd__a2bb2o_1 _4875_ (.A1_N(net268),
    .A2_N(net51),
    .B1(_1650_),
    .B2(net88),
    .X(_1651_));
 sky130_fd_sc_hd__nand2_1 _4876_ (.A(net40),
    .B(_1651_),
    .Y(_1652_));
 sky130_fd_sc_hd__o211a_1 _4877_ (.A1(net19),
    .A2(net40),
    .B1(_1652_),
    .C1(net314),
    .X(_0181_));
 sky130_fd_sc_hd__and2_1 _4878_ (.A(net20),
    .B(_1614_),
    .X(_1653_));
 sky130_fd_sc_hd__nor2_1 _4879_ (.A(net20),
    .B(_1614_),
    .Y(_1654_));
 sky130_fd_sc_hd__or2_1 _4880_ (.A(_1653_),
    .B(_1654_),
    .X(_1655_));
 sky130_fd_sc_hd__xor2_1 _4881_ (.A(net295),
    .B(_1623_),
    .X(_1656_));
 sky130_fd_sc_hd__xnor2_1 _4882_ (.A(net295),
    .B(_1618_),
    .Y(_1657_));
 sky130_fd_sc_hd__a22o_1 _4883_ (.A1(net74),
    .A2(_1656_),
    .B1(_1657_),
    .B2(_0686_),
    .X(_1658_));
 sky130_fd_sc_hd__a22o_1 _4884_ (.A1(net91),
    .A2(_1655_),
    .B1(_1658_),
    .B2(_0720_),
    .X(_1659_));
 sky130_fd_sc_hd__nor2_1 _4885_ (.A(net86),
    .B(_1659_),
    .Y(_1660_));
 sky130_fd_sc_hd__xnor2_4 _4886_ (.A(net267),
    .B(net328),
    .Y(_1661_));
 sky130_fd_sc_hd__a21oi_1 _4887_ (.A1(_1628_),
    .A2(_1636_),
    .B1(_1661_),
    .Y(_1662_));
 sky130_fd_sc_hd__a31o_1 _4888_ (.A1(_1628_),
    .A2(_1636_),
    .A3(_1661_),
    .B1(net85),
    .X(_1663_));
 sky130_fd_sc_hd__nor2_1 _4889_ (.A(_1662_),
    .B(_1663_),
    .Y(_1664_));
 sky130_fd_sc_hd__nor2_1 _4890_ (.A(net128),
    .B(_1655_),
    .Y(_1665_));
 sky130_fd_sc_hd__a221o_1 _4891_ (.A1(net20),
    .A2(_2615_),
    .B1(_1382_),
    .B2(net295),
    .C1(net149),
    .X(_1666_));
 sky130_fd_sc_hd__o22a_1 _4892_ (.A1(net267),
    .A2(net84),
    .B1(_1665_),
    .B2(_1666_),
    .X(_1667_));
 sky130_fd_sc_hd__o22a_1 _4893_ (.A1(net267),
    .A2(net50),
    .B1(_1667_),
    .B2(net75),
    .X(_1668_));
 sky130_fd_sc_hd__nand2_1 _4894_ (.A(_1628_),
    .B(_1643_),
    .Y(_1669_));
 sky130_fd_sc_hd__xnor2_2 _4895_ (.A(_1661_),
    .B(_1669_),
    .Y(_1670_));
 sky130_fd_sc_hd__a21bo_1 _4896_ (.A1(net20),
    .A2(net310),
    .B1_N(_1390_),
    .X(_1671_));
 sky130_fd_sc_hd__a211o_1 _4897_ (.A1(net324),
    .A2(_1670_),
    .B1(_1671_),
    .C1(net193),
    .X(_1672_));
 sky130_fd_sc_hd__o21a_1 _4898_ (.A1(net202),
    .A2(_1668_),
    .B1(_1672_),
    .X(_1673_));
 sky130_fd_sc_hd__o31a_1 _4899_ (.A1(_0694_),
    .A2(_1660_),
    .A3(_1664_),
    .B1(_1673_),
    .X(_1674_));
 sky130_fd_sc_hd__o22a_1 _4900_ (.A1(net267),
    .A2(net51),
    .B1(_1674_),
    .B2(net89),
    .X(_1675_));
 sky130_fd_sc_hd__or2_1 _4901_ (.A(net20),
    .B(net40),
    .X(_1676_));
 sky130_fd_sc_hd__o311a_1 _4902_ (.A1(_1319_),
    .A2(net42),
    .A3(_1675_),
    .B1(_1676_),
    .C1(net318),
    .X(_0182_));
 sky130_fd_sc_hd__nand2_1 _4903_ (.A(net21),
    .B(_1653_),
    .Y(_1677_));
 sky130_fd_sc_hd__or2_1 _4904_ (.A(net21),
    .B(_1653_),
    .X(_1678_));
 sky130_fd_sc_hd__nand2_1 _4905_ (.A(_1677_),
    .B(_1678_),
    .Y(_1679_));
 sky130_fd_sc_hd__nand2_1 _4906_ (.A(net73),
    .B(_1617_),
    .Y(_1680_));
 sky130_fd_sc_hd__and3_4 _4907_ (.A(\as2650.addr_buff[0] ),
    .B(net295),
    .C(\as2650.addr_buff[2] ),
    .X(_1681_));
 sky130_fd_sc_hd__nand2_1 _4908_ (.A(_1680_),
    .B(_1681_),
    .Y(_1682_));
 sky130_fd_sc_hd__nor2_1 _4909_ (.A(net73),
    .B(_1622_),
    .Y(_1683_));
 sky130_fd_sc_hd__a31o_1 _4910_ (.A1(net296),
    .A2(net295),
    .A3(_1680_),
    .B1(_0684_),
    .X(_1684_));
 sky130_fd_sc_hd__a31o_1 _4911_ (.A1(net296),
    .A2(net295),
    .A3(_1622_),
    .B1(net73),
    .X(_1685_));
 sky130_fd_sc_hd__a21o_1 _4912_ (.A1(_1684_),
    .A2(_1685_),
    .B1(\as2650.addr_buff[2] ),
    .X(_1686_));
 sky130_fd_sc_hd__o31ai_2 _4913_ (.A1(_0684_),
    .A2(_1682_),
    .A3(_1683_),
    .B1(_1686_),
    .Y(_1687_));
 sky130_fd_sc_hd__a22o_1 _4914_ (.A1(net91),
    .A2(_1679_),
    .B1(_1687_),
    .B2(_0720_),
    .X(_1688_));
 sky130_fd_sc_hd__nand2_1 _4915_ (.A(net266),
    .B(net328),
    .Y(_1689_));
 sky130_fd_sc_hd__or2_1 _4916_ (.A(net266),
    .B(net328),
    .X(_1690_));
 sky130_fd_sc_hd__nand2_2 _4917_ (.A(_1689_),
    .B(_1690_),
    .Y(_1691_));
 sky130_fd_sc_hd__inv_2 _4918_ (.A(_1691_),
    .Y(_1692_));
 sky130_fd_sc_hd__o21ai_2 _4919_ (.A1(net267),
    .A2(net268),
    .B1(net329),
    .Y(_1693_));
 sky130_fd_sc_hd__or2_2 _4920_ (.A(_1636_),
    .B(_1661_),
    .X(_1694_));
 sky130_fd_sc_hd__inv_2 _4921_ (.A(_1694_),
    .Y(_1695_));
 sky130_fd_sc_hd__a21oi_1 _4922_ (.A1(_1693_),
    .A2(_1694_),
    .B1(_1691_),
    .Y(_1696_));
 sky130_fd_sc_hd__a31o_1 _4923_ (.A1(_1691_),
    .A2(_1693_),
    .A3(_1694_),
    .B1(net85),
    .X(_1697_));
 sky130_fd_sc_hd__o211a_1 _4924_ (.A1(_1696_),
    .A2(_1697_),
    .B1(net53),
    .C1(net88),
    .X(_1698_));
 sky130_fd_sc_hd__o21ai_1 _4925_ (.A1(net86),
    .A2(_1688_),
    .B1(_1698_),
    .Y(_1699_));
 sky130_fd_sc_hd__or2_1 _4926_ (.A(_1643_),
    .B(_1661_),
    .X(_1700_));
 sky130_fd_sc_hd__inv_2 _4927_ (.A(_1700_),
    .Y(_1701_));
 sky130_fd_sc_hd__a21o_1 _4928_ (.A1(_1693_),
    .A2(_1700_),
    .B1(_1691_),
    .X(_1702_));
 sky130_fd_sc_hd__or3b_1 _4929_ (.A(_1692_),
    .B(_1701_),
    .C_N(_1693_),
    .X(_1703_));
 sky130_fd_sc_hd__nand2_1 _4930_ (.A(_1702_),
    .B(_1703_),
    .Y(_1704_));
 sky130_fd_sc_hd__nand2_1 _4931_ (.A(net324),
    .B(_1704_),
    .Y(_1705_));
 sky130_fd_sc_hd__o2111a_1 _4932_ (.A1(net21),
    .A2(net324),
    .B1(_1331_),
    .C1(_1705_),
    .D1(net229),
    .X(_1706_));
 sky130_fd_sc_hd__o211ai_2 _4933_ (.A1(\as2650.addr_buff[2] ),
    .A2(_1383_),
    .B1(_2603_),
    .C1(net148),
    .Y(_1707_));
 sky130_fd_sc_hd__a221o_1 _4934_ (.A1(_2539_),
    .A2(_2615_),
    .B1(_1679_),
    .B2(net123),
    .C1(_1707_),
    .X(_1708_));
 sky130_fd_sc_hd__o211ai_1 _4935_ (.A1(_2531_),
    .A2(_1339_),
    .B1(_1708_),
    .C1(net59),
    .Y(_1709_));
 sky130_fd_sc_hd__o221a_1 _4936_ (.A1(net266),
    .A2(net52),
    .B1(_1706_),
    .B2(_1709_),
    .C1(_1699_),
    .X(_1710_));
 sky130_fd_sc_hd__or2_1 _4937_ (.A(net21),
    .B(net40),
    .X(_1711_));
 sky130_fd_sc_hd__o311a_1 _4938_ (.A1(_1319_),
    .A2(_1325_),
    .A3(_1710_),
    .B1(_1711_),
    .C1(net318),
    .X(_0183_));
 sky130_fd_sc_hd__o31ai_1 _4939_ (.A1(_0684_),
    .A2(_1682_),
    .A3(_1683_),
    .B1(\as2650.addr_buff[3] ),
    .Y(_1712_));
 sky130_fd_sc_hd__nand2_1 _4940_ (.A(_1622_),
    .B(_1681_),
    .Y(_1713_));
 sky130_fd_sc_hd__a221o_1 _4941_ (.A1(_0685_),
    .A2(_1682_),
    .B1(_1713_),
    .B2(net74),
    .C1(\as2650.addr_buff[3] ),
    .X(_1714_));
 sky130_fd_sc_hd__nor2_1 _4942_ (.A(_2538_),
    .B(_1677_),
    .Y(_1715_));
 sky130_fd_sc_hd__and2_1 _4943_ (.A(_2538_),
    .B(_1677_),
    .X(_1716_));
 sky130_fd_sc_hd__or2_1 _4944_ (.A(_1715_),
    .B(_1716_),
    .X(_1717_));
 sky130_fd_sc_hd__a32o_1 _4945_ (.A1(_0720_),
    .A2(_1712_),
    .A3(_1714_),
    .B1(_1717_),
    .B2(net91),
    .X(_1718_));
 sky130_fd_sc_hd__xor2_4 _4946_ (.A(net265),
    .B(net329),
    .X(_1719_));
 sky130_fd_sc_hd__a21o_1 _4947_ (.A1(net266),
    .A2(net329),
    .B1(_1696_),
    .X(_1720_));
 sky130_fd_sc_hd__xnor2_1 _4948_ (.A(_1719_),
    .B(_1720_),
    .Y(_1721_));
 sky130_fd_sc_hd__mux2_1 _4949_ (.A0(_1718_),
    .A1(_1721_),
    .S(net87),
    .X(_1722_));
 sky130_fd_sc_hd__nor2_1 _4950_ (.A(net128),
    .B(_1717_),
    .Y(_1723_));
 sky130_fd_sc_hd__a221o_1 _4951_ (.A1(net22),
    .A2(_2615_),
    .B1(_1382_),
    .B2(\as2650.addr_buff[3] ),
    .C1(net149),
    .X(_1724_));
 sky130_fd_sc_hd__o22a_1 _4952_ (.A1(net265),
    .A2(net84),
    .B1(_1723_),
    .B2(_1724_),
    .X(_1725_));
 sky130_fd_sc_hd__o22a_1 _4953_ (.A1(net265),
    .A2(net50),
    .B1(_1725_),
    .B2(net75),
    .X(_1726_));
 sky130_fd_sc_hd__nor2_1 _4954_ (.A(net202),
    .B(_1726_),
    .Y(_1727_));
 sky130_fd_sc_hd__nand2_1 _4955_ (.A(_1689_),
    .B(_1702_),
    .Y(_1728_));
 sky130_fd_sc_hd__xor2_2 _4956_ (.A(_1719_),
    .B(_1728_),
    .X(_1729_));
 sky130_fd_sc_hd__nand2_1 _4957_ (.A(net325),
    .B(_1729_),
    .Y(_1730_));
 sky130_fd_sc_hd__o2111a_1 _4958_ (.A1(_2538_),
    .A2(net325),
    .B1(net162),
    .C1(_1390_),
    .D1(_1730_),
    .X(_1731_));
 sky130_fd_sc_hd__a211o_1 _4959_ (.A1(net53),
    .A2(_1722_),
    .B1(_1727_),
    .C1(_1731_),
    .X(_1732_));
 sky130_fd_sc_hd__a2bb2o_1 _4960_ (.A1_N(net265),
    .A2_N(net52),
    .B1(_1732_),
    .B2(net88),
    .X(_1733_));
 sky130_fd_sc_hd__mux2_1 _4961_ (.A0(_2538_),
    .A1(_1733_),
    .S(net40),
    .X(_1734_));
 sky130_fd_sc_hd__nor2_1 _4962_ (.A(net347),
    .B(_1734_),
    .Y(_0184_));
 sky130_fd_sc_hd__xnor2_1 _4963_ (.A(net24),
    .B(_1715_),
    .Y(_1735_));
 sky130_fd_sc_hd__nand2_4 _4964_ (.A(\as2650.addr_buff[3] ),
    .B(_1681_),
    .Y(_1736_));
 sky130_fd_sc_hd__nor2_1 _4965_ (.A(_1617_),
    .B(_1736_),
    .Y(_1737_));
 sky130_fd_sc_hd__xnor2_1 _4966_ (.A(\as2650.addr_buff[4] ),
    .B(_1737_),
    .Y(_1738_));
 sky130_fd_sc_hd__a211o_1 _4967_ (.A1(_1588_),
    .A2(_1589_),
    .B1(_1621_),
    .C1(_1736_),
    .X(_1739_));
 sky130_fd_sc_hd__nand2_1 _4968_ (.A(\as2650.addr_buff[4] ),
    .B(_1739_),
    .Y(_1740_));
 sky130_fd_sc_hd__or2_1 _4969_ (.A(\as2650.addr_buff[4] ),
    .B(_1739_),
    .X(_1741_));
 sky130_fd_sc_hd__a32o_1 _4970_ (.A1(net74),
    .A2(_1740_),
    .A3(_1741_),
    .B1(_0686_),
    .B2(_1738_),
    .X(_1742_));
 sky130_fd_sc_hd__a22o_1 _4971_ (.A1(_0682_),
    .A2(_1735_),
    .B1(_1742_),
    .B2(_0720_),
    .X(_1743_));
 sky130_fd_sc_hd__xnor2_4 _4972_ (.A(net264),
    .B(net329),
    .Y(_1744_));
 sky130_fd_sc_hd__o41a_1 _4973_ (.A1(net265),
    .A2(net266),
    .A3(net267),
    .A4(net268),
    .B1(net329),
    .X(_1745_));
 sky130_fd_sc_hd__a31o_1 _4974_ (.A1(_1692_),
    .A2(_1695_),
    .A3(_1719_),
    .B1(_1745_),
    .X(_1746_));
 sky130_fd_sc_hd__xor2_1 _4975_ (.A(_1744_),
    .B(_1746_),
    .X(_1747_));
 sky130_fd_sc_hd__mux2_1 _4976_ (.A0(_1743_),
    .A1(_1747_),
    .S(net87),
    .X(_1748_));
 sky130_fd_sc_hd__nor2_1 _4977_ (.A(net128),
    .B(_1735_),
    .Y(_1749_));
 sky130_fd_sc_hd__a221o_1 _4978_ (.A1(net24),
    .A2(_2615_),
    .B1(_1382_),
    .B2(\as2650.addr_buff[4] ),
    .C1(net149),
    .X(_1750_));
 sky130_fd_sc_hd__o22a_1 _4979_ (.A1(net264),
    .A2(net84),
    .B1(_1749_),
    .B2(_1750_),
    .X(_1751_));
 sky130_fd_sc_hd__o22a_1 _4980_ (.A1(net264),
    .A2(net50),
    .B1(_1751_),
    .B2(net75),
    .X(_1752_));
 sky130_fd_sc_hd__a31o_2 _4981_ (.A1(_1692_),
    .A2(_1701_),
    .A3(_1719_),
    .B1(_1745_),
    .X(_1753_));
 sky130_fd_sc_hd__xnor2_4 _4982_ (.A(_1744_),
    .B(_1753_),
    .Y(_1754_));
 sky130_fd_sc_hd__a21bo_1 _4983_ (.A1(net24),
    .A2(net310),
    .B1_N(_1390_),
    .X(_1755_));
 sky130_fd_sc_hd__a211o_1 _4984_ (.A1(net325),
    .A2(_1754_),
    .B1(_1755_),
    .C1(net193),
    .X(_1756_));
 sky130_fd_sc_hd__o21ai_1 _4985_ (.A1(net202),
    .A2(_1752_),
    .B1(_1756_),
    .Y(_1757_));
 sky130_fd_sc_hd__a21oi_1 _4986_ (.A1(net53),
    .A2(_1748_),
    .B1(_1757_),
    .Y(_1758_));
 sky130_fd_sc_hd__o22a_1 _4987_ (.A1(net264),
    .A2(net52),
    .B1(_1758_),
    .B2(net90),
    .X(_1759_));
 sky130_fd_sc_hd__or2_1 _4988_ (.A(net24),
    .B(net40),
    .X(_1760_));
 sky130_fd_sc_hd__o311a_1 _4989_ (.A1(_1319_),
    .A2(net42),
    .A3(_1759_),
    .B1(_1760_),
    .C1(net318),
    .X(_0185_));
 sky130_fd_sc_hd__a21o_1 _4990_ (.A1(_2774_),
    .A2(_0660_),
    .B1(_1298_),
    .X(_1761_));
 sky130_fd_sc_hd__or2_1 _4991_ (.A(_0803_),
    .B(_1290_),
    .X(_1762_));
 sky130_fd_sc_hd__or4_1 _4992_ (.A(net204),
    .B(net79),
    .C(_0696_),
    .D(_1313_),
    .X(_1763_));
 sky130_fd_sc_hd__or4_1 _4993_ (.A(_0719_),
    .B(_0731_),
    .C(_1286_),
    .D(_1294_),
    .X(_1764_));
 sky130_fd_sc_hd__or4b_2 _4994_ (.A(_0708_),
    .B(_1761_),
    .C(_1764_),
    .D_N(_1763_),
    .X(_1765_));
 sky130_fd_sc_hd__a211o_1 _4995_ (.A1(net121),
    .A2(_2611_),
    .B1(_2810_),
    .C1(_1762_),
    .X(_1766_));
 sky130_fd_sc_hd__or4b_2 _4996_ (.A(_1297_),
    .B(_1318_),
    .C(_1766_),
    .D_N(_0706_),
    .X(_1767_));
 sky130_fd_sc_hd__nor3_4 _4997_ (.A(_1316_),
    .B(_1765_),
    .C(_1767_),
    .Y(_1768_));
 sky130_fd_sc_hd__a21o_1 _4998_ (.A1(_1324_),
    .A2(_1768_),
    .B1(net25),
    .X(_1769_));
 sky130_fd_sc_hd__a31o_1 _4999_ (.A1(net228),
    .A2(net134),
    .A3(_2682_),
    .B1(net11),
    .X(_1770_));
 sky130_fd_sc_hd__a211o_1 _5000_ (.A1(_2692_),
    .A2(_1770_),
    .B1(_0716_),
    .C1(net80),
    .X(_1771_));
 sky130_fd_sc_hd__o31a_1 _5001_ (.A1(net230),
    .A2(net141),
    .A3(_0715_),
    .B1(_1771_),
    .X(_1772_));
 sky130_fd_sc_hd__o211ai_1 _5002_ (.A1(net90),
    .A2(_1772_),
    .B1(_1768_),
    .C1(_1324_),
    .Y(_1773_));
 sky130_fd_sc_hd__and3_1 _5003_ (.A(net316),
    .B(_1769_),
    .C(_1773_),
    .X(_0186_));
 sky130_fd_sc_hd__and3_1 _5004_ (.A(net325),
    .B(_2603_),
    .C(net116),
    .X(_1774_));
 sky130_fd_sc_hd__nor2_1 _5005_ (.A(_1313_),
    .B(net83),
    .Y(_1775_));
 sky130_fd_sc_hd__o21a_1 _5006_ (.A1(_1774_),
    .A2(_1775_),
    .B1(net225),
    .X(_1776_));
 sky130_fd_sc_hd__and3_1 _5007_ (.A(net225),
    .B(net164),
    .C(_2603_),
    .X(_1777_));
 sky130_fd_sc_hd__a21oi_1 _5008_ (.A1(net163),
    .A2(_2594_),
    .B1(net134),
    .Y(_1778_));
 sky130_fd_sc_hd__and3_1 _5009_ (.A(_1256_),
    .B(_1777_),
    .C(_1778_),
    .X(_1779_));
 sky130_fd_sc_hd__a41o_1 _5010_ (.A1(_2537_),
    .A2(net291),
    .A3(net136),
    .A4(_2594_),
    .B1(_1779_),
    .X(_1780_));
 sky130_fd_sc_hd__a311o_1 _5011_ (.A1(net228),
    .A2(_2565_),
    .A3(net121),
    .B1(_1761_),
    .C1(_1780_),
    .X(_1781_));
 sky130_fd_sc_hd__or2_1 _5012_ (.A(net293),
    .B(_2810_),
    .X(_1782_));
 sky130_fd_sc_hd__nand2_4 _5013_ (.A(net149),
    .B(net135),
    .Y(_1783_));
 sky130_fd_sc_hd__and3_1 _5014_ (.A(\as2650.cycle[0] ),
    .B(net150),
    .C(net136),
    .X(_1784_));
 sky130_fd_sc_hd__or4_1 _5015_ (.A(_2580_),
    .B(_1297_),
    .C(_1782_),
    .D(_1784_),
    .X(_1785_));
 sky130_fd_sc_hd__or4b_1 _5016_ (.A(_1290_),
    .B(_1781_),
    .C(_1785_),
    .D_N(_1314_),
    .X(_1786_));
 sky130_fd_sc_hd__or4_2 _5017_ (.A(_1286_),
    .B(_1294_),
    .C(_1776_),
    .D(_1786_),
    .X(_1787_));
 sky130_fd_sc_hd__nor2_1 _5018_ (.A(net42),
    .B(_1787_),
    .Y(_1788_));
 sky130_fd_sc_hd__a41o_1 _5019_ (.A1(net26),
    .A2(net124),
    .A3(_2607_),
    .A4(net118),
    .B1(_0694_),
    .X(_1789_));
 sky130_fd_sc_hd__nand2_1 _5020_ (.A(net134),
    .B(_2607_),
    .Y(_1790_));
 sky130_fd_sc_hd__a31o_1 _5021_ (.A1(net134),
    .A2(net124),
    .A3(_2607_),
    .B1(_1382_),
    .X(_1791_));
 sky130_fd_sc_hd__and4_1 _5022_ (.A(net26),
    .B(_2602_),
    .C(net117),
    .D(_1791_),
    .X(_1792_));
 sky130_fd_sc_hd__nor2_1 _5023_ (.A(net310),
    .B(_2602_),
    .Y(_1793_));
 sky130_fd_sc_hd__a311o_1 _5024_ (.A1(net26),
    .A2(net118),
    .A3(_0715_),
    .B1(net230),
    .C1(net79),
    .X(_1794_));
 sky130_fd_sc_hd__or3b_1 _5025_ (.A(_1792_),
    .B(_1793_),
    .C_N(net50),
    .X(_1795_));
 sky130_fd_sc_hd__a21o_1 _5026_ (.A1(_1794_),
    .A2(_1795_),
    .B1(net202),
    .X(_1796_));
 sky130_fd_sc_hd__a31o_1 _5027_ (.A1(_0712_),
    .A2(_1789_),
    .A3(_1796_),
    .B1(net90),
    .X(_1797_));
 sky130_fd_sc_hd__mux2_1 _5028_ (.A0(net26),
    .A1(_1797_),
    .S(_1788_),
    .X(_1798_));
 sky130_fd_sc_hd__and2_1 _5029_ (.A(net318),
    .B(_1798_),
    .X(_0187_));
 sky130_fd_sc_hd__o31ai_4 _5030_ (.A1(net80),
    .A2(net74),
    .A3(_0690_),
    .B1(net203),
    .Y(_1799_));
 sky130_fd_sc_hd__a211oi_4 _5031_ (.A1(_0697_),
    .A2(_1799_),
    .B1(_1306_),
    .C1(net292),
    .Y(_1800_));
 sky130_fd_sc_hd__a21bo_1 _5032_ (.A1(\as2650.addr_buff[5] ),
    .A2(net88),
    .B1_N(_1800_),
    .X(_1801_));
 sky130_fd_sc_hd__o211a_1 _5033_ (.A1(\as2650.idx_ctrl[0] ),
    .A2(_1800_),
    .B1(_1801_),
    .C1(net316),
    .X(_0188_));
 sky130_fd_sc_hd__a21bo_1 _5034_ (.A1(\as2650.addr_buff[6] ),
    .A2(_0699_),
    .B1_N(_1800_),
    .X(_1802_));
 sky130_fd_sc_hd__o211a_1 _5035_ (.A1(\as2650.idx_ctrl[1] ),
    .A2(_1800_),
    .B1(_1802_),
    .C1(net316),
    .X(_0189_));
 sky130_fd_sc_hd__a32o_1 _5036_ (.A1(net81),
    .A2(net201),
    .A3(_0775_),
    .B1(_1291_),
    .B2(net118),
    .X(_1803_));
 sky130_fd_sc_hd__a2bb2o_1 _5037_ (.A1_N(_2692_),
    .A2_N(_1292_),
    .B1(_0797_),
    .B2(net62),
    .X(_1804_));
 sky130_fd_sc_hd__or3_4 _5038_ (.A(_2674_),
    .B(_1803_),
    .C(_1804_),
    .X(_1805_));
 sky130_fd_sc_hd__and3_2 _5039_ (.A(net260),
    .B(net165),
    .C(net163),
    .X(_1806_));
 sky130_fd_sc_hd__a21o_1 _5040_ (.A1(net350),
    .A2(net145),
    .B1(_1806_),
    .X(_1807_));
 sky130_fd_sc_hd__mux2_1 _5041_ (.A0(_1807_),
    .A1(\as2650.holding_reg[0] ),
    .S(_1805_),
    .X(_0190_));
 sky130_fd_sc_hd__nand2_2 _5042_ (.A(_2550_),
    .B(net147),
    .Y(_1808_));
 sky130_fd_sc_hd__nor2_1 _5043_ (.A(net257),
    .B(net145),
    .Y(_1809_));
 sky130_fd_sc_hd__or3b_1 _5044_ (.A(_1809_),
    .B(_1805_),
    .C_N(_1808_),
    .X(_1810_));
 sky130_fd_sc_hd__a21bo_1 _5045_ (.A1(\as2650.holding_reg[1] ),
    .A2(_1805_),
    .B1_N(_1810_),
    .X(_0191_));
 sky130_fd_sc_hd__and3_1 _5046_ (.A(net253),
    .B(net165),
    .C(net163),
    .X(_1811_));
 sky130_fd_sc_hd__a21o_1 _5047_ (.A1(net343),
    .A2(net144),
    .B1(_1811_),
    .X(_1812_));
 sky130_fd_sc_hd__mux2_1 _5048_ (.A0(_1812_),
    .A1(\as2650.holding_reg[2] ),
    .S(_1805_),
    .X(_0192_));
 sky130_fd_sc_hd__and3_2 _5049_ (.A(net248),
    .B(_2564_),
    .C(_2566_),
    .X(_1813_));
 sky130_fd_sc_hd__a21o_1 _5050_ (.A1(net339),
    .A2(net144),
    .B1(_1813_),
    .X(_1814_));
 sky130_fd_sc_hd__mux2_1 _5051_ (.A0(_1814_),
    .A1(\as2650.holding_reg[3] ),
    .S(_1805_),
    .X(_0193_));
 sky130_fd_sc_hd__and3_2 _5052_ (.A(net245),
    .B(_2564_),
    .C(_2566_),
    .X(_1815_));
 sky130_fd_sc_hd__a21o_1 _5053_ (.A1(net336),
    .A2(net144),
    .B1(_1815_),
    .X(_1816_));
 sky130_fd_sc_hd__mux2_1 _5054_ (.A0(_1816_),
    .A1(\as2650.holding_reg[4] ),
    .S(_1805_),
    .X(_0194_));
 sky130_fd_sc_hd__a21o_1 _5055_ (.A1(net333),
    .A2(net145),
    .B1(_0673_),
    .X(_1817_));
 sky130_fd_sc_hd__mux2_1 _5056_ (.A0(_1817_),
    .A1(\as2650.holding_reg[5] ),
    .S(_1805_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _5057_ (.A0(net238),
    .A1(net7),
    .S(net144),
    .X(_1818_));
 sky130_fd_sc_hd__mux2_1 _5058_ (.A0(_1818_),
    .A1(\as2650.holding_reg[6] ),
    .S(_1805_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _5059_ (.A0(net234),
    .A1(net327),
    .S(net144),
    .X(_1819_));
 sky130_fd_sc_hd__mux2_1 _5060_ (.A0(_1819_),
    .A1(\as2650.holding_reg[7] ),
    .S(_1805_),
    .X(_0197_));
 sky130_fd_sc_hd__nor2_1 _5061_ (.A(net347),
    .B(_0804_),
    .Y(_0198_));
 sky130_fd_sc_hd__or2_1 _5062_ (.A(net290),
    .B(_2594_),
    .X(_1820_));
 sky130_fd_sc_hd__and2_4 _5063_ (.A(_1312_),
    .B(_1323_),
    .X(_1821_));
 sky130_fd_sc_hd__and3_2 _5064_ (.A(net77),
    .B(_1312_),
    .C(_1323_),
    .X(_1822_));
 sky130_fd_sc_hd__nand2_4 _5065_ (.A(net77),
    .B(_1821_),
    .Y(_1823_));
 sky130_fd_sc_hd__or2_1 _5066_ (.A(net291),
    .B(net150),
    .X(_1824_));
 sky130_fd_sc_hd__o211a_1 _5067_ (.A1(net128),
    .A2(_1824_),
    .B1(_1823_),
    .C1(net134),
    .X(_1825_));
 sky130_fd_sc_hd__a31o_1 _5068_ (.A1(net136),
    .A2(_1383_),
    .A3(_1820_),
    .B1(_1825_),
    .X(_1826_));
 sky130_fd_sc_hd__or4_2 _5069_ (.A(_2808_),
    .B(_0633_),
    .C(_0656_),
    .D(_0659_),
    .X(_1827_));
 sky130_fd_sc_hd__a2bb2o_1 _5070_ (.A1_N(net124),
    .A2_N(_0715_),
    .B1(_1824_),
    .B2(_1827_),
    .X(_1828_));
 sky130_fd_sc_hd__nand2_1 _5071_ (.A(_0636_),
    .B(_0668_),
    .Y(_1829_));
 sky130_fd_sc_hd__o21a_1 _5072_ (.A1(net92),
    .A2(_1824_),
    .B1(net207),
    .X(_1830_));
 sky130_fd_sc_hd__a32o_1 _5073_ (.A1(_1828_),
    .A2(_1829_),
    .A3(_1830_),
    .B1(_1826_),
    .B2(_2603_),
    .X(_1831_));
 sky130_fd_sc_hd__a22o_1 _5074_ (.A1(net290),
    .A2(net121),
    .B1(_0697_),
    .B2(_1831_),
    .X(_1832_));
 sky130_fd_sc_hd__a21oi_1 _5075_ (.A1(_2652_),
    .A2(_0707_),
    .B1(_2670_),
    .Y(_1833_));
 sky130_fd_sc_hd__nand2_1 _5076_ (.A(net312),
    .B(_2652_),
    .Y(_1834_));
 sky130_fd_sc_hd__a221o_1 _5077_ (.A1(net291),
    .A2(_2670_),
    .B1(net87),
    .B2(_1834_),
    .C1(_1833_),
    .X(_1835_));
 sky130_fd_sc_hd__or4b_1 _5078_ (.A(net79),
    .B(net131),
    .C(_1835_),
    .D_N(_1277_),
    .X(_1836_));
 sky130_fd_sc_hd__or2_2 _5079_ (.A(net208),
    .B(_0805_),
    .X(_1837_));
 sky130_fd_sc_hd__and4_1 _5080_ (.A(net203),
    .B(_0697_),
    .C(_1836_),
    .D(_1837_),
    .X(_1838_));
 sky130_fd_sc_hd__a211o_1 _5081_ (.A1(net222),
    .A2(_1832_),
    .B1(_0711_),
    .C1(net292),
    .X(_1839_));
 sky130_fd_sc_hd__o2bb2a_1 _5082_ (.A1_N(net292),
    .A2_N(net291),
    .B1(_1838_),
    .B2(_1839_),
    .X(_1840_));
 sky130_fd_sc_hd__nor2_1 _5083_ (.A(net347),
    .B(_1840_),
    .Y(_0199_));
 sky130_fd_sc_hd__nand2_2 _5084_ (.A(_2535_),
    .B(net88),
    .Y(_1841_));
 sky130_fd_sc_hd__a311o_1 _5085_ (.A1(net303),
    .A2(net163),
    .A3(_2594_),
    .B1(_1305_),
    .C1(_2590_),
    .X(_1842_));
 sky130_fd_sc_hd__or2_1 _5086_ (.A(net150),
    .B(_1305_),
    .X(_1843_));
 sky130_fd_sc_hd__o221a_1 _5087_ (.A1(net137),
    .A2(_1823_),
    .B1(_1843_),
    .B2(_1790_),
    .C1(_1842_),
    .X(_1844_));
 sky130_fd_sc_hd__o21a_1 _5088_ (.A1(_1305_),
    .A2(_1833_),
    .B1(net85),
    .X(_1845_));
 sky130_fd_sc_hd__a21o_1 _5089_ (.A1(net87),
    .A2(_1834_),
    .B1(_1845_),
    .X(_1846_));
 sky130_fd_sc_hd__or3b_1 _5090_ (.A(net79),
    .B(_1846_),
    .C_N(_2607_),
    .X(_1847_));
 sky130_fd_sc_hd__a21o_1 _5091_ (.A1(_1837_),
    .A2(_1847_),
    .B1(net222),
    .X(_1848_));
 sky130_fd_sc_hd__o211a_1 _5092_ (.A1(net141),
    .A2(_1827_),
    .B1(_1829_),
    .C1(_1843_),
    .X(_1849_));
 sky130_fd_sc_hd__o211a_1 _5093_ (.A1(net151),
    .A2(_1849_),
    .B1(_1848_),
    .C1(_0697_),
    .X(_1850_));
 sky130_fd_sc_hd__o21a_1 _5094_ (.A1(net193),
    .A2(_1844_),
    .B1(_1850_),
    .X(_1851_));
 sky130_fd_sc_hd__o22a_1 _5095_ (.A1(_2535_),
    .A2(_2537_),
    .B1(_1841_),
    .B2(_1851_),
    .X(_1852_));
 sky130_fd_sc_hd__nor2_1 _5096_ (.A(net347),
    .B(_1852_),
    .Y(_0200_));
 sky130_fd_sc_hd__and3_2 _5097_ (.A(net289),
    .B(\as2650.cycle[1] ),
    .C(net290),
    .X(_1853_));
 sky130_fd_sc_hd__a21oi_1 _5098_ (.A1(\as2650.cycle[1] ),
    .A2(net290),
    .B1(net289),
    .Y(_1854_));
 sky130_fd_sc_hd__or3_2 _5099_ (.A(net131),
    .B(_1853_),
    .C(_1854_),
    .X(_1855_));
 sky130_fd_sc_hd__o31ai_1 _5100_ (.A1(net141),
    .A2(net197),
    .A3(_0807_),
    .B1(_1855_),
    .Y(_1856_));
 sky130_fd_sc_hd__a211o_1 _5101_ (.A1(_2612_),
    .A2(net56),
    .B1(_1853_),
    .C1(_1854_),
    .X(_1857_));
 sky130_fd_sc_hd__a21oi_1 _5102_ (.A1(net126),
    .A2(net118),
    .B1(_0715_),
    .Y(_1858_));
 sky130_fd_sc_hd__or4_1 _5103_ (.A(net288),
    .B(net289),
    .C(_2608_),
    .D(net92),
    .X(_1859_));
 sky130_fd_sc_hd__xnor2_1 _5104_ (.A(_1857_),
    .B(_1858_),
    .Y(_1860_));
 sky130_fd_sc_hd__or3b_1 _5105_ (.A(net231),
    .B(_1860_),
    .C_N(_1859_),
    .X(_1861_));
 sky130_fd_sc_hd__a311o_1 _5106_ (.A1(net163),
    .A2(net136),
    .A3(_2594_),
    .B1(net116),
    .C1(_1855_),
    .X(_1862_));
 sky130_fd_sc_hd__and3_1 _5107_ (.A(net294),
    .B(net136),
    .C(net130),
    .X(_1863_));
 sky130_fd_sc_hd__o21ai_1 _5108_ (.A1(_2595_),
    .A2(net119),
    .B1(_1862_),
    .Y(_1864_));
 sky130_fd_sc_hd__o311a_1 _5109_ (.A1(net207),
    .A2(_1863_),
    .A3(_1864_),
    .B1(net222),
    .C1(_1861_),
    .X(_1865_));
 sky130_fd_sc_hd__a211o_1 _5110_ (.A1(net203),
    .A2(_1856_),
    .B1(_1865_),
    .C1(_1841_),
    .X(_1866_));
 sky130_fd_sc_hd__a21o_1 _5111_ (.A1(_2535_),
    .A2(_0699_),
    .B1(net289),
    .X(_1867_));
 sky130_fd_sc_hd__and3_1 _5112_ (.A(net316),
    .B(_1866_),
    .C(_1867_),
    .X(_0201_));
 sky130_fd_sc_hd__nor2_1 _5113_ (.A(net288),
    .B(_1853_),
    .Y(_1868_));
 sky130_fd_sc_hd__and2_2 _5114_ (.A(net288),
    .B(_1853_),
    .X(_1869_));
 sky130_fd_sc_hd__nor2_2 _5115_ (.A(_1868_),
    .B(_1869_),
    .Y(_1870_));
 sky130_fd_sc_hd__a21o_1 _5116_ (.A1(net124),
    .A2(_2607_),
    .B1(net137),
    .X(_1871_));
 sky130_fd_sc_hd__a21o_1 _5117_ (.A1(_2627_),
    .A2(_1871_),
    .B1(net206),
    .X(_1872_));
 sky130_fd_sc_hd__a31o_1 _5118_ (.A1(net230),
    .A2(_2590_),
    .A3(_1382_),
    .B1(_1774_),
    .X(_1873_));
 sky130_fd_sc_hd__nand3_1 _5119_ (.A(_2673_),
    .B(_2685_),
    .C(net85),
    .Y(_1874_));
 sky130_fd_sc_hd__a31o_1 _5120_ (.A1(_2651_),
    .A2(_0704_),
    .A3(_1874_),
    .B1(_1870_),
    .X(_1875_));
 sky130_fd_sc_hd__a221o_1 _5121_ (.A1(_2609_),
    .A2(_1793_),
    .B1(_1870_),
    .B2(_1872_),
    .C1(_1873_),
    .X(_1876_));
 sky130_fd_sc_hd__a41o_1 _5122_ (.A1(net203),
    .A2(_2607_),
    .A3(_1277_),
    .A4(_1875_),
    .B1(net292),
    .X(_1877_));
 sky130_fd_sc_hd__a21o_1 _5123_ (.A1(net222),
    .A2(_1876_),
    .B1(_1877_),
    .X(_1878_));
 sky130_fd_sc_hd__o211a_1 _5124_ (.A1(_2535_),
    .A2(net288),
    .B1(net316),
    .C1(_1878_),
    .X(_0202_));
 sky130_fd_sc_hd__a21oi_1 _5125_ (.A1(_2535_),
    .A2(_1869_),
    .B1(\as2650.cycle[4] ),
    .Y(_1879_));
 sky130_fd_sc_hd__and3_1 _5126_ (.A(_2535_),
    .B(\as2650.cycle[4] ),
    .C(_1869_),
    .X(_1880_));
 sky130_fd_sc_hd__nor3_1 _5127_ (.A(net347),
    .B(_1879_),
    .C(_1880_),
    .Y(_0203_));
 sky130_fd_sc_hd__a21oi_1 _5128_ (.A1(\as2650.cycle[5] ),
    .A2(_1880_),
    .B1(net347),
    .Y(_1881_));
 sky130_fd_sc_hd__o21a_1 _5129_ (.A1(\as2650.cycle[5] ),
    .A2(_1880_),
    .B1(_1881_),
    .X(_0204_));
 sky130_fd_sc_hd__and4_1 _5130_ (.A(\as2650.cycle[6] ),
    .B(\as2650.cycle[5] ),
    .C(\as2650.cycle[4] ),
    .D(_1869_),
    .X(_1882_));
 sky130_fd_sc_hd__a31o_1 _5131_ (.A1(\as2650.cycle[5] ),
    .A2(\as2650.cycle[4] ),
    .A3(_1869_),
    .B1(\as2650.cycle[6] ),
    .X(_1883_));
 sky130_fd_sc_hd__a31o_1 _5132_ (.A1(_2673_),
    .A2(_2685_),
    .A3(net85),
    .B1(_0701_),
    .X(_1884_));
 sky130_fd_sc_hd__and3b_1 _5133_ (.A_N(_1882_),
    .B(_1883_),
    .C(_1884_),
    .X(_1885_));
 sky130_fd_sc_hd__a311o_1 _5134_ (.A1(net303),
    .A2(_2689_),
    .A3(_0700_),
    .B1(_0705_),
    .C1(net292),
    .X(_1886_));
 sky130_fd_sc_hd__o221a_1 _5135_ (.A1(_2535_),
    .A2(\as2650.cycle[6] ),
    .B1(_1885_),
    .B2(_1886_),
    .C1(net316),
    .X(_0205_));
 sky130_fd_sc_hd__a31o_1 _5136_ (.A1(net141),
    .A2(net73),
    .A3(_0703_),
    .B1(_0701_),
    .X(_1887_));
 sky130_fd_sc_hd__xnor2_1 _5137_ (.A(_2536_),
    .B(_1882_),
    .Y(_1888_));
 sky130_fd_sc_hd__a221o_1 _5138_ (.A1(net230),
    .A2(net62),
    .B1(_1887_),
    .B2(_1888_),
    .C1(net292),
    .X(_1889_));
 sky130_fd_sc_hd__o211a_1 _5139_ (.A1(_2535_),
    .A2(\as2650.cycle[7] ),
    .B1(net316),
    .C1(_1889_),
    .X(_0206_));
 sky130_fd_sc_hd__nand2_1 _5140_ (.A(_0800_),
    .B(_0806_),
    .Y(_1890_));
 sky130_fd_sc_hd__nor2_1 _5141_ (.A(net311),
    .B(_0674_),
    .Y(_1891_));
 sky130_fd_sc_hd__a211o_1 _5142_ (.A1(\as2650.psu[7] ),
    .A2(net311),
    .B1(_0800_),
    .C1(_1891_),
    .X(_1892_));
 sky130_fd_sc_hd__o22a_1 _5143_ (.A1(net235),
    .A2(_0806_),
    .B1(_1890_),
    .B2(net9),
    .X(_1893_));
 sky130_fd_sc_hd__a21o_1 _5144_ (.A1(_1892_),
    .A2(_1893_),
    .B1(net293),
    .X(_1894_));
 sky130_fd_sc_hd__o211a_1 _5145_ (.A1(\as2650.psu[7] ),
    .A2(_2535_),
    .B1(net319),
    .C1(_1894_),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _5146_ (.A0(_2534_),
    .A1(_1329_),
    .S(net309),
    .X(_1895_));
 sky130_fd_sc_hd__o211a_1 _5147_ (.A1(_2557_),
    .A2(net127),
    .B1(net117),
    .C1(_1332_),
    .X(_1896_));
 sky130_fd_sc_hd__a221o_1 _5148_ (.A1(net285),
    .A2(_1335_),
    .B1(_1895_),
    .B2(net116),
    .C1(_1896_),
    .X(_1897_));
 sky130_fd_sc_hd__a21o_1 _5149_ (.A1(net138),
    .A2(_1897_),
    .B1(net137),
    .X(_1898_));
 sky130_fd_sc_hd__xor2_1 _5150_ (.A(net285),
    .B(net302),
    .X(_1899_));
 sky130_fd_sc_hd__mux2_1 _5151_ (.A0(net285),
    .A1(_1899_),
    .S(_1322_),
    .X(_1900_));
 sky130_fd_sc_hd__mux2_1 _5152_ (.A0(_1899_),
    .A1(net285),
    .S(_1312_),
    .X(_1901_));
 sky130_fd_sc_hd__mux2_1 _5153_ (.A0(_1900_),
    .A1(_1901_),
    .S(_2649_),
    .X(_1902_));
 sky130_fd_sc_hd__a21o_1 _5154_ (.A1(net76),
    .A2(_1902_),
    .B1(_1898_),
    .X(_1903_));
 sky130_fd_sc_hd__nand2_1 _5155_ (.A(net349),
    .B(net122),
    .Y(_1904_));
 sky130_fd_sc_hd__xnor2_2 _5156_ (.A(net349),
    .B(_2703_),
    .Y(_1905_));
 sky130_fd_sc_hd__o2111a_1 _5157_ (.A1(net122),
    .A2(_1905_),
    .B1(_2610_),
    .C1(net139),
    .D1(_1904_),
    .X(_1906_));
 sky130_fd_sc_hd__a211o_1 _5158_ (.A1(net285),
    .A2(net149),
    .B1(net134),
    .C1(_1906_),
    .X(_1907_));
 sky130_fd_sc_hd__and2_1 _5159_ (.A(net140),
    .B(_1895_),
    .X(_1908_));
 sky130_fd_sc_hd__a211o_1 _5160_ (.A1(net285),
    .A2(net76),
    .B1(net119),
    .C1(_1908_),
    .X(_1909_));
 sky130_fd_sc_hd__a31o_1 _5161_ (.A1(_1903_),
    .A2(_1907_),
    .A3(_1909_),
    .B1(net206),
    .X(_1910_));
 sky130_fd_sc_hd__and3_1 _5162_ (.A(net220),
    .B(\as2650.stack[3][0] ),
    .C(net172),
    .X(_1911_));
 sky130_fd_sc_hd__o22a_1 _5163_ (.A1(\as2650.stack[1][0] ),
    .A2(net166),
    .B1(net155),
    .B2(\as2650.stack[0][0] ),
    .X(_1912_));
 sky130_fd_sc_hd__o221a_1 _5164_ (.A1(\as2650.stack[2][0] ),
    .A2(net169),
    .B1(_1911_),
    .B2(net158),
    .C1(_1912_),
    .X(_1913_));
 sky130_fd_sc_hd__mux4_1 _5165_ (.A0(\as2650.stack[7][0] ),
    .A1(\as2650.stack[4][0] ),
    .A2(\as2650.stack[5][0] ),
    .A3(\as2650.stack[6][0] ),
    .S0(net216),
    .S1(net218),
    .X(_1914_));
 sky130_fd_sc_hd__a21o_2 _5166_ (.A1(net107),
    .A2(_1914_),
    .B1(_1913_),
    .X(_1915_));
 sky130_fd_sc_hd__o2bb2a_1 _5167_ (.A1_N(_0717_),
    .A2_N(_1915_),
    .B1(net60),
    .B2(net285),
    .X(_1916_));
 sky130_fd_sc_hd__a21oi_1 _5168_ (.A1(_1910_),
    .A2(_1916_),
    .B1(net57),
    .Y(_1917_));
 sky130_fd_sc_hd__a41o_1 _5169_ (.A1(net141),
    .A2(_0636_),
    .A3(net153),
    .A4(_0697_),
    .B1(_1863_),
    .X(_1918_));
 sky130_fd_sc_hd__or3_1 _5170_ (.A(_1297_),
    .B(_1782_),
    .C(_1918_),
    .X(_1919_));
 sky130_fd_sc_hd__nor3_1 _5171_ (.A(_2572_),
    .B(_0667_),
    .C(_1837_),
    .Y(_1920_));
 sky130_fd_sc_hd__o311a_1 _5172_ (.A1(_2536_),
    .A2(\as2650.cycle[6] ),
    .A3(net222),
    .B1(_2696_),
    .C1(_0714_),
    .X(_1921_));
 sky130_fd_sc_hd__or4b_1 _5173_ (.A(_1303_),
    .B(_1919_),
    .C(_1920_),
    .D_N(_1921_),
    .X(_1922_));
 sky130_fd_sc_hd__or4_1 _5174_ (.A(net207),
    .B(net137),
    .C(_2612_),
    .D(_0709_),
    .X(_1923_));
 sky130_fd_sc_hd__o21ai_1 _5175_ (.A1(_1313_),
    .A2(_1383_),
    .B1(_1923_),
    .Y(_1924_));
 sky130_fd_sc_hd__a211o_1 _5176_ (.A1(net162),
    .A2(_1924_),
    .B1(_1922_),
    .C1(_1781_),
    .X(_1925_));
 sky130_fd_sc_hd__or3_1 _5177_ (.A(net136),
    .B(net128),
    .C(_2606_),
    .X(_1926_));
 sky130_fd_sc_hd__or4_1 _5178_ (.A(net165),
    .B(net194),
    .C(net121),
    .D(_1926_),
    .X(_1927_));
 sky130_fd_sc_hd__or4b_1 _5179_ (.A(_1294_),
    .B(_1307_),
    .C(_1762_),
    .D_N(_1927_),
    .X(_1928_));
 sky130_fd_sc_hd__nor3_2 _5180_ (.A(_1318_),
    .B(_1925_),
    .C(_1928_),
    .Y(_1929_));
 sky130_fd_sc_hd__inv_2 _5181_ (.A(net45),
    .Y(_1930_));
 sky130_fd_sc_hd__a211o_1 _5182_ (.A1(_2534_),
    .A2(net57),
    .B1(_1917_),
    .C1(_1930_),
    .X(_1931_));
 sky130_fd_sc_hd__o211a_1 _5183_ (.A1(net286),
    .A2(net46),
    .B1(_1931_),
    .C1(net313),
    .X(_0208_));
 sky130_fd_sc_hd__xnor2_4 _5184_ (.A(net284),
    .B(net287),
    .Y(_1932_));
 sky130_fd_sc_hd__nand2_4 _5185_ (.A(_1783_),
    .B(_1823_),
    .Y(_1933_));
 sky130_fd_sc_hd__nand2_2 _5186_ (.A(net344),
    .B(_2715_),
    .Y(_1934_));
 sky130_fd_sc_hd__or2_1 _5187_ (.A(net344),
    .B(_2715_),
    .X(_1935_));
 sky130_fd_sc_hd__a22o_1 _5188_ (.A1(net349),
    .A2(_2703_),
    .B1(_1934_),
    .B2(_1935_),
    .X(_1936_));
 sky130_fd_sc_hd__nand4_2 _5189_ (.A(net349),
    .B(_2703_),
    .C(_1934_),
    .D(_1935_),
    .Y(_1937_));
 sky130_fd_sc_hd__and3_1 _5190_ (.A(net129),
    .B(_1936_),
    .C(_1937_),
    .X(_1938_));
 sky130_fd_sc_hd__a211o_1 _5191_ (.A1(net344),
    .A2(net122),
    .B1(_2612_),
    .C1(_1938_),
    .X(_1939_));
 sky130_fd_sc_hd__mux2_1 _5192_ (.A0(net344),
    .A1(net295),
    .S(net123),
    .X(_1940_));
 sky130_fd_sc_hd__mux2_1 _5193_ (.A0(net283),
    .A1(_1387_),
    .S(net309),
    .X(_1941_));
 sky130_fd_sc_hd__o21ai_1 _5194_ (.A1(net83),
    .A2(_1932_),
    .B1(net138),
    .Y(_1942_));
 sky130_fd_sc_hd__a221o_1 _5195_ (.A1(net135),
    .A2(_1939_),
    .B1(_1941_),
    .B2(net116),
    .C1(_1942_),
    .X(_1943_));
 sky130_fd_sc_hd__a21oi_1 _5196_ (.A1(_1257_),
    .A2(_1940_),
    .B1(_1943_),
    .Y(_1944_));
 sky130_fd_sc_hd__o21a_2 _5197_ (.A1(net287),
    .A2(net302),
    .B1(net282),
    .X(_1945_));
 sky130_fd_sc_hd__nor3_1 _5198_ (.A(net283),
    .B(net285),
    .C(net302),
    .Y(_1946_));
 sky130_fd_sc_hd__nor2_8 _5199_ (.A(net138),
    .B(_1821_),
    .Y(_1947_));
 sky130_fd_sc_hd__or2_2 _5200_ (.A(net139),
    .B(_1821_),
    .X(_1948_));
 sky130_fd_sc_hd__o211a_1 _5201_ (.A1(_1945_),
    .A2(_1946_),
    .B1(_1947_),
    .C1(net133),
    .X(_1949_));
 sky130_fd_sc_hd__a211o_1 _5202_ (.A1(_1932_),
    .A2(_1933_),
    .B1(_1944_),
    .C1(_1949_),
    .X(_1950_));
 sky130_fd_sc_hd__nand2_1 _5203_ (.A(net50),
    .B(_1941_),
    .Y(_1951_));
 sky130_fd_sc_hd__or2_1 _5204_ (.A(_2690_),
    .B(_1932_),
    .X(_1952_));
 sky130_fd_sc_hd__a32o_1 _5205_ (.A1(net75),
    .A2(_1951_),
    .A3(_1952_),
    .B1(_1950_),
    .B2(net119),
    .X(_1953_));
 sky130_fd_sc_hd__and3_1 _5206_ (.A(net220),
    .B(\as2650.stack[3][1] ),
    .C(net172),
    .X(_1954_));
 sky130_fd_sc_hd__o22a_1 _5207_ (.A1(\as2650.stack[1][1] ),
    .A2(net166),
    .B1(net155),
    .B2(\as2650.stack[0][1] ),
    .X(_1955_));
 sky130_fd_sc_hd__o221a_2 _5208_ (.A1(\as2650.stack[2][1] ),
    .A2(net169),
    .B1(_1954_),
    .B2(net158),
    .C1(_1955_),
    .X(_1956_));
 sky130_fd_sc_hd__mux4_2 _5209_ (.A0(\as2650.stack[7][1] ),
    .A1(\as2650.stack[4][1] ),
    .A2(\as2650.stack[5][1] ),
    .A3(\as2650.stack[6][1] ),
    .S0(net216),
    .S1(net218),
    .X(_1957_));
 sky130_fd_sc_hd__a21oi_4 _5210_ (.A1(net107),
    .A2(_1957_),
    .B1(_1956_),
    .Y(_1958_));
 sky130_fd_sc_hd__inv_2 _5211_ (.A(_1958_),
    .Y(_1959_));
 sky130_fd_sc_hd__o221a_1 _5212_ (.A1(net60),
    .A2(_1932_),
    .B1(_1958_),
    .B2(net63),
    .C1(_1953_),
    .X(_1960_));
 sky130_fd_sc_hd__nor2_1 _5213_ (.A(net58),
    .B(_1932_),
    .Y(_1961_));
 sky130_fd_sc_hd__o21ai_1 _5214_ (.A1(_1310_),
    .A2(_1960_),
    .B1(net44),
    .Y(_1962_));
 sky130_fd_sc_hd__o221a_1 _5215_ (.A1(net284),
    .A2(net44),
    .B1(_1961_),
    .B2(_1962_),
    .C1(net315),
    .X(_0209_));
 sky130_fd_sc_hd__and3_2 _5216_ (.A(net280),
    .B(net282),
    .C(net286),
    .X(_1963_));
 sky130_fd_sc_hd__a21oi_2 _5217_ (.A1(net282),
    .A2(net286),
    .B1(net281),
    .Y(_1964_));
 sky130_fd_sc_hd__nor2_4 _5218_ (.A(_1963_),
    .B(_1964_),
    .Y(_1965_));
 sky130_fd_sc_hd__mux2_1 _5219_ (.A0(net279),
    .A1(_1423_),
    .S(net309),
    .X(_1966_));
 sky130_fd_sc_hd__and2_1 _5220_ (.A(net138),
    .B(_1966_),
    .X(_1967_));
 sky130_fd_sc_hd__o21a_1 _5221_ (.A1(_2627_),
    .A2(_1966_),
    .B1(net138),
    .X(_1968_));
 sky130_fd_sc_hd__mux2_1 _5222_ (.A0(net341),
    .A1(\as2650.addr_buff[2] ),
    .S(net122),
    .X(_1969_));
 sky130_fd_sc_hd__o22a_1 _5223_ (.A1(net83),
    .A2(_1965_),
    .B1(_1969_),
    .B2(_2612_),
    .X(_1970_));
 sky130_fd_sc_hd__a21o_1 _5224_ (.A1(_1968_),
    .A2(_1970_),
    .B1(net135),
    .X(_1971_));
 sky130_fd_sc_hd__xor2_1 _5225_ (.A(net279),
    .B(_1945_),
    .X(_1972_));
 sky130_fd_sc_hd__a221o_1 _5226_ (.A1(_1822_),
    .A2(_1965_),
    .B1(_1972_),
    .B2(_1947_),
    .C1(_1971_),
    .X(_1973_));
 sky130_fd_sc_hd__and2_1 _5227_ (.A(net341),
    .B(_2823_),
    .X(_1974_));
 sky130_fd_sc_hd__nand2_1 _5228_ (.A(net343),
    .B(_2823_),
    .Y(_1975_));
 sky130_fd_sc_hd__nor2_1 _5229_ (.A(net343),
    .B(_2823_),
    .Y(_1976_));
 sky130_fd_sc_hd__o211ai_1 _5230_ (.A1(_1974_),
    .A2(_1976_),
    .B1(_1934_),
    .C1(_1937_),
    .Y(_1977_));
 sky130_fd_sc_hd__a211o_1 _5231_ (.A1(_1934_),
    .A2(_1937_),
    .B1(_1974_),
    .C1(_1976_),
    .X(_1978_));
 sky130_fd_sc_hd__and3_1 _5232_ (.A(net129),
    .B(_1977_),
    .C(_1978_),
    .X(_1979_));
 sky130_fd_sc_hd__nor2_4 _5233_ (.A(net149),
    .B(net133),
    .Y(_1980_));
 sky130_fd_sc_hd__nand2_1 _5234_ (.A(net148),
    .B(net135),
    .Y(_1981_));
 sky130_fd_sc_hd__a211o_1 _5235_ (.A1(net343),
    .A2(net125),
    .B1(_1979_),
    .C1(_1981_),
    .X(_1982_));
 sky130_fd_sc_hd__or2_1 _5236_ (.A(_1783_),
    .B(_1965_),
    .X(_1983_));
 sky130_fd_sc_hd__a31o_1 _5237_ (.A1(_1973_),
    .A2(_1982_),
    .A3(_1983_),
    .B1(net75),
    .X(_1984_));
 sky130_fd_sc_hd__a211o_1 _5238_ (.A1(net76),
    .A2(_1965_),
    .B1(_1967_),
    .C1(net119),
    .X(_1985_));
 sky130_fd_sc_hd__and3_1 _5239_ (.A(net220),
    .B(\as2650.stack[3][2] ),
    .C(net172),
    .X(_1986_));
 sky130_fd_sc_hd__o22a_1 _5240_ (.A1(\as2650.stack[1][2] ),
    .A2(net166),
    .B1(net155),
    .B2(\as2650.stack[0][2] ),
    .X(_1987_));
 sky130_fd_sc_hd__o221a_2 _5241_ (.A1(\as2650.stack[2][2] ),
    .A2(net169),
    .B1(_1986_),
    .B2(net158),
    .C1(_1987_),
    .X(_1988_));
 sky130_fd_sc_hd__o22a_1 _5242_ (.A1(\as2650.stack[7][2] ),
    .A2(net171),
    .B1(net157),
    .B2(\as2650.stack[4][2] ),
    .X(_1989_));
 sky130_fd_sc_hd__o22a_1 _5243_ (.A1(\as2650.stack[5][2] ),
    .A2(net168),
    .B1(net170),
    .B2(\as2650.stack[6][2] ),
    .X(_1990_));
 sky130_fd_sc_hd__a31o_4 _5244_ (.A1(net107),
    .A2(_1989_),
    .A3(_1990_),
    .B1(_1988_),
    .X(_1991_));
 sky130_fd_sc_hd__o221a_1 _5245_ (.A1(net60),
    .A2(_1965_),
    .B1(_1991_),
    .B2(net63),
    .C1(net59),
    .X(_1992_));
 sky130_fd_sc_hd__and3_1 _5246_ (.A(_1984_),
    .B(_1985_),
    .C(_1992_),
    .X(_1993_));
 sky130_fd_sc_hd__a211o_1 _5247_ (.A1(net57),
    .A2(_1965_),
    .B1(_1993_),
    .C1(_1930_),
    .X(_1994_));
 sky130_fd_sc_hd__o211a_1 _5248_ (.A1(net279),
    .A2(net46),
    .B1(_1994_),
    .C1(net313),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_2 _5249_ (.A0(net278),
    .A1(_1460_),
    .S(net309),
    .X(_1995_));
 sky130_fd_sc_hd__mux2_1 _5250_ (.A0(net338),
    .A1(\as2650.addr_buff[3] ),
    .S(net122),
    .X(_1996_));
 sky130_fd_sc_hd__and2_4 _5251_ (.A(net278),
    .B(_1963_),
    .X(_1997_));
 sky130_fd_sc_hd__nor2_1 _5252_ (.A(net278),
    .B(_1963_),
    .Y(_1998_));
 sky130_fd_sc_hd__nor2_1 _5253_ (.A(_1997_),
    .B(_1998_),
    .Y(_1999_));
 sky130_fd_sc_hd__or2_2 _5254_ (.A(_1997_),
    .B(_1998_),
    .X(_2000_));
 sky130_fd_sc_hd__o21a_1 _5255_ (.A1(_2612_),
    .A2(_1996_),
    .B1(net138),
    .X(_2001_));
 sky130_fd_sc_hd__o221a_1 _5256_ (.A1(_2627_),
    .A2(_1995_),
    .B1(_1999_),
    .B2(net83),
    .C1(_2001_),
    .X(_2002_));
 sky130_fd_sc_hd__and2_1 _5257_ (.A(net338),
    .B(_2871_),
    .X(_2003_));
 sky130_fd_sc_hd__nand2_1 _5258_ (.A(net338),
    .B(_2871_),
    .Y(_2004_));
 sky130_fd_sc_hd__nor2_1 _5259_ (.A(net338),
    .B(_2871_),
    .Y(_2005_));
 sky130_fd_sc_hd__a211o_2 _5260_ (.A1(_1975_),
    .A2(_1978_),
    .B1(_2003_),
    .C1(_2005_),
    .X(_2006_));
 sky130_fd_sc_hd__o211a_1 _5261_ (.A1(_2003_),
    .A2(_2005_),
    .B1(_1975_),
    .C1(_1978_),
    .X(_2007_));
 sky130_fd_sc_hd__nor2_1 _5262_ (.A(net125),
    .B(_2007_),
    .Y(_2008_));
 sky130_fd_sc_hd__a22o_1 _5263_ (.A1(net338),
    .A2(net125),
    .B1(_2006_),
    .B2(_2008_),
    .X(_2009_));
 sky130_fd_sc_hd__a2bb2o_1 _5264_ (.A1_N(_1783_),
    .A2_N(_2000_),
    .B1(_2009_),
    .B2(_1980_),
    .X(_2010_));
 sky130_fd_sc_hd__and3_2 _5265_ (.A(net278),
    .B(net280),
    .C(_1945_),
    .X(_2011_));
 sky130_fd_sc_hd__a21oi_1 _5266_ (.A1(net279),
    .A2(_1945_),
    .B1(net278),
    .Y(_2012_));
 sky130_fd_sc_hd__nor2_1 _5267_ (.A(_2011_),
    .B(_2012_),
    .Y(_2013_));
 sky130_fd_sc_hd__a221o_1 _5268_ (.A1(_1822_),
    .A2(_1999_),
    .B1(_2013_),
    .B2(_1947_),
    .C1(_2002_),
    .X(_2014_));
 sky130_fd_sc_hd__a21o_1 _5269_ (.A1(net133),
    .A2(_2014_),
    .B1(_2010_),
    .X(_2015_));
 sky130_fd_sc_hd__a221o_1 _5270_ (.A1(net50),
    .A2(_1995_),
    .B1(_1999_),
    .B2(_2689_),
    .C1(_2603_),
    .X(_2016_));
 sky130_fd_sc_hd__o21ai_2 _5271_ (.A1(net120),
    .A2(_2015_),
    .B1(_2016_),
    .Y(_2017_));
 sky130_fd_sc_hd__and3_1 _5272_ (.A(net220),
    .B(\as2650.stack[3][3] ),
    .C(net172),
    .X(_2018_));
 sky130_fd_sc_hd__o22a_1 _5273_ (.A1(\as2650.stack[1][3] ),
    .A2(net166),
    .B1(net155),
    .B2(\as2650.stack[0][3] ),
    .X(_2019_));
 sky130_fd_sc_hd__o221a_2 _5274_ (.A1(\as2650.stack[2][3] ),
    .A2(net170),
    .B1(_2018_),
    .B2(net158),
    .C1(_2019_),
    .X(_2020_));
 sky130_fd_sc_hd__mux4_2 _5275_ (.A0(\as2650.stack[7][3] ),
    .A1(\as2650.stack[4][3] ),
    .A2(\as2650.stack[5][3] ),
    .A3(\as2650.stack[6][3] ),
    .S0(net216),
    .S1(net218),
    .X(_2021_));
 sky130_fd_sc_hd__a21oi_4 _5276_ (.A1(net107),
    .A2(_2021_),
    .B1(_2020_),
    .Y(_2022_));
 sky130_fd_sc_hd__inv_2 _5277_ (.A(_2022_),
    .Y(_2023_));
 sky130_fd_sc_hd__o221a_1 _5278_ (.A1(net60),
    .A2(_2000_),
    .B1(_2022_),
    .B2(net63),
    .C1(_2017_),
    .X(_2024_));
 sky130_fd_sc_hd__nor2_1 _5279_ (.A(net58),
    .B(_2000_),
    .Y(_2025_));
 sky130_fd_sc_hd__o21ai_1 _5280_ (.A1(_1310_),
    .A2(_2024_),
    .B1(net45),
    .Y(_2026_));
 sky130_fd_sc_hd__o221a_1 _5281_ (.A1(\as2650.pc[3] ),
    .A2(net45),
    .B1(_2025_),
    .B2(_2026_),
    .C1(net315),
    .X(_0211_));
 sky130_fd_sc_hd__xnor2_4 _5282_ (.A(net275),
    .B(_1997_),
    .Y(_2027_));
 sky130_fd_sc_hd__mux2_1 _5283_ (.A0(_2533_),
    .A1(_1478_),
    .S(net309),
    .X(_2028_));
 sky130_fd_sc_hd__mux2_1 _5284_ (.A0(net337),
    .A1(\as2650.addr_buff[4] ),
    .S(net122),
    .X(_2029_));
 sky130_fd_sc_hd__o2bb2a_1 _5285_ (.A1_N(net117),
    .A2_N(_2029_),
    .B1(_2027_),
    .B2(net83),
    .X(_2030_));
 sky130_fd_sc_hd__o211a_1 _5286_ (.A1(_2627_),
    .A2(_2028_),
    .B1(_2030_),
    .C1(net133),
    .X(_2031_));
 sky130_fd_sc_hd__and2_1 _5287_ (.A(net337),
    .B(_2920_),
    .X(_2032_));
 sky130_fd_sc_hd__nor2_1 _5288_ (.A(net337),
    .B(_2920_),
    .Y(_2033_));
 sky130_fd_sc_hd__o211a_1 _5289_ (.A1(_2032_),
    .A2(_2033_),
    .B1(_2004_),
    .C1(_2006_),
    .X(_2034_));
 sky130_fd_sc_hd__a211oi_2 _5290_ (.A1(_2004_),
    .A2(_2006_),
    .B1(_2032_),
    .C1(_2033_),
    .Y(_2035_));
 sky130_fd_sc_hd__or3_2 _5291_ (.A(net125),
    .B(_2034_),
    .C(_2035_),
    .X(_2036_));
 sky130_fd_sc_hd__nand2_1 _5292_ (.A(net337),
    .B(net122),
    .Y(_2037_));
 sky130_fd_sc_hd__a31o_1 _5293_ (.A1(_1255_),
    .A2(_2036_),
    .A3(_2037_),
    .B1(_2031_),
    .X(_2038_));
 sky130_fd_sc_hd__a21o_1 _5294_ (.A1(net138),
    .A2(_2038_),
    .B1(net75),
    .X(_2039_));
 sky130_fd_sc_hd__xnor2_1 _5295_ (.A(net275),
    .B(_2011_),
    .Y(_2040_));
 sky130_fd_sc_hd__a31o_1 _5296_ (.A1(net133),
    .A2(_1947_),
    .A3(_2040_),
    .B1(_2039_),
    .X(_2041_));
 sky130_fd_sc_hd__a21o_1 _5297_ (.A1(net76),
    .A2(_2027_),
    .B1(net119),
    .X(_2042_));
 sky130_fd_sc_hd__a21o_1 _5298_ (.A1(net138),
    .A2(_2028_),
    .B1(_2042_),
    .X(_2043_));
 sky130_fd_sc_hd__a32o_1 _5299_ (.A1(net59),
    .A2(_2041_),
    .A3(_2043_),
    .B1(_1933_),
    .B2(_2027_),
    .X(_2044_));
 sky130_fd_sc_hd__mux4_2 _5300_ (.A0(\as2650.stack[7][4] ),
    .A1(\as2650.stack[4][4] ),
    .A2(\as2650.stack[5][4] ),
    .A3(\as2650.stack[6][4] ),
    .S0(net216),
    .S1(net218),
    .X(_2045_));
 sky130_fd_sc_hd__o22a_1 _5301_ (.A1(\as2650.stack[3][4] ),
    .A2(net171),
    .B1(net170),
    .B2(\as2650.stack[2][4] ),
    .X(_2046_));
 sky130_fd_sc_hd__o221a_2 _5302_ (.A1(\as2650.stack[1][4] ),
    .A2(net168),
    .B1(net157),
    .B2(\as2650.stack[0][4] ),
    .C1(_2801_),
    .X(_2047_));
 sky130_fd_sc_hd__a22oi_4 _5303_ (.A1(net107),
    .A2(_2045_),
    .B1(_2046_),
    .B2(_2047_),
    .Y(_2048_));
 sky130_fd_sc_hd__o21a_1 _5304_ (.A1(net63),
    .A2(_2048_),
    .B1(_2044_),
    .X(_2049_));
 sky130_fd_sc_hd__a21oi_1 _5305_ (.A1(net57),
    .A2(_2027_),
    .B1(_2049_),
    .Y(_2050_));
 sky130_fd_sc_hd__o21ai_1 _5306_ (.A1(net60),
    .A2(_2027_),
    .B1(net46),
    .Y(_2051_));
 sky130_fd_sc_hd__o221a_1 _5307_ (.A1(\as2650.pc[4] ),
    .A2(net46),
    .B1(_2050_),
    .B2(_2051_),
    .C1(net314),
    .X(_0212_));
 sky130_fd_sc_hd__and3_1 _5308_ (.A(net274),
    .B(net275),
    .C(_1997_),
    .X(_2052_));
 sky130_fd_sc_hd__a21oi_1 _5309_ (.A1(net275),
    .A2(_1997_),
    .B1(net274),
    .Y(_2053_));
 sky130_fd_sc_hd__nor2_1 _5310_ (.A(_2052_),
    .B(_2053_),
    .Y(_2054_));
 sky130_fd_sc_hd__or2_2 _5311_ (.A(_2052_),
    .B(_2053_),
    .X(_2055_));
 sky130_fd_sc_hd__and3_2 _5312_ (.A(net274),
    .B(net275),
    .C(_2011_),
    .X(_2056_));
 sky130_fd_sc_hd__a21oi_1 _5313_ (.A1(net275),
    .A2(_2011_),
    .B1(net274),
    .Y(_2057_));
 sky130_fd_sc_hd__nand2_1 _5314_ (.A(net334),
    .B(_0327_),
    .Y(_2058_));
 sky130_fd_sc_hd__or2_1 _5315_ (.A(net334),
    .B(_0327_),
    .X(_2059_));
 sky130_fd_sc_hd__nand2_1 _5316_ (.A(_2058_),
    .B(_2059_),
    .Y(_2060_));
 sky130_fd_sc_hd__nor2_1 _5317_ (.A(_2032_),
    .B(_2035_),
    .Y(_2061_));
 sky130_fd_sc_hd__xor2_1 _5318_ (.A(_2060_),
    .B(_2061_),
    .X(_2062_));
 sky130_fd_sc_hd__mux2_2 _5319_ (.A0(net334),
    .A1(_2062_),
    .S(net129),
    .X(_2063_));
 sky130_fd_sc_hd__mux2_2 _5320_ (.A0(net273),
    .A1(_1535_),
    .S(net309),
    .X(_2064_));
 sky130_fd_sc_hd__nor2_1 _5321_ (.A(_2627_),
    .B(_2064_),
    .Y(_2065_));
 sky130_fd_sc_hd__nand2_1 _5322_ (.A(\as2650.addr_buff[5] ),
    .B(net122),
    .Y(_2066_));
 sky130_fd_sc_hd__a32o_1 _5323_ (.A1(net117),
    .A2(_1532_),
    .A3(_2066_),
    .B1(_2055_),
    .B2(_1335_),
    .X(_2067_));
 sky130_fd_sc_hd__or3_1 _5324_ (.A(net77),
    .B(_2065_),
    .C(_2067_),
    .X(_2068_));
 sky130_fd_sc_hd__o31a_1 _5325_ (.A1(_1948_),
    .A2(_2056_),
    .A3(_2057_),
    .B1(_2068_),
    .X(_2069_));
 sky130_fd_sc_hd__a2bb2o_1 _5326_ (.A1_N(net135),
    .A2_N(_2069_),
    .B1(_2054_),
    .B2(_1933_),
    .X(_2070_));
 sky130_fd_sc_hd__a211o_1 _5327_ (.A1(_1980_),
    .A2(_2063_),
    .B1(_2070_),
    .C1(net120),
    .X(_2071_));
 sky130_fd_sc_hd__a221o_1 _5328_ (.A1(_2689_),
    .A2(_2054_),
    .B1(_2064_),
    .B2(net50),
    .C1(_2603_),
    .X(_2072_));
 sky130_fd_sc_hd__nand2_1 _5329_ (.A(_2071_),
    .B(_2072_),
    .Y(_2073_));
 sky130_fd_sc_hd__and3_1 _5330_ (.A(net220),
    .B(\as2650.stack[3][5] ),
    .C(net172),
    .X(_2074_));
 sky130_fd_sc_hd__o22a_1 _5331_ (.A1(\as2650.stack[1][5] ),
    .A2(net168),
    .B1(net157),
    .B2(\as2650.stack[0][5] ),
    .X(_2075_));
 sky130_fd_sc_hd__o221a_2 _5332_ (.A1(\as2650.stack[2][5] ),
    .A2(net170),
    .B1(_2074_),
    .B2(net158),
    .C1(_2075_),
    .X(_2076_));
 sky130_fd_sc_hd__mux4_2 _5333_ (.A0(\as2650.stack[7][5] ),
    .A1(\as2650.stack[4][5] ),
    .A2(\as2650.stack[5][5] ),
    .A3(\as2650.stack[6][5] ),
    .S0(net216),
    .S1(net218),
    .X(_2077_));
 sky130_fd_sc_hd__a21oi_4 _5334_ (.A1(net107),
    .A2(_2077_),
    .B1(_2076_),
    .Y(_2078_));
 sky130_fd_sc_hd__o221a_1 _5335_ (.A1(net60),
    .A2(_2055_),
    .B1(_2078_),
    .B2(net63),
    .C1(_2073_),
    .X(_2079_));
 sky130_fd_sc_hd__nor2_1 _5336_ (.A(net57),
    .B(_2079_),
    .Y(_2080_));
 sky130_fd_sc_hd__o21ai_1 _5337_ (.A1(net58),
    .A2(_2055_),
    .B1(net46),
    .Y(_2081_));
 sky130_fd_sc_hd__o221a_1 _5338_ (.A1(net274),
    .A2(net46),
    .B1(_2080_),
    .B2(_2081_),
    .C1(net315),
    .X(_0213_));
 sky130_fd_sc_hd__xor2_1 _5339_ (.A(\as2650.pc[6] ),
    .B(_2056_),
    .X(_2082_));
 sky130_fd_sc_hd__and2_2 _5340_ (.A(net272),
    .B(_2052_),
    .X(_2083_));
 sky130_fd_sc_hd__nor2_1 _5341_ (.A(net272),
    .B(_2052_),
    .Y(_2084_));
 sky130_fd_sc_hd__nor2_1 _5342_ (.A(_2083_),
    .B(_2084_),
    .Y(_2085_));
 sky130_fd_sc_hd__or2_1 _5343_ (.A(_2083_),
    .B(_2084_),
    .X(_2086_));
 sky130_fd_sc_hd__nand2_1 _5344_ (.A(net272),
    .B(net324),
    .Y(_2087_));
 sky130_fd_sc_hd__o21ai_2 _5345_ (.A1(net324),
    .A2(_1554_),
    .B1(_2087_),
    .Y(_2088_));
 sky130_fd_sc_hd__and2_1 _5346_ (.A(\as2650.addr_buff[6] ),
    .B(net125),
    .X(_2089_));
 sky130_fd_sc_hd__a211o_1 _5347_ (.A1(net330),
    .A2(net129),
    .B1(_2612_),
    .C1(_2089_),
    .X(_2090_));
 sky130_fd_sc_hd__o221a_1 _5348_ (.A1(net83),
    .A2(_2085_),
    .B1(_2088_),
    .B2(_2627_),
    .C1(_2090_),
    .X(_2091_));
 sky130_fd_sc_hd__a221o_1 _5349_ (.A1(_1822_),
    .A2(_2085_),
    .B1(_2091_),
    .B2(net143),
    .C1(net137),
    .X(_2092_));
 sky130_fd_sc_hd__a21oi_1 _5350_ (.A1(_1947_),
    .A2(_2082_),
    .B1(_2092_),
    .Y(_2093_));
 sky130_fd_sc_hd__nand2_1 _5351_ (.A(net330),
    .B(net125),
    .Y(_2094_));
 sky130_fd_sc_hd__and2_1 _5352_ (.A(net330),
    .B(_0382_),
    .X(_2095_));
 sky130_fd_sc_hd__nor2_1 _5353_ (.A(net330),
    .B(_0382_),
    .Y(_2096_));
 sky130_fd_sc_hd__o21a_1 _5354_ (.A1(_2060_),
    .A2(_2061_),
    .B1(_2058_),
    .X(_2097_));
 sky130_fd_sc_hd__nor3_1 _5355_ (.A(_2095_),
    .B(_2096_),
    .C(_2097_),
    .Y(_2098_));
 sky130_fd_sc_hd__o21a_1 _5356_ (.A1(_2095_),
    .A2(_2096_),
    .B1(_2097_),
    .X(_2099_));
 sky130_fd_sc_hd__o21ai_1 _5357_ (.A1(_1783_),
    .A2(_2085_),
    .B1(net229),
    .Y(_2100_));
 sky130_fd_sc_hd__nand2_1 _5358_ (.A(net143),
    .B(_2088_),
    .Y(_2101_));
 sky130_fd_sc_hd__o211a_1 _5359_ (.A1(net143),
    .A2(_2086_),
    .B1(_2101_),
    .C1(net120),
    .X(_2102_));
 sky130_fd_sc_hd__o311a_1 _5360_ (.A1(net125),
    .A2(_2098_),
    .A3(_2099_),
    .B1(_1980_),
    .C1(_2094_),
    .X(_2103_));
 sky130_fd_sc_hd__or4_1 _5361_ (.A(_2093_),
    .B(_2100_),
    .C(_2102_),
    .D(_2103_),
    .X(_2104_));
 sky130_fd_sc_hd__mux4_2 _5362_ (.A0(\as2650.stack[7][6] ),
    .A1(\as2650.stack[4][6] ),
    .A2(\as2650.stack[5][6] ),
    .A3(\as2650.stack[6][6] ),
    .S0(net216),
    .S1(net218),
    .X(_2105_));
 sky130_fd_sc_hd__o22a_1 _5363_ (.A1(\as2650.stack[3][6] ),
    .A2(net171),
    .B1(net170),
    .B2(\as2650.stack[2][6] ),
    .X(_2106_));
 sky130_fd_sc_hd__o221a_2 _5364_ (.A1(\as2650.stack[1][6] ),
    .A2(net168),
    .B1(net157),
    .B2(\as2650.stack[0][6] ),
    .C1(_2801_),
    .X(_2107_));
 sky130_fd_sc_hd__a22oi_4 _5365_ (.A1(net107),
    .A2(_2105_),
    .B1(_2106_),
    .B2(_2107_),
    .Y(_2108_));
 sky130_fd_sc_hd__o221a_1 _5366_ (.A1(net61),
    .A2(_2086_),
    .B1(_2108_),
    .B2(net63),
    .C1(_2104_),
    .X(_2109_));
 sky130_fd_sc_hd__mux2_1 _5367_ (.A0(_2086_),
    .A1(_2109_),
    .S(net58),
    .X(_2110_));
 sky130_fd_sc_hd__o21ai_1 _5368_ (.A1(\as2650.pc[6] ),
    .A2(net45),
    .B1(net321),
    .Y(_2111_));
 sky130_fd_sc_hd__a21oi_1 _5369_ (.A1(net45),
    .A2(_2110_),
    .B1(_2111_),
    .Y(_0214_));
 sky130_fd_sc_hd__and3_2 _5370_ (.A(net270),
    .B(net272),
    .C(_2056_),
    .X(_2112_));
 sky130_fd_sc_hd__a21oi_1 _5371_ (.A1(net272),
    .A2(_2056_),
    .B1(net270),
    .Y(_2113_));
 sky130_fd_sc_hd__xnor2_2 _5372_ (.A(net270),
    .B(_2083_),
    .Y(_2114_));
 sky130_fd_sc_hd__inv_2 _5373_ (.A(_2114_),
    .Y(_2115_));
 sky130_fd_sc_hd__and2_1 _5374_ (.A(net325),
    .B(_2721_),
    .X(_2116_));
 sky130_fd_sc_hd__nor2_1 _5375_ (.A(net325),
    .B(_2721_),
    .Y(_2117_));
 sky130_fd_sc_hd__nor2_1 _5376_ (.A(_2116_),
    .B(_2117_),
    .Y(_2118_));
 sky130_fd_sc_hd__nor2_1 _5377_ (.A(_2095_),
    .B(_2098_),
    .Y(_2119_));
 sky130_fd_sc_hd__xnor2_1 _5378_ (.A(_2118_),
    .B(_2119_),
    .Y(_2120_));
 sky130_fd_sc_hd__mux2_2 _5379_ (.A0(net269),
    .A1(_1608_),
    .S(net309),
    .X(_2121_));
 sky130_fd_sc_hd__mux2_1 _5380_ (.A0(net294),
    .A1(net324),
    .S(net128),
    .X(_2122_));
 sky130_fd_sc_hd__or2_1 _5381_ (.A(_2612_),
    .B(_2122_),
    .X(_2123_));
 sky130_fd_sc_hd__o211a_1 _5382_ (.A1(net83),
    .A2(_2115_),
    .B1(_2123_),
    .C1(net138),
    .X(_2124_));
 sky130_fd_sc_hd__o21ai_1 _5383_ (.A1(_2627_),
    .A2(_2121_),
    .B1(_2124_),
    .Y(_2125_));
 sky130_fd_sc_hd__o31a_1 _5384_ (.A1(_1948_),
    .A2(_2112_),
    .A3(_2113_),
    .B1(_2125_),
    .X(_2126_));
 sky130_fd_sc_hd__mux2_1 _5385_ (.A0(net325),
    .A1(_2120_),
    .S(net129),
    .X(_2127_));
 sky130_fd_sc_hd__a2bb2o_1 _5386_ (.A1_N(net135),
    .A2_N(_2126_),
    .B1(_2115_),
    .B2(_1933_),
    .X(_2128_));
 sky130_fd_sc_hd__a211o_1 _5387_ (.A1(_1980_),
    .A2(_2127_),
    .B1(_2128_),
    .C1(net120),
    .X(_2129_));
 sky130_fd_sc_hd__a221o_1 _5388_ (.A1(_2689_),
    .A2(_2115_),
    .B1(_2121_),
    .B2(_1333_),
    .C1(_2603_),
    .X(_2130_));
 sky130_fd_sc_hd__mux4_2 _5389_ (.A0(\as2650.stack[7][7] ),
    .A1(\as2650.stack[4][7] ),
    .A2(\as2650.stack[5][7] ),
    .A3(\as2650.stack[6][7] ),
    .S0(net216),
    .S1(net218),
    .X(_2131_));
 sky130_fd_sc_hd__o22a_1 _5390_ (.A1(\as2650.stack[3][7] ),
    .A2(net171),
    .B1(net170),
    .B2(\as2650.stack[2][7] ),
    .X(_2132_));
 sky130_fd_sc_hd__o221a_1 _5391_ (.A1(\as2650.stack[1][7] ),
    .A2(net168),
    .B1(net157),
    .B2(\as2650.stack[0][7] ),
    .C1(_2801_),
    .X(_2133_));
 sky130_fd_sc_hd__a22o_4 _5392_ (.A1(net107),
    .A2(_2131_),
    .B1(_2132_),
    .B2(_2133_),
    .X(_2134_));
 sky130_fd_sc_hd__a22o_1 _5393_ (.A1(_0725_),
    .A2(_2115_),
    .B1(_2134_),
    .B2(_0717_),
    .X(_2135_));
 sky130_fd_sc_hd__a21oi_1 _5394_ (.A1(_2129_),
    .A2(_2130_),
    .B1(_2135_),
    .Y(_2136_));
 sky130_fd_sc_hd__nor2_1 _5395_ (.A(net57),
    .B(_2136_),
    .Y(_2137_));
 sky130_fd_sc_hd__nor2_1 _5396_ (.A(net58),
    .B(_2114_),
    .Y(_2138_));
 sky130_fd_sc_hd__or2_1 _5397_ (.A(net270),
    .B(net45),
    .X(_2139_));
 sky130_fd_sc_hd__o311a_1 _5398_ (.A1(_1930_),
    .A2(_2137_),
    .A3(_2138_),
    .B1(_2139_),
    .C1(net315),
    .X(_0215_));
 sky130_fd_sc_hd__and2_1 _5399_ (.A(net268),
    .B(_2112_),
    .X(_2140_));
 sky130_fd_sc_hd__nor2_1 _5400_ (.A(net268),
    .B(_2112_),
    .Y(_2141_));
 sky130_fd_sc_hd__mux2_1 _5401_ (.A0(_2532_),
    .A1(_1645_),
    .S(net309),
    .X(_2142_));
 sky130_fd_sc_hd__nand2_1 _5402_ (.A(net296),
    .B(net128),
    .Y(_2143_));
 sky130_fd_sc_hd__a31o_1 _5403_ (.A1(net117),
    .A2(_1904_),
    .A3(_2143_),
    .B1(net77),
    .X(_2144_));
 sky130_fd_sc_hd__and3_1 _5404_ (.A(net268),
    .B(net270),
    .C(_2083_),
    .X(_2145_));
 sky130_fd_sc_hd__a21oi_1 _5405_ (.A1(net270),
    .A2(_2083_),
    .B1(net268),
    .Y(_2146_));
 sky130_fd_sc_hd__or2_4 _5406_ (.A(_2145_),
    .B(_2146_),
    .X(_2147_));
 sky130_fd_sc_hd__a221o_1 _5407_ (.A1(net116),
    .A2(_2142_),
    .B1(_2147_),
    .B2(_1335_),
    .C1(_2144_),
    .X(_2148_));
 sky130_fd_sc_hd__or2_1 _5408_ (.A(net148),
    .B(_2147_),
    .X(_2149_));
 sky130_fd_sc_hd__nor2_1 _5409_ (.A(net138),
    .B(_2147_),
    .Y(_2150_));
 sky130_fd_sc_hd__nand2_1 _5410_ (.A(_1821_),
    .B(_2150_),
    .Y(_2151_));
 sky130_fd_sc_hd__and3_1 _5411_ (.A(_2590_),
    .B(_2148_),
    .C(_2151_),
    .X(_2152_));
 sky130_fd_sc_hd__o31a_1 _5412_ (.A1(_1948_),
    .A2(_2140_),
    .A3(_2141_),
    .B1(_2152_),
    .X(_2153_));
 sky130_fd_sc_hd__o21ba_2 _5413_ (.A1(_2117_),
    .A2(_2119_),
    .B1_N(_2116_),
    .X(_2154_));
 sky130_fd_sc_hd__nor2_2 _5414_ (.A(net125),
    .B(_2154_),
    .Y(_2155_));
 sky130_fd_sc_hd__nor2_1 _5415_ (.A(net296),
    .B(_2155_),
    .Y(_2156_));
 sky130_fd_sc_hd__and2_1 _5416_ (.A(net296),
    .B(_2155_),
    .X(_2157_));
 sky130_fd_sc_hd__o311a_1 _5417_ (.A1(net149),
    .A2(_2156_),
    .A3(_2157_),
    .B1(net135),
    .C1(_2149_),
    .X(_2158_));
 sky130_fd_sc_hd__nor2_1 _5418_ (.A(net77),
    .B(_2142_),
    .Y(_2159_));
 sky130_fd_sc_hd__o31a_1 _5419_ (.A1(net119),
    .A2(_2150_),
    .A3(_2159_),
    .B1(net229),
    .X(_2160_));
 sky130_fd_sc_hd__or3b_2 _5420_ (.A(_2153_),
    .B(_2158_),
    .C_N(_2160_),
    .X(_2161_));
 sky130_fd_sc_hd__o2bb2a_1 _5421_ (.A1_N(_2804_),
    .A2_N(_0717_),
    .B1(net60),
    .B2(_2147_),
    .X(_2162_));
 sky130_fd_sc_hd__a21o_1 _5422_ (.A1(_2161_),
    .A2(_2162_),
    .B1(net57),
    .X(_2163_));
 sky130_fd_sc_hd__o211ai_1 _5423_ (.A1(net59),
    .A2(_2147_),
    .B1(_2163_),
    .C1(net44),
    .Y(_2164_));
 sky130_fd_sc_hd__o211a_1 _5424_ (.A1(\as2650.pc[8] ),
    .A2(net44),
    .B1(_2164_),
    .C1(net315),
    .X(_0216_));
 sky130_fd_sc_hd__nand2_1 _5425_ (.A(net295),
    .B(_2157_),
    .Y(_2165_));
 sky130_fd_sc_hd__o21a_1 _5426_ (.A1(net295),
    .A2(_2157_),
    .B1(net148),
    .X(_2166_));
 sky130_fd_sc_hd__and2_4 _5427_ (.A(net267),
    .B(_2145_),
    .X(_2167_));
 sky130_fd_sc_hd__nor2_1 _5428_ (.A(net267),
    .B(_2145_),
    .Y(_2168_));
 sky130_fd_sc_hd__or2_4 _5429_ (.A(_2167_),
    .B(_2168_),
    .X(_2169_));
 sky130_fd_sc_hd__a2bb2o_1 _5430_ (.A1_N(net148),
    .A2_N(_2169_),
    .B1(_2166_),
    .B2(_2165_),
    .X(_2170_));
 sky130_fd_sc_hd__mux2_1 _5431_ (.A0(net267),
    .A1(_1670_),
    .S(net310),
    .X(_2171_));
 sky130_fd_sc_hd__nor2_1 _5432_ (.A(net139),
    .B(_2169_),
    .Y(_2172_));
 sky130_fd_sc_hd__a211o_1 _5433_ (.A1(net139),
    .A2(_2171_),
    .B1(_2172_),
    .C1(_2602_),
    .X(_2173_));
 sky130_fd_sc_hd__and3_2 _5434_ (.A(net267),
    .B(\as2650.pc[8] ),
    .C(_2112_),
    .X(_2174_));
 sky130_fd_sc_hd__nor2_1 _5435_ (.A(\as2650.pc[9] ),
    .B(_2140_),
    .Y(_2175_));
 sky130_fd_sc_hd__mux2_1 _5436_ (.A0(net346),
    .A1(\as2650.addr_buff[1] ),
    .S(net130),
    .X(_2176_));
 sky130_fd_sc_hd__a2bb2o_1 _5437_ (.A1_N(net83),
    .A2_N(_2169_),
    .B1(_2176_),
    .B2(net117),
    .X(_2177_));
 sky130_fd_sc_hd__a21oi_1 _5438_ (.A1(_2626_),
    .A2(_2171_),
    .B1(_2177_),
    .Y(_2178_));
 sky130_fd_sc_hd__o21ba_1 _5439_ (.A1(_2174_),
    .A2(_2175_),
    .B1_N(_1821_),
    .X(_2179_));
 sky130_fd_sc_hd__a211o_1 _5440_ (.A1(_1821_),
    .A2(_2169_),
    .B1(_2179_),
    .C1(net139),
    .X(_2180_));
 sky130_fd_sc_hd__o21ai_1 _5441_ (.A1(net77),
    .A2(_2178_),
    .B1(_2180_),
    .Y(_2181_));
 sky130_fd_sc_hd__o211a_1 _5442_ (.A1(net133),
    .A2(_2170_),
    .B1(_2173_),
    .C1(net229),
    .X(_2182_));
 sky130_fd_sc_hd__o21ai_1 _5443_ (.A1(net137),
    .A2(_2181_),
    .B1(_2182_),
    .Y(_2183_));
 sky130_fd_sc_hd__o2bb2a_1 _5444_ (.A1_N(_2818_),
    .A2_N(_0717_),
    .B1(net61),
    .B2(_2169_),
    .X(_2184_));
 sky130_fd_sc_hd__a21oi_1 _5445_ (.A1(_2183_),
    .A2(_2184_),
    .B1(net57),
    .Y(_2185_));
 sky130_fd_sc_hd__o21ai_1 _5446_ (.A1(net59),
    .A2(_2169_),
    .B1(net44),
    .Y(_2186_));
 sky130_fd_sc_hd__o221a_1 _5447_ (.A1(\as2650.pc[9] ),
    .A2(net44),
    .B1(_2185_),
    .B2(_2186_),
    .C1(net319),
    .X(_0217_));
 sky130_fd_sc_hd__xor2_1 _5448_ (.A(\as2650.addr_buff[2] ),
    .B(_2165_),
    .X(_2187_));
 sky130_fd_sc_hd__mux2_2 _5449_ (.A0(_2531_),
    .A1(_1704_),
    .S(net310),
    .X(_2188_));
 sky130_fd_sc_hd__xnor2_4 _5450_ (.A(net266),
    .B(_2167_),
    .Y(_2189_));
 sky130_fd_sc_hd__mux2_1 _5451_ (.A0(net341),
    .A1(\as2650.addr_buff[2] ),
    .S(net127),
    .X(_2190_));
 sky130_fd_sc_hd__nand2_1 _5452_ (.A(net117),
    .B(_2190_),
    .Y(_2191_));
 sky130_fd_sc_hd__o221a_1 _5453_ (.A1(_2627_),
    .A2(_2188_),
    .B1(_2189_),
    .B2(net84),
    .C1(_2191_),
    .X(_2192_));
 sky130_fd_sc_hd__a22o_1 _5454_ (.A1(_1255_),
    .A2(_2187_),
    .B1(_2192_),
    .B2(net133),
    .X(_2193_));
 sky130_fd_sc_hd__xnor2_1 _5455_ (.A(net266),
    .B(_2174_),
    .Y(_2194_));
 sky130_fd_sc_hd__a31o_1 _5456_ (.A1(net134),
    .A2(_1947_),
    .A3(_2194_),
    .B1(net120),
    .X(_2195_));
 sky130_fd_sc_hd__a22o_1 _5457_ (.A1(_1933_),
    .A2(_2189_),
    .B1(_2193_),
    .B2(net139),
    .X(_2196_));
 sky130_fd_sc_hd__a221o_1 _5458_ (.A1(_1333_),
    .A2(_2188_),
    .B1(_2189_),
    .B2(_2689_),
    .C1(_2603_),
    .X(_2197_));
 sky130_fd_sc_hd__o21ai_1 _5459_ (.A1(_2195_),
    .A2(_2196_),
    .B1(_2197_),
    .Y(_2198_));
 sky130_fd_sc_hd__o2bb2a_1 _5460_ (.A1_N(_0725_),
    .A2_N(_2189_),
    .B1(_2865_),
    .B2(net63),
    .X(_2199_));
 sky130_fd_sc_hd__o21ai_1 _5461_ (.A1(net58),
    .A2(_2189_),
    .B1(net46),
    .Y(_2200_));
 sky130_fd_sc_hd__a31o_1 _5462_ (.A1(net58),
    .A2(_2198_),
    .A3(_2199_),
    .B1(_2200_),
    .X(_2201_));
 sky130_fd_sc_hd__o211a_1 _5463_ (.A1(net266),
    .A2(net46),
    .B1(_2201_),
    .C1(net319),
    .X(_0218_));
 sky130_fd_sc_hd__a21o_1 _5464_ (.A1(_1681_),
    .A2(_2155_),
    .B1(\as2650.addr_buff[3] ),
    .X(_2202_));
 sky130_fd_sc_hd__o31ai_1 _5465_ (.A1(net122),
    .A2(_1736_),
    .A3(_2154_),
    .B1(_2202_),
    .Y(_2203_));
 sky130_fd_sc_hd__mux2_2 _5466_ (.A0(net265),
    .A1(_1729_),
    .S(net310),
    .X(_2204_));
 sky130_fd_sc_hd__nand2_1 _5467_ (.A(net116),
    .B(_2204_),
    .Y(_2205_));
 sky130_fd_sc_hd__and3_1 _5468_ (.A(net265),
    .B(\as2650.pc[10] ),
    .C(_2167_),
    .X(_2206_));
 sky130_fd_sc_hd__a21oi_1 _5469_ (.A1(\as2650.pc[10] ),
    .A2(_2167_),
    .B1(\as2650.pc[11] ),
    .Y(_2207_));
 sky130_fd_sc_hd__or2_4 _5470_ (.A(_2206_),
    .B(_2207_),
    .X(_2208_));
 sky130_fd_sc_hd__mux2_1 _5471_ (.A0(net340),
    .A1(\as2650.addr_buff[3] ),
    .S(net129),
    .X(_2209_));
 sky130_fd_sc_hd__o2bb2a_1 _5472_ (.A1_N(net117),
    .A2_N(_2209_),
    .B1(_2208_),
    .B2(net83),
    .X(_2210_));
 sky130_fd_sc_hd__a32o_1 _5473_ (.A1(net133),
    .A2(_2205_),
    .A3(_2210_),
    .B1(_1255_),
    .B2(_2203_),
    .X(_2211_));
 sky130_fd_sc_hd__and3_2 _5474_ (.A(\as2650.pc[11] ),
    .B(\as2650.pc[10] ),
    .C(_2174_),
    .X(_2212_));
 sky130_fd_sc_hd__a21oi_1 _5475_ (.A1(\as2650.pc[10] ),
    .A2(_2174_),
    .B1(net265),
    .Y(_2213_));
 sky130_fd_sc_hd__o211a_1 _5476_ (.A1(_2212_),
    .A2(_2213_),
    .B1(net133),
    .C1(_1947_),
    .X(_2214_));
 sky130_fd_sc_hd__a211o_1 _5477_ (.A1(_1933_),
    .A2(_2208_),
    .B1(_2214_),
    .C1(net75),
    .X(_2215_));
 sky130_fd_sc_hd__a21o_1 _5478_ (.A1(net143),
    .A2(_2211_),
    .B1(_2215_),
    .X(_2216_));
 sky130_fd_sc_hd__o22a_1 _5479_ (.A1(_2910_),
    .A2(net63),
    .B1(net60),
    .B2(_2208_),
    .X(_2217_));
 sky130_fd_sc_hd__nor2_1 _5480_ (.A(net77),
    .B(_2204_),
    .Y(_2218_));
 sky130_fd_sc_hd__a211o_1 _5481_ (.A1(net78),
    .A2(_2208_),
    .B1(_2218_),
    .C1(net119),
    .X(_2219_));
 sky130_fd_sc_hd__a31o_1 _5482_ (.A1(_2216_),
    .A2(_2217_),
    .A3(_2219_),
    .B1(net57),
    .X(_2220_));
 sky130_fd_sc_hd__o211ai_1 _5483_ (.A1(net58),
    .A2(_2208_),
    .B1(_2220_),
    .C1(net44),
    .Y(_2221_));
 sky130_fd_sc_hd__o211a_1 _5484_ (.A1(net265),
    .A2(net44),
    .B1(_2221_),
    .C1(net319),
    .X(_0219_));
 sky130_fd_sc_hd__and2_2 _5485_ (.A(net264),
    .B(_2206_),
    .X(_2222_));
 sky130_fd_sc_hd__nor2_1 _5486_ (.A(net264),
    .B(_2206_),
    .Y(_2223_));
 sky130_fd_sc_hd__or2_4 _5487_ (.A(_2222_),
    .B(_2223_),
    .X(_2224_));
 sky130_fd_sc_hd__inv_2 _5488_ (.A(_2224_),
    .Y(_2225_));
 sky130_fd_sc_hd__a31o_1 _5489_ (.A1(\as2650.addr_buff[3] ),
    .A2(_1681_),
    .A3(_2155_),
    .B1(\as2650.addr_buff[4] ),
    .X(_2226_));
 sky130_fd_sc_hd__nand4_2 _5490_ (.A(\as2650.addr_buff[3] ),
    .B(\as2650.addr_buff[4] ),
    .C(_1681_),
    .D(_2155_),
    .Y(_2227_));
 sky130_fd_sc_hd__a21bo_1 _5491_ (.A1(_2226_),
    .A2(_2227_),
    .B1_N(_1255_),
    .X(_2228_));
 sky130_fd_sc_hd__mux2_2 _5492_ (.A0(net264),
    .A1(_1754_),
    .S(net309),
    .X(_2229_));
 sky130_fd_sc_hd__a21bo_1 _5493_ (.A1(\as2650.addr_buff[4] ),
    .A2(net129),
    .B1_N(_2037_),
    .X(_2230_));
 sky130_fd_sc_hd__a221o_1 _5494_ (.A1(_1335_),
    .A2(_2225_),
    .B1(_2230_),
    .B2(net117),
    .C1(net135),
    .X(_2231_));
 sky130_fd_sc_hd__a21o_1 _5495_ (.A1(net116),
    .A2(_2229_),
    .B1(_2231_),
    .X(_2232_));
 sky130_fd_sc_hd__a21oi_1 _5496_ (.A1(_2228_),
    .A2(_2232_),
    .B1(net77),
    .Y(_2233_));
 sky130_fd_sc_hd__and2_1 _5497_ (.A(net264),
    .B(_2212_),
    .X(_2234_));
 sky130_fd_sc_hd__nor2_1 _5498_ (.A(\as2650.pc[12] ),
    .B(_2212_),
    .Y(_2235_));
 sky130_fd_sc_hd__o211a_1 _5499_ (.A1(_2234_),
    .A2(_2235_),
    .B1(net133),
    .C1(_1947_),
    .X(_2236_));
 sky130_fd_sc_hd__nor2_1 _5500_ (.A(net76),
    .B(_2229_),
    .Y(_2237_));
 sky130_fd_sc_hd__a211o_1 _5501_ (.A1(net76),
    .A2(_2224_),
    .B1(_2237_),
    .C1(net119),
    .X(_2238_));
 sky130_fd_sc_hd__o31a_1 _5502_ (.A1(net75),
    .A2(_2233_),
    .A3(_2236_),
    .B1(net59),
    .X(_2239_));
 sky130_fd_sc_hd__a22o_1 _5503_ (.A1(_1933_),
    .A2(_2224_),
    .B1(_2238_),
    .B2(_2239_),
    .X(_2240_));
 sky130_fd_sc_hd__o21a_1 _5504_ (.A1(_0317_),
    .A2(net63),
    .B1(_2240_),
    .X(_2241_));
 sky130_fd_sc_hd__a21oi_1 _5505_ (.A1(_1310_),
    .A2(_2224_),
    .B1(_2241_),
    .Y(_2242_));
 sky130_fd_sc_hd__o21ai_1 _5506_ (.A1(net60),
    .A2(_2224_),
    .B1(net44),
    .Y(_2243_));
 sky130_fd_sc_hd__o221a_1 _5507_ (.A1(net264),
    .A2(net44),
    .B1(_2242_),
    .B2(_2243_),
    .C1(net315),
    .X(_0220_));
 sky130_fd_sc_hd__nand2_4 _5508_ (.A(\as2650.pc[13] ),
    .B(_2222_),
    .Y(_2244_));
 sky130_fd_sc_hd__or2_1 _5509_ (.A(\as2650.pc[13] ),
    .B(_2222_),
    .X(_2245_));
 sky130_fd_sc_hd__nand2_2 _5510_ (.A(_2244_),
    .B(_2245_),
    .Y(_2246_));
 sky130_fd_sc_hd__or2_1 _5511_ (.A(_1335_),
    .B(_1822_),
    .X(_2247_));
 sky130_fd_sc_hd__a21o_1 _5512_ (.A1(net83),
    .A2(_1823_),
    .B1(_2246_),
    .X(_2248_));
 sky130_fd_sc_hd__xnor2_1 _5513_ (.A(\as2650.pc[13] ),
    .B(_2234_),
    .Y(_2249_));
 sky130_fd_sc_hd__a31o_1 _5514_ (.A1(\as2650.pc[13] ),
    .A2(net327),
    .A3(net116),
    .B1(net135),
    .X(_2250_));
 sky130_fd_sc_hd__a21oi_1 _5515_ (.A1(\as2650.addr_buff[5] ),
    .A2(net129),
    .B1(_2250_),
    .Y(_2251_));
 sky130_fd_sc_hd__o211a_1 _5516_ (.A1(_1948_),
    .A2(_2249_),
    .B1(_2251_),
    .C1(_2248_),
    .X(_2252_));
 sky130_fd_sc_hd__a31o_1 _5517_ (.A1(net149),
    .A2(net136),
    .A3(_2246_),
    .B1(net75),
    .X(_2253_));
 sky130_fd_sc_hd__a311o_1 _5518_ (.A1(_1980_),
    .A2(_2066_),
    .A3(_2227_),
    .B1(_2252_),
    .C1(_2253_),
    .X(_2254_));
 sky130_fd_sc_hd__o22a_1 _5519_ (.A1(_0370_),
    .A2(net63),
    .B1(net60),
    .B2(_2246_),
    .X(_2255_));
 sky130_fd_sc_hd__a21oi_1 _5520_ (.A1(\as2650.pc[13] ),
    .A2(net327),
    .B1(net78),
    .Y(_2256_));
 sky130_fd_sc_hd__a211o_1 _5521_ (.A1(net78),
    .A2(_2246_),
    .B1(_2256_),
    .C1(net119),
    .X(_2257_));
 sky130_fd_sc_hd__a31o_1 _5522_ (.A1(_2254_),
    .A2(_2255_),
    .A3(_2257_),
    .B1(net57),
    .X(_2258_));
 sky130_fd_sc_hd__o211ai_1 _5523_ (.A1(net58),
    .A2(_2246_),
    .B1(_2258_),
    .C1(net45),
    .Y(_2259_));
 sky130_fd_sc_hd__o211a_1 _5524_ (.A1(\as2650.pc[13] ),
    .A2(net45),
    .B1(_2259_),
    .C1(net315),
    .X(_0221_));
 sky130_fd_sc_hd__xnor2_4 _5525_ (.A(\as2650.pc[14] ),
    .B(_2244_),
    .Y(_2260_));
 sky130_fd_sc_hd__nand3_1 _5526_ (.A(\as2650.pc[14] ),
    .B(\as2650.pc[13] ),
    .C(_2234_),
    .Y(_2261_));
 sky130_fd_sc_hd__a31o_1 _5527_ (.A1(\as2650.pc[13] ),
    .A2(\as2650.pc[12] ),
    .A3(_2212_),
    .B1(\as2650.pc[14] ),
    .X(_2262_));
 sky130_fd_sc_hd__and3_1 _5528_ (.A(_1947_),
    .B(_2261_),
    .C(_2262_),
    .X(_2263_));
 sky130_fd_sc_hd__and3_1 _5529_ (.A(\as2650.pc[14] ),
    .B(net327),
    .C(net116),
    .X(_2264_));
 sky130_fd_sc_hd__a2111o_1 _5530_ (.A1(\as2650.addr_buff[6] ),
    .A2(net129),
    .B1(_2263_),
    .C1(_2264_),
    .D1(net137),
    .X(_2265_));
 sky130_fd_sc_hd__a21o_1 _5531_ (.A1(_2247_),
    .A2(_2260_),
    .B1(_2265_),
    .X(_2266_));
 sky130_fd_sc_hd__and3_1 _5532_ (.A(\as2650.pc[14] ),
    .B(net327),
    .C(net143),
    .X(_2267_));
 sky130_fd_sc_hd__a211o_1 _5533_ (.A1(net78),
    .A2(_2260_),
    .B1(_2267_),
    .C1(net119),
    .X(_2268_));
 sky130_fd_sc_hd__o221a_1 _5534_ (.A1(_1981_),
    .A2(_2089_),
    .B1(_2260_),
    .B2(_1783_),
    .C1(net229),
    .X(_2269_));
 sky130_fd_sc_hd__and3_1 _5535_ (.A(_2266_),
    .B(_2268_),
    .C(_2269_),
    .X(_2270_));
 sky130_fd_sc_hd__a221o_1 _5536_ (.A1(_0422_),
    .A2(_0717_),
    .B1(_0725_),
    .B2(_2260_),
    .C1(_2270_),
    .X(_2271_));
 sky130_fd_sc_hd__mux2_1 _5537_ (.A0(_2260_),
    .A1(_2271_),
    .S(net58),
    .X(_2272_));
 sky130_fd_sc_hd__or2_1 _5538_ (.A(\as2650.pc[14] ),
    .B(net45),
    .X(_2273_));
 sky130_fd_sc_hd__o211a_1 _5539_ (.A1(_1930_),
    .A2(_2272_),
    .B1(_2273_),
    .C1(net315),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _5540_ (.A0(_2736_),
    .A1(_2746_),
    .S(net72),
    .X(_2274_));
 sky130_fd_sc_hd__or2_1 _5541_ (.A(net131),
    .B(_2274_),
    .X(_2275_));
 sky130_fd_sc_hd__o211a_1 _5542_ (.A1(net126),
    .A2(_2771_),
    .B1(net53),
    .C1(_2275_),
    .X(_2276_));
 sky130_fd_sc_hd__a21oi_1 _5543_ (.A1(\as2650.psu[0] ),
    .A2(net64),
    .B1(_2780_),
    .Y(_2277_));
 sky130_fd_sc_hd__o21ai_1 _5544_ (.A1(_2526_),
    .A2(net64),
    .B1(_2277_),
    .Y(_2278_));
 sky130_fd_sc_hd__o211a_1 _5545_ (.A1(net192),
    .A2(_2775_),
    .B1(_0631_),
    .C1(_2278_),
    .X(_2279_));
 sky130_fd_sc_hd__o21a_1 _5546_ (.A1(net66),
    .A2(_1915_),
    .B1(_2279_),
    .X(_2280_));
 sky130_fd_sc_hd__a211o_1 _5547_ (.A1(_2727_),
    .A2(_0630_),
    .B1(_2280_),
    .C1(_2662_),
    .X(_2281_));
 sky130_fd_sc_hd__o21a_1 _5548_ (.A1(_2663_),
    .A2(net111),
    .B1(_2681_),
    .X(_2282_));
 sky130_fd_sc_hd__a22o_1 _5549_ (.A1(net350),
    .A2(net115),
    .B1(_2281_),
    .B2(_2282_),
    .X(_2283_));
 sky130_fd_sc_hd__and4bb_1 _5550_ (.A_N(_0723_),
    .B_N(_0797_),
    .C(_0802_),
    .D(_0774_),
    .X(_2284_));
 sky130_fd_sc_hd__o21ai_2 _5551_ (.A1(_2684_),
    .A2(_1369_),
    .B1(net202),
    .Y(_2285_));
 sky130_fd_sc_hd__o221a_1 _5552_ (.A1(net118),
    .A2(_2682_),
    .B1(net56),
    .B2(_0805_),
    .C1(_2285_),
    .X(_2286_));
 sky130_fd_sc_hd__nor2_1 _5553_ (.A(net177),
    .B(_2286_),
    .Y(_2287_));
 sky130_fd_sc_hd__a31o_1 _5554_ (.A1(net299),
    .A2(net80),
    .A3(net177),
    .B1(net194),
    .X(_2288_));
 sky130_fd_sc_hd__nor2_1 _5555_ (.A(net121),
    .B(_2288_),
    .Y(_2289_));
 sky130_fd_sc_hd__nand2_1 _5556_ (.A(_0692_),
    .B(_0798_),
    .Y(_2290_));
 sky130_fd_sc_hd__o32ai_4 _5557_ (.A1(_2685_),
    .A2(_2687_),
    .A3(_0799_),
    .B1(_2698_),
    .B2(_2696_),
    .Y(_2291_));
 sky130_fd_sc_hd__or4_1 _5558_ (.A(_2589_),
    .B(_0731_),
    .C(_0788_),
    .D(_0803_),
    .X(_2292_));
 sky130_fd_sc_hd__or3b_1 _5559_ (.A(_2292_),
    .B(_0695_),
    .C_N(_0792_),
    .X(_2293_));
 sky130_fd_sc_hd__o211a_1 _5560_ (.A1(net142),
    .A2(_2682_),
    .B1(_1260_),
    .C1(_1299_),
    .X(_2294_));
 sky130_fd_sc_hd__a21oi_1 _5561_ (.A1(_2596_),
    .A2(_2697_),
    .B1(_1362_),
    .Y(_2295_));
 sky130_fd_sc_hd__o211a_1 _5562_ (.A1(net224),
    .A2(_2295_),
    .B1(_2294_),
    .C1(_1317_),
    .X(_2296_));
 sky130_fd_sc_hd__or4b_1 _5563_ (.A(_2580_),
    .B(_2284_),
    .C(_2289_),
    .D_N(_2296_),
    .X(_2297_));
 sky130_fd_sc_hd__or4_2 _5564_ (.A(_0721_),
    .B(_2287_),
    .C(_2293_),
    .D(_2297_),
    .X(_2298_));
 sky130_fd_sc_hd__nor4_4 _5565_ (.A(_0785_),
    .B(_2290_),
    .C(_2291_),
    .D(_2298_),
    .Y(_2299_));
 sky130_fd_sc_hd__clkinv_2 _5566_ (.A(_2299_),
    .Y(_2300_));
 sky130_fd_sc_hd__a221o_1 _5567_ (.A1(net113),
    .A2(net62),
    .B1(_2283_),
    .B2(net153),
    .C1(_2300_),
    .X(_2301_));
 sky130_fd_sc_hd__a211o_1 _5568_ (.A1(net162),
    .A2(_2709_),
    .B1(_2276_),
    .C1(_2301_),
    .X(_2302_));
 sky130_fd_sc_hd__o211a_1 _5569_ (.A1(net262),
    .A2(_2299_),
    .B1(_2302_),
    .C1(net317),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _5570_ (.A0(_2834_),
    .A1(_2838_),
    .S(net72),
    .X(_2303_));
 sky130_fd_sc_hd__or2_1 _5571_ (.A(net131),
    .B(_2303_),
    .X(_2304_));
 sky130_fd_sc_hd__o211a_1 _5572_ (.A1(net126),
    .A2(_2856_),
    .B1(net53),
    .C1(_2304_),
    .X(_2305_));
 sky130_fd_sc_hd__mux2_1 _5573_ (.A0(\as2650.psl[1] ),
    .A1(net218),
    .S(net64),
    .X(_2306_));
 sky130_fd_sc_hd__o21a_1 _5574_ (.A1(_2632_),
    .A2(_2775_),
    .B1(net55),
    .X(_2307_));
 sky130_fd_sc_hd__o221a_2 _5575_ (.A1(net66),
    .A2(_1959_),
    .B1(_2306_),
    .B2(_2780_),
    .C1(_2307_),
    .X(_2308_));
 sky130_fd_sc_hd__mux2_1 _5576_ (.A0(net105),
    .A1(net114),
    .S(net297),
    .X(_2309_));
 sky130_fd_sc_hd__a21o_1 _5577_ (.A1(_0633_),
    .A2(_2309_),
    .B1(net115),
    .X(_2310_));
 sky130_fd_sc_hd__o221a_1 _5578_ (.A1(net346),
    .A2(_2681_),
    .B1(_2308_),
    .B2(_2310_),
    .C1(_0638_),
    .X(_2311_));
 sky130_fd_sc_hd__a221o_1 _5579_ (.A1(net162),
    .A2(_2822_),
    .B1(net62),
    .B2(net112),
    .C1(_2311_),
    .X(_2312_));
 sky130_fd_sc_hd__or3_1 _5580_ (.A(_2300_),
    .B(_2305_),
    .C(_2312_),
    .X(_2313_));
 sky130_fd_sc_hd__o211a_1 _5581_ (.A1(net258),
    .A2(_2299_),
    .B1(_2313_),
    .C1(net316),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _5582_ (.A0(_2882_),
    .A1(_2886_),
    .S(net72),
    .X(_2314_));
 sky130_fd_sc_hd__or2_1 _5583_ (.A(net132),
    .B(_2314_),
    .X(_2315_));
 sky130_fd_sc_hd__o211a_1 _5584_ (.A1(net126),
    .A2(_2903_),
    .B1(net53),
    .C1(_2315_),
    .X(_2316_));
 sky130_fd_sc_hd__mux2_1 _5585_ (.A0(\as2650.overflow ),
    .A1(net221),
    .S(net64),
    .X(_2317_));
 sky130_fd_sc_hd__o221a_1 _5586_ (.A1(_2634_),
    .A2(_2775_),
    .B1(net66),
    .B2(_1991_),
    .C1(net55),
    .X(_2318_));
 sky130_fd_sc_hd__o21a_2 _5587_ (.A1(_2780_),
    .A2(_2317_),
    .B1(_2318_),
    .X(_2319_));
 sky130_fd_sc_hd__mux2_1 _5588_ (.A0(net103),
    .A1(net111),
    .S(net297),
    .X(_2320_));
 sky130_fd_sc_hd__a211o_1 _5589_ (.A1(_0633_),
    .A2(_2320_),
    .B1(_2319_),
    .C1(net115),
    .X(_2321_));
 sky130_fd_sc_hd__o211a_1 _5590_ (.A1(net343),
    .A2(_2681_),
    .B1(net153),
    .C1(_2321_),
    .X(_2322_));
 sky130_fd_sc_hd__a221o_1 _5591_ (.A1(net162),
    .A2(_2870_),
    .B1(net62),
    .B2(net105),
    .C1(_2322_),
    .X(_2323_));
 sky130_fd_sc_hd__or2_1 _5592_ (.A(net253),
    .B(_2299_),
    .X(_2324_));
 sky130_fd_sc_hd__o311a_1 _5593_ (.A1(_2300_),
    .A2(_2316_),
    .A3(_2323_),
    .B1(_2324_),
    .C1(net320),
    .X(_0225_));
 sky130_fd_sc_hd__nor2_1 _5594_ (.A(net72),
    .B(_0284_),
    .Y(_2325_));
 sky130_fd_sc_hd__a211o_1 _5595_ (.A1(net73),
    .A2(_0288_),
    .B1(_2325_),
    .C1(net131),
    .X(_2326_));
 sky130_fd_sc_hd__o211a_1 _5596_ (.A1(net126),
    .A2(_0309_),
    .B1(net53),
    .C1(_2326_),
    .X(_2327_));
 sky130_fd_sc_hd__mux2_1 _5597_ (.A0(\as2650.psl[3] ),
    .A1(\as2650.psu[3] ),
    .S(net64),
    .X(_2328_));
 sky130_fd_sc_hd__o21a_1 _5598_ (.A1(_2636_),
    .A2(_2775_),
    .B1(net56),
    .X(_2329_));
 sky130_fd_sc_hd__o221a_2 _5599_ (.A1(net66),
    .A2(_2023_),
    .B1(_2328_),
    .B2(_2780_),
    .C1(_2329_),
    .X(_2330_));
 sky130_fd_sc_hd__mux2_1 _5600_ (.A0(net99),
    .A1(net105),
    .S(net297),
    .X(_2331_));
 sky130_fd_sc_hd__a211o_1 _5601_ (.A1(_0633_),
    .A2(_2331_),
    .B1(_2330_),
    .C1(_2680_),
    .X(_2332_));
 sky130_fd_sc_hd__o211a_1 _5602_ (.A1(net339),
    .A2(_2681_),
    .B1(net153),
    .C1(_2332_),
    .X(_2333_));
 sky130_fd_sc_hd__a211o_1 _5603_ (.A1(net102),
    .A2(_0722_),
    .B1(_2300_),
    .C1(_2333_),
    .X(_2334_));
 sky130_fd_sc_hd__a211o_1 _5604_ (.A1(net162),
    .A2(_2914_),
    .B1(_2327_),
    .C1(_2334_),
    .X(_2335_));
 sky130_fd_sc_hd__o211a_1 _5605_ (.A1(net246),
    .A2(_2299_),
    .B1(_2335_),
    .C1(net317),
    .X(_0226_));
 sky130_fd_sc_hd__nand2_1 _5606_ (.A(net131),
    .B(_0360_),
    .Y(_2336_));
 sky130_fd_sc_hd__nor2_1 _5607_ (.A(_2671_),
    .B(_0341_),
    .Y(_2337_));
 sky130_fd_sc_hd__a211o_1 _5608_ (.A1(_2671_),
    .A2(_0337_),
    .B1(_2337_),
    .C1(net132),
    .X(_2338_));
 sky130_fd_sc_hd__mux2_1 _5609_ (.A0(net213),
    .A1(\as2650.psu[4] ),
    .S(net64),
    .X(_2339_));
 sky130_fd_sc_hd__nand2_1 _5610_ (.A(net70),
    .B(_2048_),
    .Y(_2340_));
 sky130_fd_sc_hd__o211a_1 _5611_ (.A1(net70),
    .A2(_2339_),
    .B1(_2340_),
    .C1(_2775_),
    .X(_2341_));
 sky130_fd_sc_hd__mux2_1 _5612_ (.A0(net97),
    .A1(net103),
    .S(net298),
    .X(_2342_));
 sky130_fd_sc_hd__a211o_1 _5613_ (.A1(_2638_),
    .A2(_2774_),
    .B1(_0633_),
    .C1(_2341_),
    .X(_2343_));
 sky130_fd_sc_hd__o21ai_2 _5614_ (.A1(net55),
    .A2(_2342_),
    .B1(_2343_),
    .Y(_2344_));
 sky130_fd_sc_hd__a21o_1 _5615_ (.A1(_2553_),
    .A2(_2680_),
    .B1(net152),
    .X(_2345_));
 sky130_fd_sc_hd__a21oi_2 _5616_ (.A1(_2681_),
    .A2(_2344_),
    .B1(_2345_),
    .Y(_2346_));
 sky130_fd_sc_hd__a221o_1 _5617_ (.A1(net162),
    .A2(_0321_),
    .B1(_0722_),
    .B2(net98),
    .C1(_2346_),
    .X(_2347_));
 sky130_fd_sc_hd__a311o_1 _5618_ (.A1(net54),
    .A2(_2336_),
    .A3(_2338_),
    .B1(_2347_),
    .C1(_2300_),
    .X(_2348_));
 sky130_fd_sc_hd__o211a_1 _5619_ (.A1(net245),
    .A2(_2299_),
    .B1(_2348_),
    .C1(net317),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _5620_ (.A0(_0394_),
    .A1(_0396_),
    .S(net73),
    .X(_2349_));
 sky130_fd_sc_hd__or2_1 _5621_ (.A(net132),
    .B(_2349_),
    .X(_2350_));
 sky130_fd_sc_hd__o211a_1 _5622_ (.A1(net126),
    .A2(_0414_),
    .B1(net54),
    .C1(_2350_),
    .X(_2351_));
 sky130_fd_sc_hd__mux2_1 _5623_ (.A0(\as2650.psl[5] ),
    .A1(\as2650.psu[5] ),
    .S(net64),
    .X(_2352_));
 sky130_fd_sc_hd__nand2_1 _5624_ (.A(net70),
    .B(_2078_),
    .Y(_2353_));
 sky130_fd_sc_hd__o221a_1 _5625_ (.A1(net182),
    .A2(_2775_),
    .B1(_2780_),
    .B2(_2352_),
    .C1(_0631_),
    .X(_2354_));
 sky130_fd_sc_hd__a22o_1 _5626_ (.A1(net100),
    .A2(_0630_),
    .B1(_2353_),
    .B2(_2354_),
    .X(_2355_));
 sky130_fd_sc_hd__mux2_1 _5627_ (.A0(net94),
    .A1(_2355_),
    .S(_2663_),
    .X(_2356_));
 sky130_fd_sc_hd__nor2_1 _5628_ (.A(net333),
    .B(_2681_),
    .Y(_2357_));
 sky130_fd_sc_hd__o21ai_1 _5629_ (.A1(net115),
    .A2(_2356_),
    .B1(net153),
    .Y(_2358_));
 sky130_fd_sc_hd__o221a_1 _5630_ (.A1(net194),
    .A2(_0381_),
    .B1(_2357_),
    .B2(_2358_),
    .C1(_2299_),
    .X(_2359_));
 sky130_fd_sc_hd__o21ai_1 _5631_ (.A1(_0329_),
    .A2(_0723_),
    .B1(_2359_),
    .Y(_2360_));
 sky130_fd_sc_hd__o221a_1 _5632_ (.A1(net240),
    .A2(_2299_),
    .B1(_2351_),
    .B2(_2360_),
    .C1(net317),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _5633_ (.A0(_0436_),
    .A1(_0439_),
    .S(net72),
    .X(_2361_));
 sky130_fd_sc_hd__or2_1 _5634_ (.A(net131),
    .B(_2361_),
    .X(_2362_));
 sky130_fd_sc_hd__o211a_1 _5635_ (.A1(net126),
    .A2(_0458_),
    .B1(net54),
    .C1(_2362_),
    .X(_2363_));
 sky130_fd_sc_hd__mux2_1 _5636_ (.A0(\as2650.psl[6] ),
    .A1(net30),
    .S(net64),
    .X(_2364_));
 sky130_fd_sc_hd__nand2_1 _5637_ (.A(net70),
    .B(_2108_),
    .Y(_2365_));
 sky130_fd_sc_hd__o221a_1 _5638_ (.A1(net180),
    .A2(_2775_),
    .B1(_2780_),
    .B2(_2364_),
    .C1(_2365_),
    .X(_2366_));
 sky130_fd_sc_hd__nand2_1 _5639_ (.A(_0329_),
    .B(_0630_),
    .Y(_2367_));
 sky130_fd_sc_hd__o211a_1 _5640_ (.A1(_0630_),
    .A2(_2366_),
    .B1(_2367_),
    .C1(_2663_),
    .X(_2368_));
 sky130_fd_sc_hd__a211o_1 _5641_ (.A1(_2662_),
    .A2(net109),
    .B1(_2368_),
    .C1(_2680_),
    .X(_2369_));
 sky130_fd_sc_hd__o211a_1 _5642_ (.A1(net7),
    .A2(_2681_),
    .B1(net153),
    .C1(_2369_),
    .X(_2370_));
 sky130_fd_sc_hd__a211o_1 _5643_ (.A1(_2587_),
    .A2(_0426_),
    .B1(_2300_),
    .C1(_2370_),
    .X(_2371_));
 sky130_fd_sc_hd__a211o_1 _5644_ (.A1(net93),
    .A2(net62),
    .B1(_2363_),
    .C1(_2371_),
    .X(_2372_));
 sky130_fd_sc_hd__o211a_1 _5645_ (.A1(net238),
    .A2(_2299_),
    .B1(_2372_),
    .C1(net317),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _5646_ (.A0(_0474_),
    .A1(_0477_),
    .S(net72),
    .X(_2373_));
 sky130_fd_sc_hd__or2_1 _5647_ (.A(net132),
    .B(_2373_),
    .X(_2374_));
 sky130_fd_sc_hd__o211a_1 _5648_ (.A1(net126),
    .A2(_0494_),
    .B1(net54),
    .C1(_2374_),
    .X(_2375_));
 sky130_fd_sc_hd__mux2_1 _5649_ (.A0(\as2650.psl[7] ),
    .A1(\as2650.psu[7] ),
    .S(net64),
    .X(_2376_));
 sky130_fd_sc_hd__o221a_1 _5650_ (.A1(_2722_),
    .A2(_2775_),
    .B1(_2780_),
    .B2(_2376_),
    .C1(net56),
    .X(_2377_));
 sky130_fd_sc_hd__o21ai_2 _5651_ (.A1(net66),
    .A2(_2134_),
    .B1(_2377_),
    .Y(_2378_));
 sky130_fd_sc_hd__nand2_1 _5652_ (.A(_0853_),
    .B(_2378_),
    .Y(_2379_));
 sky130_fd_sc_hd__mux2_1 _5653_ (.A0(net326),
    .A1(_2379_),
    .S(_2681_),
    .X(_2380_));
 sky130_fd_sc_hd__a221o_1 _5654_ (.A1(_2587_),
    .A2(_0463_),
    .B1(net153),
    .B2(_2380_),
    .C1(_2300_),
    .X(_2381_));
 sky130_fd_sc_hd__a211o_1 _5655_ (.A1(net110),
    .A2(net62),
    .B1(_2375_),
    .C1(_2381_),
    .X(_2382_));
 sky130_fd_sc_hd__o211a_1 _5656_ (.A1(net235),
    .A2(_2299_),
    .B1(_2382_),
    .C1(net317),
    .X(_0230_));
 sky130_fd_sc_hd__or2_4 _5657_ (.A(_2529_),
    .B(net170),
    .X(_2383_));
 sky130_fd_sc_hd__nor2_8 _5658_ (.A(net49),
    .B(_2383_),
    .Y(_2384_));
 sky130_fd_sc_hd__nor2_8 _5659_ (.A(_2559_),
    .B(net47),
    .Y(_2385_));
 sky130_fd_sc_hd__mux2_1 _5660_ (.A0(\as2650.stack[6][0] ),
    .A1(net286),
    .S(_2385_),
    .X(_2386_));
 sky130_fd_sc_hd__mux2_1 _5661_ (.A0(_2386_),
    .A1(net259),
    .S(_2384_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _5662_ (.A0(\as2650.stack[6][1] ),
    .A1(net282),
    .S(_2385_),
    .X(_2387_));
 sky130_fd_sc_hd__mux2_1 _5663_ (.A0(_2387_),
    .A1(net254),
    .S(_2384_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _5664_ (.A0(\as2650.stack[6][2] ),
    .A1(net280),
    .S(_2385_),
    .X(_2388_));
 sky130_fd_sc_hd__mux2_1 _5665_ (.A0(_2388_),
    .A1(net250),
    .S(_2384_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _5666_ (.A0(\as2650.stack[6][3] ),
    .A1(net277),
    .S(_2385_),
    .X(_2389_));
 sky130_fd_sc_hd__mux2_1 _5667_ (.A0(_2389_),
    .A1(net246),
    .S(_2384_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _5668_ (.A0(\as2650.stack[6][4] ),
    .A1(net276),
    .S(_2385_),
    .X(_2390_));
 sky130_fd_sc_hd__mux2_1 _5669_ (.A0(_2390_),
    .A1(net243),
    .S(_2384_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _5670_ (.A0(\as2650.stack[6][5] ),
    .A1(net273),
    .S(_2385_),
    .X(_2391_));
 sky130_fd_sc_hd__mux2_1 _5671_ (.A0(_2391_),
    .A1(net240),
    .S(_2384_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _5672_ (.A0(\as2650.stack[6][6] ),
    .A1(net271),
    .S(_2385_),
    .X(_2392_));
 sky130_fd_sc_hd__mux2_1 _5673_ (.A0(_2392_),
    .A1(net237),
    .S(_2384_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _5674_ (.A0(\as2650.stack[6][7] ),
    .A1(net269),
    .S(_2385_),
    .X(_2393_));
 sky130_fd_sc_hd__mux2_1 _5675_ (.A0(_2393_),
    .A1(net232),
    .S(_2384_),
    .X(_0238_));
 sky130_fd_sc_hd__nor2_8 _5676_ (.A(net47),
    .B(_2383_),
    .Y(_2394_));
 sky130_fd_sc_hd__mux2_1 _5677_ (.A0(\as2650.stack[7][0] ),
    .A1(net286),
    .S(_2394_),
    .X(_2395_));
 sky130_fd_sc_hd__mux2_1 _5678_ (.A0(net259),
    .A1(_2395_),
    .S(_0869_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _5679_ (.A0(\as2650.stack[7][1] ),
    .A1(net282),
    .S(_2394_),
    .X(_2396_));
 sky130_fd_sc_hd__mux2_1 _5680_ (.A0(net254),
    .A1(_2396_),
    .S(_0869_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _5681_ (.A0(\as2650.stack[7][2] ),
    .A1(net280),
    .S(_2394_),
    .X(_2397_));
 sky130_fd_sc_hd__mux2_1 _5682_ (.A0(net250),
    .A1(_2397_),
    .S(_0869_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _5683_ (.A0(\as2650.stack[7][3] ),
    .A1(net277),
    .S(_2394_),
    .X(_2398_));
 sky130_fd_sc_hd__mux2_1 _5684_ (.A0(net246),
    .A1(_2398_),
    .S(_0869_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _5685_ (.A0(\as2650.stack[7][4] ),
    .A1(net276),
    .S(_2394_),
    .X(_2399_));
 sky130_fd_sc_hd__mux2_1 _5686_ (.A0(net243),
    .A1(_2399_),
    .S(_0869_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _5687_ (.A0(\as2650.stack[7][5] ),
    .A1(net273),
    .S(_2394_),
    .X(_2400_));
 sky130_fd_sc_hd__mux2_1 _5688_ (.A0(net240),
    .A1(_2400_),
    .S(_0869_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _5689_ (.A0(\as2650.stack[7][6] ),
    .A1(net271),
    .S(_2394_),
    .X(_2401_));
 sky130_fd_sc_hd__mux2_1 _5690_ (.A0(net237),
    .A1(_2401_),
    .S(_0869_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _5691_ (.A0(\as2650.stack[7][7] ),
    .A1(net269),
    .S(_2394_),
    .X(_2402_));
 sky130_fd_sc_hd__mux2_1 _5692_ (.A0(net232),
    .A1(_2402_),
    .S(_0869_),
    .X(_0246_));
 sky130_fd_sc_hd__a21o_4 _5693_ (.A1(net48),
    .A2(_2618_),
    .B1(_2383_),
    .X(_2403_));
 sky130_fd_sc_hd__mux2_1 _5694_ (.A0(_2625_),
    .A1(\as2650.stack[7][8] ),
    .S(_2403_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _5695_ (.A0(_2633_),
    .A1(\as2650.stack[7][9] ),
    .S(_2403_),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _5696_ (.A0(_2635_),
    .A1(\as2650.stack[7][10] ),
    .S(_2403_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _5697_ (.A0(_2637_),
    .A1(\as2650.stack[7][11] ),
    .S(_2403_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _5698_ (.A0(_2639_),
    .A1(\as2650.stack[7][12] ),
    .S(_2403_),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _5699_ (.A0(_2641_),
    .A1(\as2650.stack[7][13] ),
    .S(_2403_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _5700_ (.A0(_2643_),
    .A1(\as2650.stack[7][14] ),
    .S(_2403_),
    .X(_0253_));
 sky130_fd_sc_hd__a21o_4 _5701_ (.A1(_2646_),
    .A2(_0871_),
    .B1(net348),
    .X(_2404_));
 sky130_fd_sc_hd__nor2_8 _5702_ (.A(net307),
    .B(_2785_),
    .Y(_2405_));
 sky130_fd_sc_hd__nor2_8 _5703_ (.A(_2404_),
    .B(_2405_),
    .Y(_2406_));
 sky130_fd_sc_hd__o21a_2 _5704_ (.A1(_2404_),
    .A2(_2405_),
    .B1(_2809_),
    .X(_2407_));
 sky130_fd_sc_hd__or3_4 _5705_ (.A(_2647_),
    .B(_2807_),
    .C(_2406_),
    .X(_2408_));
 sky130_fd_sc_hd__a32o_1 _5706_ (.A1(net260),
    .A2(net192),
    .A3(_2407_),
    .B1(_2405_),
    .B2(_2772_),
    .X(_2409_));
 sky130_fd_sc_hd__a21o_1 _5707_ (.A1(\as2650.r123[1][0] ),
    .A2(_2406_),
    .B1(_2409_),
    .X(_0254_));
 sky130_fd_sc_hd__a22oi_1 _5708_ (.A1(_2857_),
    .A2(_2405_),
    .B1(_2406_),
    .B2(\as2650.r123[1][1] ),
    .Y(_2410_));
 sky130_fd_sc_hd__o21ai_1 _5709_ (.A1(_0880_),
    .A2(net41),
    .B1(_2410_),
    .Y(_0255_));
 sky130_fd_sc_hd__a22oi_1 _5710_ (.A1(_2904_),
    .A2(_2405_),
    .B1(_2406_),
    .B2(\as2650.r123[1][2] ),
    .Y(_2411_));
 sky130_fd_sc_hd__o21ai_1 _5711_ (.A1(_0890_),
    .A2(net41),
    .B1(_2411_),
    .Y(_0256_));
 sky130_fd_sc_hd__nor2_1 _5712_ (.A(_0907_),
    .B(net41),
    .Y(_2412_));
 sky130_fd_sc_hd__a221o_1 _5713_ (.A1(_0310_),
    .A2(_2405_),
    .B1(_2406_),
    .B2(\as2650.r123[1][3] ),
    .C1(_2412_),
    .X(_0257_));
 sky130_fd_sc_hd__and2_1 _5714_ (.A(_0931_),
    .B(_2407_),
    .X(_2413_));
 sky130_fd_sc_hd__a221o_1 _5715_ (.A1(_0362_),
    .A2(_2405_),
    .B1(_2406_),
    .B2(\as2650.r123[1][4] ),
    .C1(_2413_),
    .X(_0258_));
 sky130_fd_sc_hd__nor2_1 _5716_ (.A(_0959_),
    .B(net41),
    .Y(_2414_));
 sky130_fd_sc_hd__a221o_1 _5717_ (.A1(_0415_),
    .A2(_2405_),
    .B1(_2406_),
    .B2(\as2650.r123[1][5] ),
    .C1(_2414_),
    .X(_0259_));
 sky130_fd_sc_hd__nor2_1 _5718_ (.A(_0993_),
    .B(_2408_),
    .Y(_2415_));
 sky130_fd_sc_hd__a221o_1 _5719_ (.A1(_0459_),
    .A2(_2405_),
    .B1(_2406_),
    .B2(\as2650.r123[1][6] ),
    .C1(_2415_),
    .X(_0260_));
 sky130_fd_sc_hd__nor2_1 _5720_ (.A(_1034_),
    .B(net41),
    .Y(_2416_));
 sky130_fd_sc_hd__a221o_1 _5721_ (.A1(_0495_),
    .A2(_2405_),
    .B1(_2406_),
    .B2(\as2650.r123[1][7] ),
    .C1(_2416_),
    .X(_0261_));
 sky130_fd_sc_hd__nor2_1 _5722_ (.A(_1077_),
    .B(_2408_),
    .Y(_2417_));
 sky130_fd_sc_hd__nor2_8 _5723_ (.A(_2584_),
    .B(_2785_),
    .Y(_2418_));
 sky130_fd_sc_hd__nor2_8 _5724_ (.A(_2404_),
    .B(_2418_),
    .Y(_2419_));
 sky130_fd_sc_hd__a221o_1 _5725_ (.A1(_2772_),
    .A2(_2418_),
    .B1(_2419_),
    .B2(\as2650.r123[2][0] ),
    .C1(_2417_),
    .X(_0262_));
 sky130_fd_sc_hd__nor2_1 _5726_ (.A(_1112_),
    .B(net41),
    .Y(_2420_));
 sky130_fd_sc_hd__a221o_1 _5727_ (.A1(_2857_),
    .A2(_2418_),
    .B1(_2419_),
    .B2(\as2650.r123[2][1] ),
    .C1(_2420_),
    .X(_0263_));
 sky130_fd_sc_hd__nor2_1 _5728_ (.A(_1144_),
    .B(net41),
    .Y(_2421_));
 sky130_fd_sc_hd__a221o_1 _5729_ (.A1(_2904_),
    .A2(_2418_),
    .B1(_2419_),
    .B2(\as2650.r123[2][2] ),
    .C1(_2421_),
    .X(_0264_));
 sky130_fd_sc_hd__nor2_1 _5730_ (.A(_1173_),
    .B(net41),
    .Y(_2422_));
 sky130_fd_sc_hd__a221o_1 _5731_ (.A1(_0310_),
    .A2(_2418_),
    .B1(_2419_),
    .B2(\as2650.r123[2][3] ),
    .C1(_2422_),
    .X(_0265_));
 sky130_fd_sc_hd__a2bb2o_1 _5732_ (.A1_N(_1195_),
    .A2_N(net41),
    .B1(_2419_),
    .B2(\as2650.r123[2][4] ),
    .X(_2423_));
 sky130_fd_sc_hd__a21o_1 _5733_ (.A1(_0362_),
    .A2(_2418_),
    .B1(_2423_),
    .X(_0266_));
 sky130_fd_sc_hd__nor2_1 _5734_ (.A(_1210_),
    .B(net41),
    .Y(_2424_));
 sky130_fd_sc_hd__a221o_1 _5735_ (.A1(_0415_),
    .A2(_2418_),
    .B1(_2419_),
    .B2(\as2650.r123[2][5] ),
    .C1(_2424_),
    .X(_0267_));
 sky130_fd_sc_hd__a22o_1 _5736_ (.A1(_0459_),
    .A2(_2418_),
    .B1(_2419_),
    .B2(\as2650.r123[2][6] ),
    .X(_2425_));
 sky130_fd_sc_hd__a21o_1 _5737_ (.A1(_1220_),
    .A2(_2407_),
    .B1(_2425_),
    .X(_0268_));
 sky130_fd_sc_hd__a22o_1 _5738_ (.A1(_0495_),
    .A2(_2418_),
    .B1(_2419_),
    .B2(\as2650.r123[2][7] ),
    .X(_2426_));
 sky130_fd_sc_hd__a21o_1 _5739_ (.A1(_1223_),
    .A2(_2407_),
    .B1(_2426_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _5740_ (.A0(net229),
    .A1(net340),
    .S(_0865_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _5741_ (.A0(net228),
    .A1(net337),
    .S(_0865_),
    .X(_0271_));
 sky130_fd_sc_hd__o21ai_1 _5742_ (.A1(net79),
    .A2(net92),
    .B1(_0661_),
    .Y(_2427_));
 sky130_fd_sc_hd__a2111o_1 _5743_ (.A1(net77),
    .A2(net65),
    .B1(_1775_),
    .C1(_1841_),
    .D1(_2620_),
    .X(_2428_));
 sky130_fd_sc_hd__or4b_1 _5744_ (.A(_0781_),
    .B(_1920_),
    .C(_2428_),
    .D_N(_1923_),
    .X(_2429_));
 sky130_fd_sc_hd__and3b_1 _5745_ (.A_N(_1926_),
    .B(_2568_),
    .C(_2603_),
    .X(_2430_));
 sky130_fd_sc_hd__a31o_1 _5746_ (.A1(_2609_),
    .A2(_0642_),
    .A3(_0725_),
    .B1(_2430_),
    .X(_2431_));
 sky130_fd_sc_hd__a311o_1 _5747_ (.A1(net225),
    .A2(net300),
    .A3(_2599_),
    .B1(_2591_),
    .C1(net206),
    .X(_2432_));
 sky130_fd_sc_hd__o221a_1 _5748_ (.A1(net134),
    .A2(net130),
    .B1(net56),
    .B2(net230),
    .C1(_2432_),
    .X(_2433_));
 sky130_fd_sc_hd__or4_1 _5749_ (.A(_2774_),
    .B(_0649_),
    .C(_0711_),
    .D(_0790_),
    .X(_2434_));
 sky130_fd_sc_hd__a31o_1 _5750_ (.A1(_2543_),
    .A2(net308),
    .A3(_0640_),
    .B1(_2689_),
    .X(_2435_));
 sky130_fd_sc_hd__or4_1 _5751_ (.A(_1261_),
    .B(_1298_),
    .C(_2434_),
    .D(_2435_),
    .X(_2436_));
 sky130_fd_sc_hd__or3b_1 _5752_ (.A(_2436_),
    .B(_1873_),
    .C_N(_2433_),
    .X(_2437_));
 sky130_fd_sc_hd__a2111o_4 _5753_ (.A1(net207),
    .A2(_2427_),
    .B1(_2429_),
    .C1(_2431_),
    .D1(_2437_),
    .X(_2438_));
 sky130_fd_sc_hd__a21oi_2 _5754_ (.A1(_2551_),
    .A2(_0794_),
    .B1(_2438_),
    .Y(_2439_));
 sky130_fd_sc_hd__or2_1 _5755_ (.A(_2610_),
    .B(_0793_),
    .X(_2440_));
 sky130_fd_sc_hd__o21ai_1 _5756_ (.A1(_2551_),
    .A2(_0674_),
    .B1(net143),
    .Y(_2441_));
 sky130_fd_sc_hd__nand2_1 _5757_ (.A(net221),
    .B(net169),
    .Y(_2442_));
 sky130_fd_sc_hd__nand2_2 _5758_ (.A(_0679_),
    .B(_2442_),
    .Y(_2443_));
 sky130_fd_sc_hd__mux2_1 _5759_ (.A0(net250),
    .A1(_2443_),
    .S(_2579_),
    .X(_2444_));
 sky130_fd_sc_hd__o31a_1 _5760_ (.A1(net143),
    .A2(net68),
    .A3(_2444_),
    .B1(_2441_),
    .X(_2445_));
 sky130_fd_sc_hd__nor2_1 _5761_ (.A(_2810_),
    .B(_0636_),
    .Y(_2446_));
 sky130_fd_sc_hd__o221a_1 _5762_ (.A1(_0636_),
    .A2(_2445_),
    .B1(_2446_),
    .B2(net107),
    .C1(net207),
    .X(_2447_));
 sky130_fd_sc_hd__a21oi_1 _5763_ (.A1(net229),
    .A2(_2443_),
    .B1(_2447_),
    .Y(_2448_));
 sky130_fd_sc_hd__a21oi_1 _5764_ (.A1(_2439_),
    .A2(_2448_),
    .B1(net348),
    .Y(_2449_));
 sky130_fd_sc_hd__o21a_1 _5765_ (.A1(net221),
    .A2(_2439_),
    .B1(_2449_),
    .X(_0272_));
 sky130_fd_sc_hd__a21oi_1 _5766_ (.A1(_2550_),
    .A2(_0794_),
    .B1(_2438_),
    .Y(_2450_));
 sky130_fd_sc_hd__o21ai_1 _5767_ (.A1(net217),
    .A2(_2450_),
    .B1(net319),
    .Y(_2451_));
 sky130_fd_sc_hd__mux2_1 _5768_ (.A0(net254),
    .A1(_2798_),
    .S(_2579_),
    .X(_2452_));
 sky130_fd_sc_hd__or3_1 _5769_ (.A(net147),
    .B(net68),
    .C(_2452_),
    .X(_2453_));
 sky130_fd_sc_hd__nand2_1 _5770_ (.A(net147),
    .B(_0674_),
    .Y(_2454_));
 sky130_fd_sc_hd__a31o_1 _5771_ (.A1(_1808_),
    .A2(_2453_),
    .A3(_2454_),
    .B1(_0636_),
    .X(_2455_));
 sky130_fd_sc_hd__o31a_1 _5772_ (.A1(net173),
    .A2(_2796_),
    .A3(_2446_),
    .B1(net207),
    .X(_2456_));
 sky130_fd_sc_hd__a22oi_1 _5773_ (.A1(net229),
    .A2(_2798_),
    .B1(_2455_),
    .B2(_2456_),
    .Y(_2457_));
 sky130_fd_sc_hd__a21oi_1 _5774_ (.A1(_2450_),
    .A2(_2457_),
    .B1(_2451_),
    .Y(_0273_));
 sky130_fd_sc_hd__o21ba_1 _5775_ (.A1(net349),
    .A2(_0793_),
    .B1_N(_2438_),
    .X(_2458_));
 sky130_fd_sc_hd__nor2_2 _5776_ (.A(net78),
    .B(_0674_),
    .Y(_2459_));
 sky130_fd_sc_hd__a22oi_2 _5777_ (.A1(_0647_),
    .A2(_1806_),
    .B1(_2459_),
    .B2(net1),
    .Y(_2460_));
 sky130_fd_sc_hd__a211o_1 _5778_ (.A1(_0647_),
    .A2(_0725_),
    .B1(_0794_),
    .C1(net216),
    .X(_2461_));
 sky130_fd_sc_hd__o211ai_1 _5779_ (.A1(net61),
    .A2(_2460_),
    .B1(_2461_),
    .C1(_2458_),
    .Y(_2462_));
 sky130_fd_sc_hd__o211a_1 _5780_ (.A1(net216),
    .A2(_2458_),
    .B1(_2462_),
    .C1(net319),
    .X(_0274_));
 sky130_fd_sc_hd__o22a_1 _5781_ (.A1(net146),
    .A2(_0654_),
    .B1(_0793_),
    .B2(_0631_),
    .X(_2463_));
 sky130_fd_sc_hd__a21oi_1 _5782_ (.A1(net79),
    .A2(net65),
    .B1(_0789_),
    .Y(_2464_));
 sky130_fd_sc_hd__and4b_1 _5783_ (.A_N(_2580_),
    .B(_1275_),
    .C(_2463_),
    .D(_2464_),
    .X(_2465_));
 sky130_fd_sc_hd__o31a_1 _5784_ (.A1(\as2650.psl[3] ),
    .A2(net231),
    .A3(net55),
    .B1(_2465_),
    .X(_2466_));
 sky130_fd_sc_hd__or4_1 _5785_ (.A(net204),
    .B(_0635_),
    .C(_0640_),
    .D(_2440_),
    .X(_2467_));
 sky130_fd_sc_hd__o211a_1 _5786_ (.A1(net195),
    .A2(_2696_),
    .B1(_0718_),
    .C1(_0799_),
    .X(_2468_));
 sky130_fd_sc_hd__and4_1 _5787_ (.A(net52),
    .B(_0801_),
    .C(_1299_),
    .D(_2468_),
    .X(_2469_));
 sky130_fd_sc_hd__and4b_1 _5788_ (.A_N(_0790_),
    .B(_2467_),
    .C(_2469_),
    .D(_0787_),
    .X(_2470_));
 sky130_fd_sc_hd__and3_1 _5789_ (.A(_1295_),
    .B(_2466_),
    .C(_2470_),
    .X(_2471_));
 sky130_fd_sc_hd__o31a_1 _5790_ (.A1(net333),
    .A2(_0633_),
    .A3(_0795_),
    .B1(_2471_),
    .X(_2472_));
 sky130_fd_sc_hd__o21a_1 _5791_ (.A1(_0645_),
    .A2(_0673_),
    .B1(_0631_),
    .X(_2473_));
 sky130_fd_sc_hd__a22o_1 _5792_ (.A1(net101),
    .A2(_0630_),
    .B1(_1817_),
    .B2(_2473_),
    .X(_2474_));
 sky130_fd_sc_hd__mux2_1 _5793_ (.A0(net95),
    .A1(_2474_),
    .S(_2663_),
    .X(_2475_));
 sky130_fd_sc_hd__and2_1 _5794_ (.A(net226),
    .B(_2475_),
    .X(_2476_));
 sky130_fd_sc_hd__o21ai_1 _5795_ (.A1(net227),
    .A2(_0360_),
    .B1(_2472_),
    .Y(_2477_));
 sky130_fd_sc_hd__o221a_1 _5796_ (.A1(\as2650.psl[5] ),
    .A2(_2472_),
    .B1(_2476_),
    .B2(_2477_),
    .C1(net320),
    .X(_0275_));
 sky130_fd_sc_hd__or2_1 _5797_ (.A(_0494_),
    .B(_0756_),
    .X(_2478_));
 sky130_fd_sc_hd__a211o_1 _5798_ (.A1(_2852_),
    .A2(_2854_),
    .B1(_2751_),
    .C1(_2771_),
    .X(_2479_));
 sky130_fd_sc_hd__o21a_1 _5799_ (.A1(_2854_),
    .A2(_2856_),
    .B1(_2479_),
    .X(_2480_));
 sky130_fd_sc_hd__or2_1 _5800_ (.A(_2903_),
    .B(_2480_),
    .X(_2481_));
 sky130_fd_sc_hd__a22o_1 _5801_ (.A1(_0304_),
    .A2(_0309_),
    .B1(_2480_),
    .B2(_2903_),
    .X(_2482_));
 sky130_fd_sc_hd__a31o_1 _5802_ (.A1(_0294_),
    .A2(_0295_),
    .A3(_2481_),
    .B1(_2482_),
    .X(_2483_));
 sky130_fd_sc_hd__o221a_1 _5803_ (.A1(_0304_),
    .A2(_0309_),
    .B1(_0354_),
    .B2(_0361_),
    .C1(_2483_),
    .X(_2484_));
 sky130_fd_sc_hd__a221o_1 _5804_ (.A1(_0354_),
    .A2(_0361_),
    .B1(_0408_),
    .B2(_0414_),
    .C1(_2484_),
    .X(_2485_));
 sky130_fd_sc_hd__o221a_1 _5805_ (.A1(_0408_),
    .A2(_0414_),
    .B1(_0452_),
    .B2(_0458_),
    .C1(_2485_),
    .X(_2486_));
 sky130_fd_sc_hd__nand2_1 _5806_ (.A(_0494_),
    .B(_0756_),
    .Y(_2487_));
 sky130_fd_sc_hd__a221o_1 _5807_ (.A1(_0452_),
    .A2(_0458_),
    .B1(_0494_),
    .B2(_0756_),
    .C1(_2486_),
    .X(_2488_));
 sky130_fd_sc_hd__a21o_1 _5808_ (.A1(_2478_),
    .A2(_2488_),
    .B1(net227),
    .X(_2489_));
 sky130_fd_sc_hd__o31a_2 _5809_ (.A1(net1),
    .A2(_0633_),
    .A3(_0795_),
    .B1(_2471_),
    .X(_2490_));
 sky130_fd_sc_hd__mux2_1 _5810_ (.A0(net114),
    .A1(net110),
    .S(net298),
    .X(_2491_));
 sky130_fd_sc_hd__o21a_1 _5811_ (.A1(_0645_),
    .A2(_1806_),
    .B1(_1807_),
    .X(_2492_));
 sky130_fd_sc_hd__mux2_1 _5812_ (.A0(_2491_),
    .A1(_2492_),
    .S(net55),
    .X(_2493_));
 sky130_fd_sc_hd__nand2_1 _5813_ (.A(net227),
    .B(_2493_),
    .Y(_2494_));
 sky130_fd_sc_hd__a31o_1 _5814_ (.A1(_2489_),
    .A2(_2490_),
    .A3(_2494_),
    .B1(net348),
    .X(_2495_));
 sky130_fd_sc_hd__o21ba_1 _5815_ (.A1(\as2650.carry ),
    .A2(_2490_),
    .B1_N(_2495_),
    .X(_0276_));
 sky130_fd_sc_hd__and2_1 _5816_ (.A(_2478_),
    .B(_2487_),
    .X(_2496_));
 sky130_fd_sc_hd__o22a_1 _5817_ (.A1(net231),
    .A2(net55),
    .B1(_0795_),
    .B2(net343),
    .X(_2497_));
 sky130_fd_sc_hd__and3_1 _5818_ (.A(_0657_),
    .B(_1275_),
    .C(_2497_),
    .X(_2498_));
 sky130_fd_sc_hd__o211ai_1 _5819_ (.A1(_0645_),
    .A2(_1811_),
    .B1(_1812_),
    .C1(net227),
    .Y(_2499_));
 sky130_fd_sc_hd__and3_2 _5820_ (.A(_1295_),
    .B(_2470_),
    .C(_2498_),
    .X(_2500_));
 sky130_fd_sc_hd__o311a_1 _5821_ (.A1(net227),
    .A2(_0481_),
    .A3(_2496_),
    .B1(_2499_),
    .C1(_2500_),
    .X(_2501_));
 sky130_fd_sc_hd__nor2_1 _5822_ (.A(net348),
    .B(_2501_),
    .Y(_2502_));
 sky130_fd_sc_hd__o21a_1 _5823_ (.A1(\as2650.overflow ),
    .A2(_2500_),
    .B1(_2502_),
    .X(_0277_));
 sky130_fd_sc_hd__a211oi_2 _5824_ (.A1(net291),
    .A2(_0641_),
    .B1(_2568_),
    .C1(net293),
    .Y(_2503_));
 sky130_fd_sc_hd__and3b_1 _5825_ (.A_N(_2702_),
    .B(_0800_),
    .C(_2503_),
    .X(_2504_));
 sky130_fd_sc_hd__o2111a_4 _5826_ (.A1(net146),
    .A2(_0783_),
    .B1(_2504_),
    .C1(_0648_),
    .D1(_0652_),
    .X(_2505_));
 sky130_fd_sc_hd__o21ai_1 _5827_ (.A1(net336),
    .A2(net81),
    .B1(_2505_),
    .Y(_2506_));
 sky130_fd_sc_hd__a31o_1 _5828_ (.A1(net336),
    .A2(net144),
    .A3(_0645_),
    .B1(_1815_),
    .X(_2507_));
 sky130_fd_sc_hd__a22o_1 _5829_ (.A1(net213),
    .A2(_2506_),
    .B1(_2507_),
    .B2(_2505_),
    .X(_2508_));
 sky130_fd_sc_hd__and2_1 _5830_ (.A(net320),
    .B(_2508_),
    .X(_0278_));
 sky130_fd_sc_hd__o21ai_1 _5831_ (.A1(net340),
    .A2(net81),
    .B1(_2505_),
    .Y(_2509_));
 sky130_fd_sc_hd__a31o_1 _5832_ (.A1(net340),
    .A2(net144),
    .A3(_0645_),
    .B1(_1813_),
    .X(_2510_));
 sky130_fd_sc_hd__a22o_1 _5833_ (.A1(\as2650.psl[3] ),
    .A2(_2509_),
    .B1(_2510_),
    .B2(_2505_),
    .X(_2511_));
 sky130_fd_sc_hd__and2_1 _5834_ (.A(net320),
    .B(_2511_),
    .X(_0279_));
 sky130_fd_sc_hd__a21oi_1 _5835_ (.A1(_1808_),
    .A2(_2505_),
    .B1(\as2650.psl[1] ),
    .Y(_2512_));
 sky130_fd_sc_hd__a31o_1 _5836_ (.A1(net346),
    .A2(net145),
    .A3(_0644_),
    .B1(_1809_),
    .X(_2513_));
 sky130_fd_sc_hd__a211oi_1 _5837_ (.A1(_2505_),
    .A2(_2513_),
    .B1(_2512_),
    .C1(net348),
    .Y(_0280_));
 sky130_fd_sc_hd__a21o_1 _5838_ (.A1(_0655_),
    .A2(_0658_),
    .B1(net146),
    .X(_2514_));
 sky130_fd_sc_hd__and4b_4 _5839_ (.A_N(net308),
    .B(_2776_),
    .C(_2503_),
    .D(_2514_),
    .X(_2515_));
 sky130_fd_sc_hd__o21ai_1 _5840_ (.A1(net330),
    .A2(net78),
    .B1(_2515_),
    .Y(_2516_));
 sky130_fd_sc_hd__o22ai_1 _5841_ (.A1(net238),
    .A2(net147),
    .B1(_2454_),
    .B2(_2556_),
    .Y(_2517_));
 sky130_fd_sc_hd__a221oi_1 _5842_ (.A1(_2524_),
    .A2(_2516_),
    .B1(_2517_),
    .B2(_2515_),
    .C1(net348),
    .Y(_0281_));
 sky130_fd_sc_hd__o21a_1 _5843_ (.A1(net336),
    .A2(net81),
    .B1(_2515_),
    .X(_2518_));
 sky130_fd_sc_hd__a21o_1 _5844_ (.A1(net336),
    .A2(_2459_),
    .B1(_1815_),
    .X(_2519_));
 sky130_fd_sc_hd__mux2_1 _5845_ (.A0(\as2650.psu[4] ),
    .A1(_2519_),
    .S(_2518_),
    .X(_2520_));
 sky130_fd_sc_hd__and2_1 _5846_ (.A(net319),
    .B(_2520_),
    .X(_0282_));
 sky130_fd_sc_hd__o21a_1 _5847_ (.A1(net340),
    .A2(net81),
    .B1(_2515_),
    .X(_2521_));
 sky130_fd_sc_hd__a21o_1 _5848_ (.A1(net340),
    .A2(_2459_),
    .B1(_1813_),
    .X(_2522_));
 sky130_fd_sc_hd__mux2_1 _5849_ (.A0(\as2650.psu[3] ),
    .A1(_2522_),
    .S(_2521_),
    .X(_2523_));
 sky130_fd_sc_hd__and2_1 _5850_ (.A(net319),
    .B(_2523_),
    .X(_0283_));
 sky130_fd_sc_hd__clkbuf_2 _5851_ (.A(\as2650.r123_2[3][0] ),
    .X(_0098_));
 sky130_fd_sc_hd__clkbuf_2 _5852_ (.A(\as2650.r123_2[3][1] ),
    .X(_0099_));
 sky130_fd_sc_hd__clkbuf_2 _5853_ (.A(\as2650.r123_2[3][2] ),
    .X(_0100_));
 sky130_fd_sc_hd__clkbuf_2 _5854_ (.A(\as2650.r123_2[3][3] ),
    .X(_0101_));
 sky130_fd_sc_hd__clkbuf_2 _5855_ (.A(\as2650.r123_2[3][4] ),
    .X(_0102_));
 sky130_fd_sc_hd__clkbuf_2 _5856_ (.A(\as2650.r123_2[3][5] ),
    .X(_0103_));
 sky130_fd_sc_hd__clkbuf_2 _5857_ (.A(\as2650.r123_2[3][6] ),
    .X(_0104_));
 sky130_fd_sc_hd__clkbuf_2 _5858_ (.A(\as2650.r123_2[3][7] ),
    .X(_0105_));
 sky130_fd_sc_hd__clkbuf_2 _5859_ (.A(\as2650.r123[3][0] ),
    .X(_0146_));
 sky130_fd_sc_hd__clkbuf_2 _5860_ (.A(\as2650.r123[3][1] ),
    .X(_0147_));
 sky130_fd_sc_hd__clkbuf_2 _5861_ (.A(\as2650.r123[3][2] ),
    .X(_0148_));
 sky130_fd_sc_hd__clkbuf_2 _5862_ (.A(\as2650.r123[3][3] ),
    .X(_0149_));
 sky130_fd_sc_hd__clkbuf_2 _5863_ (.A(\as2650.r123[3][4] ),
    .X(_0150_));
 sky130_fd_sc_hd__clkbuf_2 _5864_ (.A(\as2650.r123[3][5] ),
    .X(_0151_));
 sky130_fd_sc_hd__clkbuf_2 _5865_ (.A(\as2650.r123[3][6] ),
    .X(_0152_));
 sky130_fd_sc_hd__clkbuf_2 _5866_ (.A(\as2650.r123[3][7] ),
    .X(_0153_));
 sky130_fd_sc_hd__dfxtp_1 _5867_ (.CLK(clknet_leaf_18_clk),
    .D(_0000_),
    .Q(\as2650.stack[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _5868_ (.CLK(clknet_leaf_21_clk),
    .D(_0001_),
    .Q(\as2650.stack[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _5869_ (.CLK(clknet_leaf_30_clk),
    .D(_0002_),
    .Q(\as2650.stack[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _5870_ (.CLK(clknet_leaf_21_clk),
    .D(_0003_),
    .Q(\as2650.stack[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _5871_ (.CLK(clknet_leaf_23_clk),
    .D(_0004_),
    .Q(\as2650.stack[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _5872_ (.CLK(clknet_leaf_24_clk),
    .D(_0005_),
    .Q(\as2650.stack[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _5873_ (.CLK(clknet_leaf_24_clk),
    .D(_0006_),
    .Q(\as2650.stack[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _5874_ (.CLK(clknet_leaf_11_clk),
    .D(_0007_),
    .Q(\as2650.r123[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5875_ (.CLK(clknet_leaf_14_clk),
    .D(_0008_),
    .Q(\as2650.r123[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5876_ (.CLK(clknet_leaf_15_clk),
    .D(_0009_),
    .Q(\as2650.r123[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5877_ (.CLK(clknet_leaf_19_clk),
    .D(_0010_),
    .Q(\as2650.r123[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5878_ (.CLK(clknet_leaf_17_clk),
    .D(_0011_),
    .Q(\as2650.r123[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5879_ (.CLK(clknet_leaf_19_clk),
    .D(_0012_),
    .Q(\as2650.r123[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5880_ (.CLK(clknet_leaf_13_clk),
    .D(_0013_),
    .Q(\as2650.r123[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5881_ (.CLK(clknet_leaf_14_clk),
    .D(_0014_),
    .Q(\as2650.r123[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5882_ (.CLK(clknet_leaf_18_clk),
    .D(_0015_),
    .Q(\as2650.stack[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _5883_ (.CLK(clknet_leaf_21_clk),
    .D(_0016_),
    .Q(\as2650.stack[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _5884_ (.CLK(clknet_leaf_17_clk),
    .D(_0017_),
    .Q(\as2650.stack[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _5885_ (.CLK(clknet_leaf_21_clk),
    .D(_0018_),
    .Q(\as2650.stack[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _5886_ (.CLK(clknet_leaf_24_clk),
    .D(_0019_),
    .Q(\as2650.stack[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _5887_ (.CLK(clknet_leaf_24_clk),
    .D(_0020_),
    .Q(\as2650.stack[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _5888_ (.CLK(clknet_leaf_24_clk),
    .D(_0021_),
    .Q(\as2650.stack[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _5889_ (.CLK(clknet_leaf_37_clk),
    .D(_0022_),
    .Q(\as2650.stack[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5890_ (.CLK(clknet_leaf_37_clk),
    .D(_0023_),
    .Q(\as2650.stack[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5891_ (.CLK(clknet_leaf_36_clk),
    .D(_0024_),
    .Q(\as2650.stack[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5892_ (.CLK(clknet_leaf_38_clk),
    .D(_0025_),
    .Q(\as2650.stack[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5893_ (.CLK(clknet_leaf_37_clk),
    .D(_0026_),
    .Q(\as2650.stack[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5894_ (.CLK(clknet_leaf_40_clk),
    .D(_0027_),
    .Q(\as2650.stack[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5895_ (.CLK(clknet_leaf_38_clk),
    .D(_0028_),
    .Q(\as2650.stack[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5896_ (.CLK(clknet_leaf_39_clk),
    .D(_0029_),
    .Q(\as2650.stack[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5897_ (.CLK(clknet_leaf_18_clk),
    .D(_0030_),
    .Q(\as2650.stack[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _5898_ (.CLK(clknet_leaf_22_clk),
    .D(_0031_),
    .Q(\as2650.stack[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _5899_ (.CLK(clknet_leaf_18_clk),
    .D(_0032_),
    .Q(\as2650.stack[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _5900_ (.CLK(clknet_leaf_22_clk),
    .D(_0033_),
    .Q(\as2650.stack[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _5901_ (.CLK(clknet_leaf_23_clk),
    .D(_0034_),
    .Q(\as2650.stack[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _5902_ (.CLK(clknet_leaf_24_clk),
    .D(_0035_),
    .Q(\as2650.stack[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _5903_ (.CLK(clknet_leaf_22_clk),
    .D(_0036_),
    .Q(\as2650.stack[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _5904_ (.CLK(clknet_leaf_15_clk),
    .D(_0037_),
    .Q(\as2650.r123_2[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5905_ (.CLK(clknet_leaf_14_clk),
    .D(_0038_),
    .Q(\as2650.r123_2[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5906_ (.CLK(clknet_leaf_15_clk),
    .D(_0039_),
    .Q(\as2650.r123_2[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5907_ (.CLK(clknet_leaf_14_clk),
    .D(_0040_),
    .Q(\as2650.r123_2[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5908_ (.CLK(clknet_leaf_17_clk),
    .D(_0041_),
    .Q(\as2650.r123_2[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5909_ (.CLK(clknet_leaf_19_clk),
    .D(_0042_),
    .Q(\as2650.r123_2[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5910_ (.CLK(clknet_leaf_14_clk),
    .D(_0043_),
    .Q(\as2650.r123_2[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5911_ (.CLK(clknet_leaf_14_clk),
    .D(_0044_),
    .Q(\as2650.r123_2[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5912_ (.CLK(clknet_leaf_6_clk),
    .D(_0045_),
    .Q(\as2650.psu[5] ));
 sky130_fd_sc_hd__dfxtp_1 _5913_ (.CLK(clknet_leaf_25_clk),
    .D(_0046_),
    .Q(\as2650.stack[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _5914_ (.CLK(clknet_leaf_22_clk),
    .D(_0047_),
    .Q(\as2650.stack[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _5915_ (.CLK(clknet_leaf_30_clk),
    .D(_0048_),
    .Q(\as2650.stack[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _5916_ (.CLK(clknet_leaf_21_clk),
    .D(_0049_),
    .Q(\as2650.stack[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _5917_ (.CLK(clknet_leaf_25_clk),
    .D(_0050_),
    .Q(\as2650.stack[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _5918_ (.CLK(clknet_leaf_25_clk),
    .D(_0051_),
    .Q(\as2650.stack[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _5919_ (.CLK(clknet_leaf_25_clk),
    .D(_0052_),
    .Q(\as2650.stack[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _5920_ (.CLK(clknet_leaf_39_clk),
    .D(_0053_),
    .Q(net12));
 sky130_fd_sc_hd__dfxtp_1 _5921_ (.CLK(clknet_leaf_38_clk),
    .D(_0054_),
    .Q(net23));
 sky130_fd_sc_hd__dfxtp_1 _5922_ (.CLK(clknet_leaf_39_clk),
    .D(_0055_),
    .Q(net31));
 sky130_fd_sc_hd__dfxtp_1 _5923_ (.CLK(clknet_leaf_39_clk),
    .D(_0056_),
    .Q(net32));
 sky130_fd_sc_hd__dfxtp_1 _5924_ (.CLK(clknet_leaf_40_clk),
    .D(_0057_),
    .Q(net33));
 sky130_fd_sc_hd__dfxtp_1 _5925_ (.CLK(clknet_leaf_40_clk),
    .D(_0058_),
    .Q(net34));
 sky130_fd_sc_hd__dfxtp_1 _5926_ (.CLK(clknet_leaf_40_clk),
    .D(_0059_),
    .Q(net35));
 sky130_fd_sc_hd__dfxtp_1 _5927_ (.CLK(clknet_leaf_40_clk),
    .D(_0060_),
    .Q(net36));
 sky130_fd_sc_hd__dfxtp_1 _5928_ (.CLK(clknet_leaf_30_clk),
    .D(_0061_),
    .Q(\as2650.stack[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _5929_ (.CLK(clknet_leaf_25_clk),
    .D(_0062_),
    .Q(\as2650.stack[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _5930_ (.CLK(clknet_leaf_30_clk),
    .D(_0063_),
    .Q(\as2650.stack[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _5931_ (.CLK(clknet_leaf_18_clk),
    .D(_0064_),
    .Q(\as2650.stack[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _5932_ (.CLK(clknet_leaf_25_clk),
    .D(_0065_),
    .Q(\as2650.stack[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _5933_ (.CLK(clknet_leaf_26_clk),
    .D(_0066_),
    .Q(\as2650.stack[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _5934_ (.CLK(clknet_leaf_25_clk),
    .D(_0067_),
    .Q(\as2650.stack[2][14] ));
 sky130_fd_sc_hd__dfxtp_2 _5935_ (.CLK(clknet_leaf_7_clk),
    .D(_0068_),
    .Q(\as2650.psl[6] ));
 sky130_fd_sc_hd__dfxtp_2 _5936_ (.CLK(clknet_leaf_7_clk),
    .D(_0069_),
    .Q(\as2650.psl[7] ));
 sky130_fd_sc_hd__dfxtp_1 _5937_ (.CLK(clknet_leaf_25_clk),
    .D(_0070_),
    .Q(\as2650.stack[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _5938_ (.CLK(clknet_leaf_24_clk),
    .D(_0071_),
    .Q(\as2650.stack[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _5939_ (.CLK(clknet_leaf_29_clk),
    .D(_0072_),
    .Q(\as2650.stack[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _5940_ (.CLK(clknet_leaf_21_clk),
    .D(_0073_),
    .Q(\as2650.stack[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _5941_ (.CLK(clknet_leaf_26_clk),
    .D(_0074_),
    .Q(\as2650.stack[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _5942_ (.CLK(clknet_leaf_26_clk),
    .D(_0075_),
    .Q(\as2650.stack[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _5943_ (.CLK(clknet_leaf_24_clk),
    .D(_0076_),
    .Q(\as2650.stack[1][14] ));
 sky130_fd_sc_hd__dfxtp_2 _5944_ (.CLK(clknet_leaf_5_clk),
    .D(_0077_),
    .Q(\as2650.ins_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _5945_ (.CLK(clknet_leaf_5_clk),
    .D(_0078_),
    .Q(\as2650.ins_reg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _5946_ (.CLK(clknet_leaf_5_clk),
    .D(_0079_),
    .Q(\as2650.ins_reg[2] ));
 sky130_fd_sc_hd__dfxtp_4 _5947_ (.CLK(clknet_leaf_5_clk),
    .D(_0080_),
    .Q(\as2650.ins_reg[5] ));
 sky130_fd_sc_hd__dfxtp_4 _5948_ (.CLK(clknet_leaf_5_clk),
    .D(_0081_),
    .Q(\as2650.ins_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _5949_ (.CLK(clknet_leaf_5_clk),
    .D(_0082_),
    .Q(\as2650.ins_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _5950_ (.CLK(clknet_leaf_25_clk),
    .D(_0083_),
    .Q(\as2650.stack[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _5951_ (.CLK(clknet_leaf_24_clk),
    .D(_0084_),
    .Q(\as2650.stack[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _5952_ (.CLK(clknet_leaf_29_clk),
    .D(_0085_),
    .Q(\as2650.stack[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _5953_ (.CLK(clknet_leaf_21_clk),
    .D(_0086_),
    .Q(\as2650.stack[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _5954_ (.CLK(clknet_leaf_26_clk),
    .D(_0087_),
    .Q(\as2650.stack[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _5955_ (.CLK(clknet_leaf_26_clk),
    .D(_0088_),
    .Q(\as2650.stack[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _5956_ (.CLK(clknet_leaf_24_clk),
    .D(_0089_),
    .Q(\as2650.stack[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _5957_ (.CLK(clknet_leaf_11_clk),
    .D(_0090_),
    .Q(\as2650.r123_2[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5958_ (.CLK(clknet_leaf_10_clk),
    .D(_0091_),
    .Q(\as2650.r123_2[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5959_ (.CLK(clknet_leaf_12_clk),
    .D(_0092_),
    .Q(\as2650.r123_2[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5960_ (.CLK(clknet_leaf_10_clk),
    .D(_0093_),
    .Q(\as2650.r123_2[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5961_ (.CLK(clknet_leaf_10_clk),
    .D(_0094_),
    .Q(\as2650.r123_2[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5962_ (.CLK(clknet_leaf_11_clk),
    .D(_0095_),
    .Q(\as2650.r123_2[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5963_ (.CLK(clknet_leaf_12_clk),
    .D(_0096_),
    .Q(\as2650.r123_2[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5964_ (.CLK(clknet_leaf_12_clk),
    .D(_0097_),
    .Q(\as2650.r123_2[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5965_ (.CLK(clknet_leaf_23_clk),
    .D(_0098_),
    .Q(\as2650.r123_2[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5966_ (.CLK(clknet_leaf_22_clk),
    .D(_0099_),
    .Q(\as2650.r123_2[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5967_ (.CLK(clknet_leaf_23_clk),
    .D(_0100_),
    .Q(\as2650.r123_2[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5968_ (.CLK(clknet_leaf_23_clk),
    .D(_0101_),
    .Q(\as2650.r123_2[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5969_ (.CLK(clknet_leaf_22_clk),
    .D(_0102_),
    .Q(\as2650.r123_2[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5970_ (.CLK(clknet_leaf_22_clk),
    .D(_0103_),
    .Q(\as2650.r123_2[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5971_ (.CLK(clknet_leaf_21_clk),
    .D(_0104_),
    .Q(\as2650.r123_2[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5972_ (.CLK(clknet_leaf_22_clk),
    .D(_0105_),
    .Q(\as2650.r123_2[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5973_ (.CLK(clknet_leaf_28_clk),
    .D(_0106_),
    .Q(\as2650.stack[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5974_ (.CLK(clknet_leaf_28_clk),
    .D(_0107_),
    .Q(\as2650.stack[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5975_ (.CLK(clknet_leaf_27_clk),
    .D(_0108_),
    .Q(\as2650.stack[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5976_ (.CLK(clknet_leaf_33_clk),
    .D(_0109_),
    .Q(\as2650.stack[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5977_ (.CLK(clknet_leaf_35_clk),
    .D(_0110_),
    .Q(\as2650.stack[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5978_ (.CLK(clknet_leaf_32_clk),
    .D(_0111_),
    .Q(\as2650.stack[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5979_ (.CLK(clknet_leaf_33_clk),
    .D(_0112_),
    .Q(\as2650.stack[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5980_ (.CLK(clknet_leaf_35_clk),
    .D(_0113_),
    .Q(\as2650.stack[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5981_ (.CLK(clknet_leaf_12_clk),
    .D(_0114_),
    .Q(\as2650.r123_2[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5982_ (.CLK(clknet_leaf_12_clk),
    .D(_0115_),
    .Q(\as2650.r123_2[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5983_ (.CLK(clknet_leaf_13_clk),
    .D(_0116_),
    .Q(\as2650.r123_2[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5984_ (.CLK(clknet_leaf_13_clk),
    .D(_0117_),
    .Q(\as2650.r123_2[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5985_ (.CLK(clknet_leaf_19_clk),
    .D(_0118_),
    .Q(\as2650.r123_2[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5986_ (.CLK(clknet_leaf_19_clk),
    .D(_0119_),
    .Q(\as2650.r123_2[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5987_ (.CLK(clknet_leaf_13_clk),
    .D(_0120_),
    .Q(\as2650.r123_2[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5988_ (.CLK(clknet_leaf_13_clk),
    .D(_0121_),
    .Q(\as2650.r123_2[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5989_ (.CLK(clknet_leaf_37_clk),
    .D(_0122_),
    .Q(\as2650.stack[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5990_ (.CLK(clknet_leaf_37_clk),
    .D(_0123_),
    .Q(\as2650.stack[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5991_ (.CLK(clknet_leaf_35_clk),
    .D(_0124_),
    .Q(\as2650.stack[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5992_ (.CLK(clknet_leaf_38_clk),
    .D(_0125_),
    .Q(\as2650.stack[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5993_ (.CLK(clknet_leaf_36_clk),
    .D(_0126_),
    .Q(\as2650.stack[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5994_ (.CLK(clknet_leaf_40_clk),
    .D(_0127_),
    .Q(\as2650.stack[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5995_ (.CLK(clknet_leaf_38_clk),
    .D(_0128_),
    .Q(\as2650.stack[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5996_ (.CLK(clknet_leaf_38_clk),
    .D(_0129_),
    .Q(\as2650.stack[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5997_ (.CLK(clknet_leaf_29_clk),
    .D(_0130_),
    .Q(\as2650.stack[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5998_ (.CLK(clknet_leaf_27_clk),
    .D(_0131_),
    .Q(\as2650.stack[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5999_ (.CLK(clknet_leaf_27_clk),
    .D(_0132_),
    .Q(\as2650.stack[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6000_ (.CLK(clknet_leaf_27_clk),
    .D(_0133_),
    .Q(\as2650.stack[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6001_ (.CLK(clknet_leaf_35_clk),
    .D(_0134_),
    .Q(\as2650.stack[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6002_ (.CLK(clknet_leaf_32_clk),
    .D(_0135_),
    .Q(\as2650.stack[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6003_ (.CLK(clknet_leaf_34_clk),
    .D(_0136_),
    .Q(\as2650.stack[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6004_ (.CLK(clknet_leaf_35_clk),
    .D(_0137_),
    .Q(\as2650.stack[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6005_ (.CLK(clknet_leaf_29_clk),
    .D(_0138_),
    .Q(\as2650.stack[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6006_ (.CLK(clknet_leaf_28_clk),
    .D(_0139_),
    .Q(\as2650.stack[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6007_ (.CLK(clknet_leaf_26_clk),
    .D(_0140_),
    .Q(\as2650.stack[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6008_ (.CLK(clknet_leaf_26_clk),
    .D(_0141_),
    .Q(\as2650.stack[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6009_ (.CLK(clknet_leaf_34_clk),
    .D(_0142_),
    .Q(\as2650.stack[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6010_ (.CLK(clknet_leaf_33_clk),
    .D(_0143_),
    .Q(\as2650.stack[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6011_ (.CLK(clknet_leaf_27_clk),
    .D(_0144_),
    .Q(\as2650.stack[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6012_ (.CLK(clknet_leaf_33_clk),
    .D(_0145_),
    .Q(\as2650.stack[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6013_ (.CLK(clknet_leaf_23_clk),
    .D(_0146_),
    .Q(\as2650.r123[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6014_ (.CLK(clknet_leaf_23_clk),
    .D(_0147_),
    .Q(\as2650.r123[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6015_ (.CLK(clknet_leaf_23_clk),
    .D(_0148_),
    .Q(\as2650.r123[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6016_ (.CLK(clknet_leaf_23_clk),
    .D(_0149_),
    .Q(\as2650.r123[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6017_ (.CLK(clknet_leaf_23_clk),
    .D(_0150_),
    .Q(\as2650.r123[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6018_ (.CLK(clknet_leaf_22_clk),
    .D(_0151_),
    .Q(\as2650.r123[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6019_ (.CLK(clknet_leaf_22_clk),
    .D(_0152_),
    .Q(\as2650.r123[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6020_ (.CLK(clknet_leaf_23_clk),
    .D(_0153_),
    .Q(\as2650.r123[3][7] ));
 sky130_fd_sc_hd__dfxtp_2 _6021_ (.CLK(clknet_leaf_0_clk),
    .D(_0154_),
    .Q(\as2650.addr_buff[0] ));
 sky130_fd_sc_hd__dfxtp_2 _6022_ (.CLK(clknet_leaf_0_clk),
    .D(_0155_),
    .Q(\as2650.addr_buff[1] ));
 sky130_fd_sc_hd__dfxtp_4 _6023_ (.CLK(clknet_leaf_0_clk),
    .D(_0156_),
    .Q(\as2650.addr_buff[2] ));
 sky130_fd_sc_hd__dfxtp_4 _6024_ (.CLK(clknet_leaf_1_clk),
    .D(_0157_),
    .Q(\as2650.addr_buff[3] ));
 sky130_fd_sc_hd__dfxtp_4 _6025_ (.CLK(clknet_leaf_1_clk),
    .D(_0158_),
    .Q(\as2650.addr_buff[4] ));
 sky130_fd_sc_hd__dfxtp_4 _6026_ (.CLK(clknet_leaf_3_clk),
    .D(_0159_),
    .Q(\as2650.addr_buff[5] ));
 sky130_fd_sc_hd__dfxtp_4 _6027_ (.CLK(clknet_leaf_3_clk),
    .D(_0160_),
    .Q(\as2650.addr_buff[6] ));
 sky130_fd_sc_hd__dfxtp_4 _6028_ (.CLK(clknet_leaf_3_clk),
    .D(_0161_),
    .Q(\as2650.addr_buff[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6029_ (.CLK(clknet_leaf_28_clk),
    .D(_0162_),
    .Q(\as2650.stack[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6030_ (.CLK(clknet_leaf_25_clk),
    .D(_0163_),
    .Q(\as2650.stack[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6031_ (.CLK(clknet_leaf_27_clk),
    .D(_0164_),
    .Q(\as2650.stack[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6032_ (.CLK(clknet_leaf_27_clk),
    .D(_0165_),
    .Q(\as2650.stack[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6033_ (.CLK(clknet_leaf_34_clk),
    .D(_0166_),
    .Q(\as2650.stack[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6034_ (.CLK(clknet_leaf_33_clk),
    .D(_0167_),
    .Q(\as2650.stack[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6035_ (.CLK(clknet_leaf_34_clk),
    .D(_0168_),
    .Q(\as2650.stack[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6036_ (.CLK(clknet_leaf_33_clk),
    .D(_0169_),
    .Q(\as2650.stack[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6037_ (.CLK(clknet_leaf_3_clk),
    .D(_0170_),
    .Q(net27));
 sky130_fd_sc_hd__dfxtp_1 _6038_ (.CLK(clknet_leaf_2_clk),
    .D(_0171_),
    .Q(net29));
 sky130_fd_sc_hd__dfxtp_1 _6039_ (.CLK(clknet_leaf_2_clk),
    .D(_0172_),
    .Q(net28));
 sky130_fd_sc_hd__dfxtp_4 _6040_ (.CLK(clknet_leaf_41_clk),
    .D(_0173_),
    .Q(net37));
 sky130_fd_sc_hd__dfxtp_4 _6041_ (.CLK(clknet_leaf_41_clk),
    .D(_0174_),
    .Q(net38));
 sky130_fd_sc_hd__dfxtp_2 _6042_ (.CLK(clknet_leaf_41_clk),
    .D(_0175_),
    .Q(net13));
 sky130_fd_sc_hd__dfxtp_4 _6043_ (.CLK(clknet_leaf_41_clk),
    .D(_0176_),
    .Q(net14));
 sky130_fd_sc_hd__dfxtp_4 _6044_ (.CLK(clknet_leaf_40_clk),
    .D(_0177_),
    .Q(net15));
 sky130_fd_sc_hd__dfxtp_2 _6045_ (.CLK(clknet_leaf_41_clk),
    .D(_0178_),
    .Q(net16));
 sky130_fd_sc_hd__dfxtp_4 _6046_ (.CLK(clknet_leaf_41_clk),
    .D(_0179_),
    .Q(net17));
 sky130_fd_sc_hd__dfxtp_4 _6047_ (.CLK(clknet_leaf_42_clk),
    .D(_0180_),
    .Q(net18));
 sky130_fd_sc_hd__dfxtp_4 _6048_ (.CLK(clknet_leaf_42_clk),
    .D(_0181_),
    .Q(net19));
 sky130_fd_sc_hd__dfxtp_2 _6049_ (.CLK(clknet_leaf_0_clk),
    .D(_0182_),
    .Q(net20));
 sky130_fd_sc_hd__dfxtp_4 _6050_ (.CLK(clknet_leaf_0_clk),
    .D(_0183_),
    .Q(net21));
 sky130_fd_sc_hd__dfxtp_2 _6051_ (.CLK(clknet_leaf_0_clk),
    .D(_0184_),
    .Q(net22));
 sky130_fd_sc_hd__dfxtp_4 _6052_ (.CLK(clknet_leaf_0_clk),
    .D(_0185_),
    .Q(net24));
 sky130_fd_sc_hd__dfxtp_1 _6053_ (.CLK(clknet_leaf_2_clk),
    .D(_0186_),
    .Q(net25));
 sky130_fd_sc_hd__dfxtp_4 _6054_ (.CLK(clknet_leaf_2_clk),
    .D(_0187_),
    .Q(net26));
 sky130_fd_sc_hd__dfxtp_4 _6055_ (.CLK(clknet_leaf_4_clk),
    .D(_0188_),
    .Q(\as2650.idx_ctrl[0] ));
 sky130_fd_sc_hd__dfxtp_4 _6056_ (.CLK(clknet_leaf_4_clk),
    .D(_0189_),
    .Q(\as2650.idx_ctrl[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6057_ (.CLK(clknet_leaf_7_clk),
    .D(_0190_),
    .Q(\as2650.holding_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6058_ (.CLK(clknet_leaf_7_clk),
    .D(_0191_),
    .Q(\as2650.holding_reg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _6059_ (.CLK(clknet_leaf_9_clk),
    .D(_0192_),
    .Q(\as2650.holding_reg[2] ));
 sky130_fd_sc_hd__dfxtp_4 _6060_ (.CLK(clknet_leaf_9_clk),
    .D(_0193_),
    .Q(\as2650.holding_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6061_ (.CLK(clknet_leaf_9_clk),
    .D(_0194_),
    .Q(\as2650.holding_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6062_ (.CLK(clknet_leaf_9_clk),
    .D(_0195_),
    .Q(\as2650.holding_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6063_ (.CLK(clknet_leaf_9_clk),
    .D(_0196_),
    .Q(\as2650.holding_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6064_ (.CLK(clknet_leaf_9_clk),
    .D(_0197_),
    .Q(\as2650.holding_reg[7] ));
 sky130_fd_sc_hd__dfxtp_4 _6065_ (.CLK(clknet_leaf_3_clk),
    .D(_0198_),
    .Q(\as2650.halted ));
 sky130_fd_sc_hd__dfxtp_2 _6066_ (.CLK(clknet_leaf_2_clk),
    .D(_0199_),
    .Q(\as2650.cycle[0] ));
 sky130_fd_sc_hd__dfxtp_4 _6067_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0200_),
    .Q(\as2650.cycle[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6068_ (.CLK(clknet_leaf_2_clk),
    .D(_0201_),
    .Q(\as2650.cycle[2] ));
 sky130_fd_sc_hd__dfxtp_4 _6069_ (.CLK(clknet_leaf_2_clk),
    .D(_0202_),
    .Q(\as2650.cycle[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6070_ (.CLK(clknet_leaf_2_clk),
    .D(_0203_),
    .Q(\as2650.cycle[4] ));
 sky130_fd_sc_hd__dfxtp_2 _6071_ (.CLK(clknet_leaf_2_clk),
    .D(_0204_),
    .Q(\as2650.cycle[5] ));
 sky130_fd_sc_hd__dfxtp_4 _6072_ (.CLK(clknet_leaf_3_clk),
    .D(_0205_),
    .Q(\as2650.cycle[6] ));
 sky130_fd_sc_hd__dfxtp_4 _6073_ (.CLK(clknet_leaf_3_clk),
    .D(_0206_),
    .Q(\as2650.cycle[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6074_ (.CLK(clknet_leaf_5_clk),
    .D(_0207_),
    .Q(\as2650.psu[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6075_ (.CLK(clknet_leaf_32_clk),
    .D(_0208_),
    .Q(\as2650.pc[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6076_ (.CLK(clknet_leaf_16_clk),
    .D(_0209_),
    .Q(\as2650.pc[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6077_ (.CLK(clknet_leaf_32_clk),
    .D(_0210_),
    .Q(\as2650.pc[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6078_ (.CLK(clknet_leaf_31_clk),
    .D(_0211_),
    .Q(\as2650.pc[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6079_ (.CLK(clknet_leaf_32_clk),
    .D(_0212_),
    .Q(\as2650.pc[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6080_ (.CLK(clknet_leaf_32_clk),
    .D(_0213_),
    .Q(\as2650.pc[5] ));
 sky130_fd_sc_hd__dfxtp_2 _6081_ (.CLK(clknet_leaf_29_clk),
    .D(_0214_),
    .Q(\as2650.pc[6] ));
 sky130_fd_sc_hd__dfxtp_2 _6082_ (.CLK(clknet_leaf_31_clk),
    .D(_0215_),
    .Q(\as2650.pc[7] ));
 sky130_fd_sc_hd__dfxtp_2 _6083_ (.CLK(clknet_leaf_16_clk),
    .D(_0216_),
    .Q(\as2650.pc[8] ));
 sky130_fd_sc_hd__dfxtp_4 _6084_ (.CLK(clknet_leaf_5_clk),
    .D(_0217_),
    .Q(\as2650.pc[9] ));
 sky130_fd_sc_hd__dfxtp_2 _6085_ (.CLK(clknet_leaf_16_clk),
    .D(_0218_),
    .Q(\as2650.pc[10] ));
 sky130_fd_sc_hd__dfxtp_2 _6086_ (.CLK(clknet_leaf_16_clk),
    .D(_0219_),
    .Q(\as2650.pc[11] ));
 sky130_fd_sc_hd__dfxtp_2 _6087_ (.CLK(clknet_leaf_16_clk),
    .D(_0220_),
    .Q(\as2650.pc[12] ));
 sky130_fd_sc_hd__dfxtp_4 _6088_ (.CLK(clknet_leaf_31_clk),
    .D(_0221_),
    .Q(\as2650.pc[13] ));
 sky130_fd_sc_hd__dfxtp_4 _6089_ (.CLK(clknet_leaf_31_clk),
    .D(_0222_),
    .Q(\as2650.pc[14] ));
 sky130_fd_sc_hd__dfxtp_1 _6090_ (.CLK(clknet_leaf_4_clk),
    .D(_0223_),
    .Q(\as2650.r0[0] ));
 sky130_fd_sc_hd__dfxtp_4 _6091_ (.CLK(clknet_leaf_4_clk),
    .D(_0224_),
    .Q(\as2650.r0[1] ));
 sky130_fd_sc_hd__dfxtp_4 _6092_ (.CLK(clknet_leaf_4_clk),
    .D(_0225_),
    .Q(\as2650.r0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6093_ (.CLK(clknet_leaf_4_clk),
    .D(_0226_),
    .Q(\as2650.r0[3] ));
 sky130_fd_sc_hd__dfxtp_4 _6094_ (.CLK(clknet_leaf_4_clk),
    .D(_0227_),
    .Q(\as2650.r0[4] ));
 sky130_fd_sc_hd__dfxtp_4 _6095_ (.CLK(clknet_leaf_4_clk),
    .D(_0228_),
    .Q(\as2650.r0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6096_ (.CLK(clknet_leaf_4_clk),
    .D(_0229_),
    .Q(\as2650.r0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6097_ (.CLK(clknet_leaf_4_clk),
    .D(_0230_),
    .Q(\as2650.r0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6098_ (.CLK(clknet_leaf_37_clk),
    .D(_0231_),
    .Q(\as2650.stack[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6099_ (.CLK(clknet_leaf_37_clk),
    .D(_0232_),
    .Q(\as2650.stack[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6100_ (.CLK(clknet_leaf_36_clk),
    .D(_0233_),
    .Q(\as2650.stack[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6101_ (.CLK(clknet_leaf_38_clk),
    .D(_0234_),
    .Q(\as2650.stack[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6102_ (.CLK(clknet_leaf_37_clk),
    .D(_0235_),
    .Q(\as2650.stack[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6103_ (.CLK(clknet_leaf_40_clk),
    .D(_0236_),
    .Q(\as2650.stack[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6104_ (.CLK(clknet_leaf_38_clk),
    .D(_0237_),
    .Q(\as2650.stack[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6105_ (.CLK(clknet_leaf_39_clk),
    .D(_0238_),
    .Q(\as2650.stack[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6106_ (.CLK(clknet_leaf_37_clk),
    .D(_0239_),
    .Q(\as2650.stack[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6107_ (.CLK(clknet_leaf_37_clk),
    .D(_0240_),
    .Q(\as2650.stack[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6108_ (.CLK(clknet_leaf_35_clk),
    .D(_0241_),
    .Q(\as2650.stack[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6109_ (.CLK(clknet_leaf_38_clk),
    .D(_0242_),
    .Q(\as2650.stack[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6110_ (.CLK(clknet_leaf_35_clk),
    .D(_0243_),
    .Q(\as2650.stack[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6111_ (.CLK(clknet_leaf_37_clk),
    .D(_0244_),
    .Q(\as2650.stack[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6112_ (.CLK(clknet_leaf_38_clk),
    .D(_0245_),
    .Q(\as2650.stack[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6113_ (.CLK(clknet_leaf_38_clk),
    .D(_0246_),
    .Q(\as2650.stack[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6114_ (.CLK(clknet_leaf_21_clk),
    .D(_0247_),
    .Q(\as2650.stack[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6115_ (.CLK(clknet_leaf_22_clk),
    .D(_0248_),
    .Q(\as2650.stack[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6116_ (.CLK(clknet_leaf_17_clk),
    .D(_0249_),
    .Q(\as2650.stack[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6117_ (.CLK(clknet_leaf_21_clk),
    .D(_0250_),
    .Q(\as2650.stack[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6118_ (.CLK(clknet_leaf_23_clk),
    .D(_0251_),
    .Q(\as2650.stack[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6119_ (.CLK(clknet_leaf_24_clk),
    .D(_0252_),
    .Q(\as2650.stack[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _6120_ (.CLK(clknet_leaf_22_clk),
    .D(_0253_),
    .Q(\as2650.stack[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _6121_ (.CLK(clknet_leaf_11_clk),
    .D(_0254_),
    .Q(\as2650.r123[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6122_ (.CLK(clknet_leaf_9_clk),
    .D(_0255_),
    .Q(\as2650.r123[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6123_ (.CLK(clknet_leaf_12_clk),
    .D(_0256_),
    .Q(\as2650.r123[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6124_ (.CLK(clknet_leaf_10_clk),
    .D(_0257_),
    .Q(\as2650.r123[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6125_ (.CLK(clknet_leaf_10_clk),
    .D(_0258_),
    .Q(\as2650.r123[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6126_ (.CLK(clknet_leaf_11_clk),
    .D(_0259_),
    .Q(\as2650.r123[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6127_ (.CLK(clknet_leaf_12_clk),
    .D(_0260_),
    .Q(\as2650.r123[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6128_ (.CLK(clknet_leaf_12_clk),
    .D(_0261_),
    .Q(\as2650.r123[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6129_ (.CLK(clknet_leaf_12_clk),
    .D(_0262_),
    .Q(\as2650.r123[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6130_ (.CLK(clknet_leaf_13_clk),
    .D(_0263_),
    .Q(\as2650.r123[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6131_ (.CLK(clknet_leaf_13_clk),
    .D(_0264_),
    .Q(\as2650.r123[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6132_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0265_),
    .Q(\as2650.r123[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6133_ (.CLK(clknet_leaf_19_clk),
    .D(_0266_),
    .Q(\as2650.r123[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6134_ (.CLK(clknet_leaf_19_clk),
    .D(_0267_),
    .Q(\as2650.r123[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6135_ (.CLK(clknet_leaf_13_clk),
    .D(_0268_),
    .Q(\as2650.r123[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6136_ (.CLK(clknet_leaf_13_clk),
    .D(_0269_),
    .Q(\as2650.r123[2][7] ));
 sky130_fd_sc_hd__dfxtp_4 _6137_ (.CLK(clknet_leaf_5_clk),
    .D(_0270_),
    .Q(\as2650.ins_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6138_ (.CLK(clknet_leaf_5_clk),
    .D(_0271_),
    .Q(\as2650.ins_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6139_ (.CLK(clknet_leaf_15_clk),
    .D(_0272_),
    .Q(\as2650.psu[2] ));
 sky130_fd_sc_hd__dfxtp_2 _6140_ (.CLK(clknet_leaf_15_clk),
    .D(_0273_),
    .Q(\as2650.psu[1] ));
 sky130_fd_sc_hd__dfxtp_2 _6141_ (.CLK(clknet_leaf_15_clk),
    .D(_0274_),
    .Q(\as2650.psu[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6142_ (.CLK(clknet_leaf_7_clk),
    .D(_0275_),
    .Q(\as2650.psl[5] ));
 sky130_fd_sc_hd__dfxtp_2 _6143_ (.CLK(clknet_leaf_7_clk),
    .D(_0276_),
    .Q(\as2650.carry ));
 sky130_fd_sc_hd__dfxtp_1 _6144_ (.CLK(clknet_leaf_8_clk),
    .D(_0277_),
    .Q(\as2650.overflow ));
 sky130_fd_sc_hd__dfxtp_2 _6145_ (.CLK(clknet_leaf_8_clk),
    .D(_0278_),
    .Q(\as2650.psl[4] ));
 sky130_fd_sc_hd__dfxtp_4 _6146_ (.CLK(clknet_leaf_8_clk),
    .D(_0279_),
    .Q(\as2650.psl[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6147_ (.CLK(clknet_leaf_8_clk),
    .D(_0280_),
    .Q(\as2650.psl[1] ));
 sky130_fd_sc_hd__dfxtp_4 _6148_ (.CLK(clknet_leaf_15_clk),
    .D(_0281_),
    .Q(net30));
 sky130_fd_sc_hd__dfxtp_1 _6149_ (.CLK(clknet_leaf_6_clk),
    .D(_0282_),
    .Q(\as2650.psu[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6150_ (.CLK(clknet_leaf_8_clk),
    .D(_0283_),
    .Q(\as2650.psu[3] ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__buf_12 input1 (.A(io_in[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(io_in[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(io_in[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(io_in[3]),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input5 (.A(io_in[4]),
    .X(net5));
 sky130_fd_sc_hd__buf_2 input6 (.A(io_in[5]),
    .X(net6));
 sky130_fd_sc_hd__buf_6 input7 (.A(io_in[6]),
    .X(net7));
 sky130_fd_sc_hd__buf_2 input8 (.A(io_in[7]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_4 input9 (.A(io_in[8]),
    .X(net9));
 sky130_fd_sc_hd__buf_6 input10 (.A(rst),
    .X(net10));
 sky130_fd_sc_hd__buf_4 output11 (.A(net11),
    .X(io_oeb));
 sky130_fd_sc_hd__buf_4 output12 (.A(net12),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_4 output13 (.A(net13),
    .X(io_out[10]));
 sky130_fd_sc_hd__buf_4 output14 (.A(net14),
    .X(io_out[11]));
 sky130_fd_sc_hd__buf_4 output15 (.A(net15),
    .X(io_out[12]));
 sky130_fd_sc_hd__buf_4 output16 (.A(net16),
    .X(io_out[13]));
 sky130_fd_sc_hd__buf_4 output17 (.A(net17),
    .X(io_out[14]));
 sky130_fd_sc_hd__buf_4 output18 (.A(net18),
    .X(io_out[15]));
 sky130_fd_sc_hd__buf_4 output19 (.A(net19),
    .X(io_out[16]));
 sky130_fd_sc_hd__buf_4 output20 (.A(net20),
    .X(io_out[17]));
 sky130_fd_sc_hd__buf_4 output21 (.A(net21),
    .X(io_out[18]));
 sky130_fd_sc_hd__buf_4 output22 (.A(net22),
    .X(io_out[19]));
 sky130_fd_sc_hd__buf_4 output23 (.A(net23),
    .X(io_out[1]));
 sky130_fd_sc_hd__buf_4 output24 (.A(net24),
    .X(io_out[20]));
 sky130_fd_sc_hd__buf_4 output25 (.A(net25),
    .X(io_out[21]));
 sky130_fd_sc_hd__buf_4 output26 (.A(net26),
    .X(io_out[22]));
 sky130_fd_sc_hd__buf_4 output27 (.A(net27),
    .X(io_out[23]));
 sky130_fd_sc_hd__buf_4 output28 (.A(net28),
    .X(io_out[24]));
 sky130_fd_sc_hd__buf_4 output29 (.A(net29),
    .X(io_out[25]));
 sky130_fd_sc_hd__buf_4 output30 (.A(net30),
    .X(io_out[26]));
 sky130_fd_sc_hd__buf_4 output31 (.A(net31),
    .X(io_out[2]));
 sky130_fd_sc_hd__buf_4 output32 (.A(net32),
    .X(io_out[3]));
 sky130_fd_sc_hd__buf_4 output33 (.A(net33),
    .X(io_out[4]));
 sky130_fd_sc_hd__buf_4 output34 (.A(net34),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_4 output35 (.A(net35),
    .X(io_out[6]));
 sky130_fd_sc_hd__buf_4 output36 (.A(net36),
    .X(io_out[7]));
 sky130_fd_sc_hd__buf_4 output37 (.A(net37),
    .X(io_out[8]));
 sky130_fd_sc_hd__buf_4 output38 (.A(net38),
    .X(io_out[9]));
 sky130_fd_sc_hd__buf_4 fanout39 (.A(_1326_),
    .X(net39));
 sky130_fd_sc_hd__buf_2 fanout40 (.A(_1326_),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_8 fanout41 (.A(_2408_),
    .X(net41));
 sky130_fd_sc_hd__buf_4 fanout42 (.A(_1325_),
    .X(net42));
 sky130_fd_sc_hd__buf_4 fanout43 (.A(_0876_),
    .X(net43));
 sky130_fd_sc_hd__buf_4 fanout44 (.A(net45),
    .X(net44));
 sky130_fd_sc_hd__buf_4 fanout45 (.A(net46),
    .X(net45));
 sky130_fd_sc_hd__buf_4 fanout46 (.A(_1929_),
    .X(net46));
 sky130_fd_sc_hd__buf_12 max_cap47 (.A(_2623_),
    .X(net47));
 sky130_fd_sc_hd__buf_8 fanout48 (.A(net49),
    .X(net48));
 sky130_fd_sc_hd__buf_8 fanout49 (.A(_2581_),
    .X(net49));
 sky130_fd_sc_hd__buf_6 fanout50 (.A(_1333_),
    .X(net50));
 sky130_fd_sc_hd__buf_6 fanout51 (.A(net52),
    .X(net51));
 sky130_fd_sc_hd__buf_4 fanout52 (.A(_0724_),
    .X(net52));
 sky130_fd_sc_hd__buf_8 fanout53 (.A(_0693_),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_4 fanout54 (.A(_0693_),
    .X(net54));
 sky130_fd_sc_hd__buf_6 fanout55 (.A(net56),
    .X(net55));
 sky130_fd_sc_hd__buf_6 fanout56 (.A(_0632_),
    .X(net56));
 sky130_fd_sc_hd__buf_6 fanout57 (.A(_1310_),
    .X(net57));
 sky130_fd_sc_hd__buf_4 fanout58 (.A(net59),
    .X(net58));
 sky130_fd_sc_hd__buf_4 fanout59 (.A(_1309_),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_8 fanout60 (.A(net61),
    .X(net60));
 sky130_fd_sc_hd__buf_4 fanout61 (.A(_0726_),
    .X(net61));
 sky130_fd_sc_hd__buf_6 fanout62 (.A(_0722_),
    .X(net62));
 sky130_fd_sc_hd__buf_4 fanout63 (.A(_0718_),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_8 fanout64 (.A(net65),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_4 fanout65 (.A(_0650_),
    .X(net65));
 sky130_fd_sc_hd__buf_8 fanout66 (.A(_2778_),
    .X(net66));
 sky130_fd_sc_hd__buf_2 fanout67 (.A(_2778_),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_4 fanout68 (.A(net70),
    .X(net68));
 sky130_fd_sc_hd__buf_2 fanout69 (.A(net70),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_4 fanout70 (.A(_2777_),
    .X(net70));
 sky130_fd_sc_hd__buf_6 max_cap71 (.A(_2749_),
    .X(net71));
 sky130_fd_sc_hd__buf_8 fanout72 (.A(net73),
    .X(net72));
 sky130_fd_sc_hd__buf_6 fanout73 (.A(_2672_),
    .X(net73));
 sky130_fd_sc_hd__buf_8 fanout74 (.A(_2671_),
    .X(net74));
 sky130_fd_sc_hd__buf_6 fanout75 (.A(_2604_),
    .X(net75));
 sky130_fd_sc_hd__buf_6 fanout76 (.A(net77),
    .X(net76));
 sky130_fd_sc_hd__buf_6 fanout77 (.A(net78),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_8 fanout78 (.A(_2569_),
    .X(net78));
 sky130_fd_sc_hd__buf_6 fanout79 (.A(net82),
    .X(net79));
 sky130_fd_sc_hd__buf_4 fanout80 (.A(net82),
    .X(net80));
 sky130_fd_sc_hd__buf_6 fanout81 (.A(net82),
    .X(net81));
 sky130_fd_sc_hd__buf_4 fanout82 (.A(_2569_),
    .X(net82));
 sky130_fd_sc_hd__buf_6 fanout83 (.A(net84),
    .X(net83));
 sky130_fd_sc_hd__buf_6 fanout84 (.A(_1336_),
    .X(net84));
 sky130_fd_sc_hd__buf_6 fanout85 (.A(_0703_),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_8 fanout86 (.A(_0702_),
    .X(net86));
 sky130_fd_sc_hd__buf_4 fanout87 (.A(_0702_),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_16 fanout88 (.A(_0699_),
    .X(net88));
 sky130_fd_sc_hd__buf_8 fanout89 (.A(_0698_),
    .X(net89));
 sky130_fd_sc_hd__buf_4 fanout90 (.A(_0698_),
    .X(net90));
 sky130_fd_sc_hd__buf_4 fanout91 (.A(_0682_),
    .X(net91));
 sky130_fd_sc_hd__buf_8 fanout92 (.A(_0637_),
    .X(net92));
 sky130_fd_sc_hd__buf_12 fanout93 (.A(net95),
    .X(net93));
 sky130_fd_sc_hd__buf_4 fanout94 (.A(net95),
    .X(net94));
 sky130_fd_sc_hd__buf_8 fanout95 (.A(_0385_),
    .X(net95));
 sky130_fd_sc_hd__buf_8 fanout96 (.A(_0328_),
    .X(net96));
 sky130_fd_sc_hd__buf_4 fanout97 (.A(_0328_),
    .X(net97));
 sky130_fd_sc_hd__buf_12 fanout98 (.A(net100),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_4 fanout99 (.A(net100),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_8 fanout100 (.A(net101),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_8 fanout101 (.A(_2921_),
    .X(net101));
 sky130_fd_sc_hd__buf_12 fanout102 (.A(_2874_),
    .X(net102));
 sky130_fd_sc_hd__buf_8 fanout103 (.A(_2874_),
    .X(net103));
 sky130_fd_sc_hd__buf_6 fanout104 (.A(net105),
    .X(net104));
 sky130_fd_sc_hd__buf_6 fanout105 (.A(net106),
    .X(net105));
 sky130_fd_sc_hd__buf_4 fanout106 (.A(_2826_),
    .X(net106));
 sky130_fd_sc_hd__buf_12 fanout107 (.A(_2800_),
    .X(net107));
 sky130_fd_sc_hd__buf_4 fanout108 (.A(_2800_),
    .X(net108));
 sky130_fd_sc_hd__buf_6 fanout109 (.A(net110),
    .X(net109));
 sky130_fd_sc_hd__buf_12 fanout110 (.A(_2725_),
    .X(net110));
 sky130_fd_sc_hd__buf_6 fanout111 (.A(net112),
    .X(net111));
 sky130_fd_sc_hd__buf_12 fanout112 (.A(_2718_),
    .X(net112));
 sky130_fd_sc_hd__buf_12 fanout113 (.A(_2708_),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_4 fanout114 (.A(_2708_),
    .X(net114));
 sky130_fd_sc_hd__buf_6 fanout115 (.A(_2680_),
    .X(net115));
 sky130_fd_sc_hd__buf_6 fanout116 (.A(_2626_),
    .X(net116));
 sky130_fd_sc_hd__buf_6 fanout117 (.A(_2613_),
    .X(net117));
 sky130_fd_sc_hd__buf_6 fanout118 (.A(_2613_),
    .X(net118));
 sky130_fd_sc_hd__buf_6 fanout119 (.A(_2602_),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_16 fanout120 (.A(_2601_),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_4 fanout121 (.A(_2601_),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_8 fanout122 (.A(net123),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_8 fanout123 (.A(net124),
    .X(net123));
 sky130_fd_sc_hd__buf_4 fanout124 (.A(net125),
    .X(net124));
 sky130_fd_sc_hd__buf_6 fanout125 (.A(_2597_),
    .X(net125));
 sky130_fd_sc_hd__buf_6 fanout126 (.A(_2597_),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_8 fanout127 (.A(net128),
    .X(net127));
 sky130_fd_sc_hd__buf_8 fanout128 (.A(net130),
    .X(net128));
 sky130_fd_sc_hd__buf_6 fanout129 (.A(net130),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_8 fanout130 (.A(_2596_),
    .X(net130));
 sky130_fd_sc_hd__buf_4 fanout131 (.A(_2596_),
    .X(net131));
 sky130_fd_sc_hd__buf_4 fanout132 (.A(_2596_),
    .X(net132));
 sky130_fd_sc_hd__buf_6 fanout133 (.A(net134),
    .X(net133));
 sky130_fd_sc_hd__buf_6 fanout134 (.A(_2592_),
    .X(net134));
 sky130_fd_sc_hd__buf_6 fanout135 (.A(net136),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_8 fanout136 (.A(_2591_),
    .X(net136));
 sky130_fd_sc_hd__buf_6 fanout137 (.A(_2589_),
    .X(net137));
 sky130_fd_sc_hd__buf_6 fanout138 (.A(net139),
    .X(net138));
 sky130_fd_sc_hd__buf_6 fanout139 (.A(net140),
    .X(net139));
 sky130_fd_sc_hd__buf_8 fanout140 (.A(_2570_),
    .X(net140));
 sky130_fd_sc_hd__buf_6 fanout141 (.A(_2570_),
    .X(net141));
 sky130_fd_sc_hd__buf_2 fanout142 (.A(_2570_),
    .X(net142));
 sky130_fd_sc_hd__buf_6 fanout143 (.A(net147),
    .X(net143));
 sky130_fd_sc_hd__buf_8 fanout144 (.A(net146),
    .X(net144));
 sky130_fd_sc_hd__buf_2 fanout145 (.A(net146),
    .X(net145));
 sky130_fd_sc_hd__buf_6 fanout146 (.A(net147),
    .X(net146));
 sky130_fd_sc_hd__buf_4 fanout147 (.A(_2570_),
    .X(net147));
 sky130_fd_sc_hd__buf_6 fanout148 (.A(_2568_),
    .X(net148));
 sky130_fd_sc_hd__buf_8 fanout149 (.A(_2567_),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_4 fanout150 (.A(_2567_),
    .X(net150));
 sky130_fd_sc_hd__buf_8 fanout151 (.A(_0639_),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_4 fanout152 (.A(_0639_),
    .X(net152));
 sky130_fd_sc_hd__buf_4 fanout153 (.A(_0638_),
    .X(net153));
 sky130_fd_sc_hd__buf_6 fanout154 (.A(_0520_),
    .X(net154));
 sky130_fd_sc_hd__buf_6 fanout155 (.A(net157),
    .X(net155));
 sky130_fd_sc_hd__buf_2 fanout156 (.A(net157),
    .X(net156));
 sky130_fd_sc_hd__buf_6 fanout157 (.A(_2795_),
    .X(net157));
 sky130_fd_sc_hd__buf_6 fanout158 (.A(_2792_),
    .X(net158));
 sky130_fd_sc_hd__buf_8 fanout159 (.A(_2769_),
    .X(net159));
 sky130_fd_sc_hd__buf_4 fanout160 (.A(_2661_),
    .X(net160));
 sky130_fd_sc_hd__buf_6 wire161 (.A(_2609_),
    .X(net161));
 sky130_fd_sc_hd__buf_6 fanout162 (.A(_2587_),
    .X(net162));
 sky130_fd_sc_hd__buf_8 fanout163 (.A(_2566_),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_16 fanout164 (.A(_2565_),
    .X(net164));
 sky130_fd_sc_hd__buf_12 fanout165 (.A(_2564_),
    .X(net165));
 sky130_fd_sc_hd__buf_6 fanout166 (.A(net168),
    .X(net166));
 sky130_fd_sc_hd__buf_2 fanout167 (.A(net168),
    .X(net167));
 sky130_fd_sc_hd__buf_6 fanout168 (.A(_2558_),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_8 fanout169 (.A(net170),
    .X(net169));
 sky130_fd_sc_hd__buf_6 fanout170 (.A(_2797_),
    .X(net170));
 sky130_fd_sc_hd__buf_6 fanout171 (.A(_2791_),
    .X(net171));
 sky130_fd_sc_hd__buf_6 fanout172 (.A(net173),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_4 fanout173 (.A(_2790_),
    .X(net173));
 sky130_fd_sc_hd__buf_4 fanout174 (.A(net175),
    .X(net174));
 sky130_fd_sc_hd__buf_4 fanout175 (.A(_2722_),
    .X(net175));
 sky130_fd_sc_hd__buf_4 fanout176 (.A(_2686_),
    .X(net176));
 sky130_fd_sc_hd__buf_8 fanout177 (.A(_2644_),
    .X(net177));
 sky130_fd_sc_hd__buf_4 fanout178 (.A(_2644_),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_8 fanout179 (.A(net180),
    .X(net179));
 sky130_fd_sc_hd__buf_8 fanout180 (.A(_2642_),
    .X(net180));
 sky130_fd_sc_hd__buf_6 fanout181 (.A(net182),
    .X(net181));
 sky130_fd_sc_hd__buf_12 fanout182 (.A(_2640_),
    .X(net182));
 sky130_fd_sc_hd__buf_4 fanout183 (.A(_2638_),
    .X(net183));
 sky130_fd_sc_hd__buf_4 fanout184 (.A(_2638_),
    .X(net184));
 sky130_fd_sc_hd__buf_6 fanout185 (.A(_2636_),
    .X(net185));
 sky130_fd_sc_hd__buf_2 fanout186 (.A(_2636_),
    .X(net186));
 sky130_fd_sc_hd__buf_4 fanout187 (.A(net188),
    .X(net187));
 sky130_fd_sc_hd__buf_4 fanout188 (.A(_2634_),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_4 fanout189 (.A(net190),
    .X(net189));
 sky130_fd_sc_hd__buf_6 fanout190 (.A(_2632_),
    .X(net190));
 sky130_fd_sc_hd__buf_6 fanout191 (.A(net192),
    .X(net191));
 sky130_fd_sc_hd__buf_6 fanout192 (.A(_2624_),
    .X(net192));
 sky130_fd_sc_hd__buf_6 fanout193 (.A(_2588_),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_4 fanout194 (.A(_2588_),
    .X(net194));
 sky130_fd_sc_hd__buf_8 fanout195 (.A(_2585_),
    .X(net195));
 sky130_fd_sc_hd__buf_8 fanout196 (.A(_2583_),
    .X(net196));
 sky130_fd_sc_hd__buf_6 fanout197 (.A(_2576_),
    .X(net197));
 sky130_fd_sc_hd__buf_2 fanout198 (.A(_2576_),
    .X(net198));
 sky130_fd_sc_hd__buf_8 fanout199 (.A(net200),
    .X(net199));
 sky130_fd_sc_hd__buf_6 fanout200 (.A(net201),
    .X(net200));
 sky130_fd_sc_hd__buf_8 fanout201 (.A(_2575_),
    .X(net201));
 sky130_fd_sc_hd__buf_12 fanout202 (.A(net205),
    .X(net202));
 sky130_fd_sc_hd__buf_8 fanout203 (.A(net205),
    .X(net203));
 sky130_fd_sc_hd__buf_12 fanout204 (.A(net205),
    .X(net204));
 sky130_fd_sc_hd__buf_6 fanout205 (.A(_2546_),
    .X(net205));
 sky130_fd_sc_hd__buf_12 fanout206 (.A(net207),
    .X(net206));
 sky130_fd_sc_hd__buf_12 fanout207 (.A(_2545_),
    .X(net207));
 sky130_fd_sc_hd__buf_12 fanout208 (.A(_2544_),
    .X(net208));
 sky130_fd_sc_hd__buf_6 fanout209 (.A(_2544_),
    .X(net209));
 sky130_fd_sc_hd__buf_8 fanout210 (.A(net212),
    .X(net210));
 sky130_fd_sc_hd__buf_4 fanout211 (.A(net212),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_16 fanout212 (.A(\as2650.psl[4] ),
    .X(net212));
 sky130_fd_sc_hd__buf_6 fanout213 (.A(\as2650.psl[4] ),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_4 fanout214 (.A(\as2650.psl[4] ),
    .X(net214));
 sky130_fd_sc_hd__buf_8 fanout215 (.A(net216),
    .X(net215));
 sky130_fd_sc_hd__buf_12 fanout216 (.A(\as2650.psu[0] ),
    .X(net216));
 sky130_fd_sc_hd__buf_8 fanout217 (.A(net218),
    .X(net217));
 sky130_fd_sc_hd__buf_12 fanout218 (.A(\as2650.psu[1] ),
    .X(net218));
 sky130_fd_sc_hd__buf_6 fanout219 (.A(net220),
    .X(net219));
 sky130_fd_sc_hd__buf_8 fanout220 (.A(net221),
    .X(net220));
 sky130_fd_sc_hd__buf_4 fanout221 (.A(\as2650.psu[2] ),
    .X(net221));
 sky130_fd_sc_hd__buf_4 fanout222 (.A(net224),
    .X(net222));
 sky130_fd_sc_hd__buf_6 fanout223 (.A(net224),
    .X(net223));
 sky130_fd_sc_hd__buf_8 fanout224 (.A(net225),
    .X(net224));
 sky130_fd_sc_hd__buf_6 fanout225 (.A(net228),
    .X(net225));
 sky130_fd_sc_hd__buf_8 fanout226 (.A(net228),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_4 fanout227 (.A(net228),
    .X(net227));
 sky130_fd_sc_hd__buf_6 fanout228 (.A(\as2650.ins_reg[4] ),
    .X(net228));
 sky130_fd_sc_hd__buf_6 fanout229 (.A(\as2650.ins_reg[3] ),
    .X(net229));
 sky130_fd_sc_hd__buf_6 fanout230 (.A(net231),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_16 fanout231 (.A(\as2650.ins_reg[3] ),
    .X(net231));
 sky130_fd_sc_hd__buf_8 fanout232 (.A(net235),
    .X(net232));
 sky130_fd_sc_hd__buf_6 fanout233 (.A(net234),
    .X(net233));
 sky130_fd_sc_hd__buf_8 fanout234 (.A(net235),
    .X(net234));
 sky130_fd_sc_hd__buf_6 fanout235 (.A(\as2650.r0[7] ),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_8 fanout236 (.A(net237),
    .X(net236));
 sky130_fd_sc_hd__buf_6 fanout237 (.A(net239),
    .X(net237));
 sky130_fd_sc_hd__buf_12 fanout238 (.A(net239),
    .X(net238));
 sky130_fd_sc_hd__buf_8 fanout239 (.A(\as2650.r0[6] ),
    .X(net239));
 sky130_fd_sc_hd__buf_6 fanout240 (.A(\as2650.r0[5] ),
    .X(net240));
 sky130_fd_sc_hd__buf_6 fanout241 (.A(net242),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_16 fanout242 (.A(\as2650.r0[5] ),
    .X(net242));
 sky130_fd_sc_hd__buf_6 fanout243 (.A(\as2650.r0[4] ),
    .X(net243));
 sky130_fd_sc_hd__buf_4 fanout244 (.A(\as2650.r0[4] ),
    .X(net244));
 sky130_fd_sc_hd__buf_8 fanout245 (.A(\as2650.r0[4] ),
    .X(net245));
 sky130_fd_sc_hd__buf_12 fanout246 (.A(net249),
    .X(net246));
 sky130_fd_sc_hd__buf_6 fanout247 (.A(net248),
    .X(net247));
 sky130_fd_sc_hd__buf_8 fanout248 (.A(net249),
    .X(net248));
 sky130_fd_sc_hd__buf_8 fanout249 (.A(\as2650.r0[3] ),
    .X(net249));
 sky130_fd_sc_hd__buf_6 fanout250 (.A(\as2650.r0[2] ),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_8 fanout251 (.A(\as2650.r0[2] ),
    .X(net251));
 sky130_fd_sc_hd__buf_6 fanout252 (.A(net253),
    .X(net252));
 sky130_fd_sc_hd__buf_6 fanout253 (.A(\as2650.r0[2] ),
    .X(net253));
 sky130_fd_sc_hd__buf_6 fanout254 (.A(\as2650.r0[1] ),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_8 fanout255 (.A(\as2650.r0[1] ),
    .X(net255));
 sky130_fd_sc_hd__buf_4 fanout256 (.A(net257),
    .X(net256));
 sky130_fd_sc_hd__buf_2 fanout257 (.A(net258),
    .X(net257));
 sky130_fd_sc_hd__buf_6 fanout258 (.A(\as2650.r0[1] ),
    .X(net258));
 sky130_fd_sc_hd__buf_6 fanout259 (.A(net263),
    .X(net259));
 sky130_fd_sc_hd__buf_4 fanout260 (.A(net261),
    .X(net260));
 sky130_fd_sc_hd__buf_6 fanout261 (.A(net262),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_8 fanout262 (.A(net263),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_16 fanout263 (.A(\as2650.r0[0] ),
    .X(net263));
 sky130_fd_sc_hd__buf_8 fanout264 (.A(\as2650.pc[12] ),
    .X(net264));
 sky130_fd_sc_hd__buf_8 fanout265 (.A(\as2650.pc[11] ),
    .X(net265));
 sky130_fd_sc_hd__buf_8 fanout266 (.A(\as2650.pc[10] ),
    .X(net266));
 sky130_fd_sc_hd__buf_8 fanout267 (.A(\as2650.pc[9] ),
    .X(net267));
 sky130_fd_sc_hd__buf_4 fanout268 (.A(\as2650.pc[8] ),
    .X(net268));
 sky130_fd_sc_hd__buf_8 fanout269 (.A(\as2650.pc[7] ),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_8 fanout270 (.A(\as2650.pc[7] ),
    .X(net270));
 sky130_fd_sc_hd__buf_4 fanout271 (.A(net272),
    .X(net271));
 sky130_fd_sc_hd__buf_6 fanout272 (.A(\as2650.pc[6] ),
    .X(net272));
 sky130_fd_sc_hd__buf_4 fanout273 (.A(\as2650.pc[5] ),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_4 fanout274 (.A(\as2650.pc[5] ),
    .X(net274));
 sky130_fd_sc_hd__buf_6 fanout275 (.A(\as2650.pc[4] ),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_8 fanout276 (.A(\as2650.pc[4] ),
    .X(net276));
 sky130_fd_sc_hd__buf_4 fanout277 (.A(net278),
    .X(net277));
 sky130_fd_sc_hd__buf_4 fanout278 (.A(\as2650.pc[3] ),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_8 fanout279 (.A(net280),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_4 fanout280 (.A(net281),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_4 fanout281 (.A(\as2650.pc[2] ),
    .X(net281));
 sky130_fd_sc_hd__buf_4 fanout282 (.A(net284),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_2 fanout283 (.A(net284),
    .X(net283));
 sky130_fd_sc_hd__buf_6 fanout284 (.A(\as2650.pc[1] ),
    .X(net284));
 sky130_fd_sc_hd__buf_4 fanout285 (.A(net286),
    .X(net285));
 sky130_fd_sc_hd__buf_4 fanout286 (.A(net287),
    .X(net286));
 sky130_fd_sc_hd__buf_6 fanout287 (.A(\as2650.pc[0] ),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_8 fanout288 (.A(\as2650.cycle[3] ),
    .X(net288));
 sky130_fd_sc_hd__buf_6 fanout289 (.A(\as2650.cycle[2] ),
    .X(net289));
 sky130_fd_sc_hd__buf_6 fanout290 (.A(net291),
    .X(net290));
 sky130_fd_sc_hd__buf_8 fanout291 (.A(\as2650.cycle[0] ),
    .X(net291));
 sky130_fd_sc_hd__buf_6 fanout292 (.A(net293),
    .X(net292));
 sky130_fd_sc_hd__buf_12 fanout293 (.A(\as2650.halted ),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_16 fanout294 (.A(\as2650.addr_buff[7] ),
    .X(net294));
 sky130_fd_sc_hd__buf_6 fanout295 (.A(\as2650.addr_buff[1] ),
    .X(net295));
 sky130_fd_sc_hd__buf_6 fanout296 (.A(\as2650.addr_buff[0] ),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_16 fanout297 (.A(net298),
    .X(net297));
 sky130_fd_sc_hd__buf_12 fanout298 (.A(\as2650.ins_reg[7] ),
    .X(net298));
 sky130_fd_sc_hd__buf_12 fanout299 (.A(\as2650.ins_reg[6] ),
    .X(net299));
 sky130_fd_sc_hd__buf_6 fanout300 (.A(net301),
    .X(net300));
 sky130_fd_sc_hd__buf_12 fanout301 (.A(\as2650.ins_reg[5] ),
    .X(net301));
 sky130_fd_sc_hd__buf_8 fanout302 (.A(\as2650.ins_reg[2] ),
    .X(net302));
 sky130_fd_sc_hd__buf_8 fanout303 (.A(\as2650.ins_reg[2] ),
    .X(net303));
 sky130_fd_sc_hd__buf_6 fanout304 (.A(\as2650.ins_reg[1] ),
    .X(net304));
 sky130_fd_sc_hd__buf_8 fanout305 (.A(\as2650.ins_reg[1] ),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_16 fanout306 (.A(net307),
    .X(net306));
 sky130_fd_sc_hd__buf_12 fanout307 (.A(\as2650.ins_reg[0] ),
    .X(net307));
 sky130_fd_sc_hd__buf_4 fanout308 (.A(\as2650.ins_reg[0] ),
    .X(net308));
 sky130_fd_sc_hd__buf_6 fanout309 (.A(net311),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_4 fanout310 (.A(net311),
    .X(net310));
 sky130_fd_sc_hd__buf_4 fanout311 (.A(net312),
    .X(net311));
 sky130_fd_sc_hd__buf_6 fanout312 (.A(_2548_),
    .X(net312));
 sky130_fd_sc_hd__buf_4 fanout313 (.A(net314),
    .X(net313));
 sky130_fd_sc_hd__buf_4 fanout314 (.A(net315),
    .X(net314));
 sky130_fd_sc_hd__buf_6 fanout315 (.A(net321),
    .X(net315));
 sky130_fd_sc_hd__buf_4 fanout316 (.A(net318),
    .X(net316));
 sky130_fd_sc_hd__buf_2 fanout317 (.A(net318),
    .X(net317));
 sky130_fd_sc_hd__buf_4 fanout318 (.A(net321),
    .X(net318));
 sky130_fd_sc_hd__buf_6 fanout319 (.A(net321),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_4 fanout320 (.A(net321),
    .X(net320));
 sky130_fd_sc_hd__buf_6 fanout321 (.A(_2547_),
    .X(net321));
 sky130_fd_sc_hd__buf_4 fanout322 (.A(net323),
    .X(net322));
 sky130_fd_sc_hd__buf_2 fanout323 (.A(net324),
    .X(net323));
 sky130_fd_sc_hd__buf_6 fanout324 (.A(net325),
    .X(net324));
 sky130_fd_sc_hd__buf_8 fanout325 (.A(net327),
    .X(net325));
 sky130_fd_sc_hd__buf_6 fanout326 (.A(net327),
    .X(net326));
 sky130_fd_sc_hd__buf_8 fanout327 (.A(net8),
    .X(net327));
 sky130_fd_sc_hd__buf_8 fanout328 (.A(net330),
    .X(net328));
 sky130_fd_sc_hd__buf_6 fanout329 (.A(net330),
    .X(net329));
 sky130_fd_sc_hd__buf_8 fanout330 (.A(net7),
    .X(net330));
 sky130_fd_sc_hd__buf_8 fanout331 (.A(net7),
    .X(net331));
 sky130_fd_sc_hd__buf_6 fanout332 (.A(net334),
    .X(net332));
 sky130_fd_sc_hd__clkbuf_4 fanout333 (.A(net334),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_16 fanout334 (.A(net6),
    .X(net334));
 sky130_fd_sc_hd__clkbuf_16 fanout335 (.A(net337),
    .X(net335));
 sky130_fd_sc_hd__clkbuf_2 fanout336 (.A(net337),
    .X(net336));
 sky130_fd_sc_hd__buf_12 fanout337 (.A(net5),
    .X(net337));
 sky130_fd_sc_hd__buf_6 fanout338 (.A(net340),
    .X(net338));
 sky130_fd_sc_hd__buf_8 fanout339 (.A(net340),
    .X(net339));
 sky130_fd_sc_hd__buf_8 fanout340 (.A(net4),
    .X(net340));
 sky130_fd_sc_hd__buf_8 fanout341 (.A(net343),
    .X(net341));
 sky130_fd_sc_hd__buf_4 fanout342 (.A(net343),
    .X(net342));
 sky130_fd_sc_hd__buf_12 fanout343 (.A(net3),
    .X(net343));
 sky130_fd_sc_hd__buf_8 fanout344 (.A(net346),
    .X(net344));
 sky130_fd_sc_hd__buf_6 fanout345 (.A(net346),
    .X(net345));
 sky130_fd_sc_hd__buf_8 fanout346 (.A(net2),
    .X(net346));
 sky130_fd_sc_hd__buf_12 fanout347 (.A(net10),
    .X(net347));
 sky130_fd_sc_hd__buf_6 fanout348 (.A(net10),
    .X(net348));
 sky130_fd_sc_hd__clkbuf_16 fanout349 (.A(net1),
    .X(net349));
 sky130_fd_sc_hd__buf_8 fanout350 (.A(net1),
    .X(net350));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__5595__A2 (.DIODE(_0288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4653__B (.DIODE(_0288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4652__B (.DIODE(_0288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3690__A1 (.DIODE(_0288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3358__B1 (.DIODE(_0288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5803__A2 (.DIODE(_0309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5801__A2 (.DIODE(_0309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__A2 (.DIODE(_0309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3897__D (.DIODE(_0309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3691__A0 (.DIODE(_0309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3379__A1 (.DIODE(_0309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5731__A1 (.DIODE(_0310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5713__A1 (.DIODE(_0310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3380__A2 (.DIODE(_0310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5504__A1 (.DIODE(_0317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3693__A (.DIODE(_0317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3388__B (.DIODE(_0317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__A2 (.DIODE(_0321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4537__A (.DIODE(_0321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3695__A (.DIODE(_0321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3392__B (.DIODE(_0321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__B (.DIODE(_0327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__B (.DIODE(_0327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3398__B1 (.DIODE(_0327_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout97_A (.DIODE(_0328_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout96_A (.DIODE(_0328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5639__A (.DIODE(_0329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5631__A1 (.DIODE(_0329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3479__A1 (.DIODE(_0329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3470__B (.DIODE(_0329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3463__A (.DIODE(_0329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3451__A2 (.DIODE(_0329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5608__A2 (.DIODE(_0337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__B (.DIODE(_0337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4710__B (.DIODE(_0337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3700__A (.DIODE(_0337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3408__A1 (.DIODE(_0337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__B (.DIODE(_0340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3412__A1 (.DIODE(_0340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5607__B (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__B (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3702__A1 (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__A2 (.DIODE(_0360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5606__B (.DIODE(_0360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3431__A (.DIODE(_0360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5733__A1 (.DIODE(_0362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5715__A1 (.DIODE(_0362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3433__A2 (.DIODE(_0362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__A1 (.DIODE(_0370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3442__B (.DIODE(_0370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__A2 (.DIODE(_0374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3504__A (.DIODE(_0374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3464__A (.DIODE(_0374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3446__A (.DIODE(_0374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__A2 (.DIODE(_0381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4537__D_N (.DIODE(_0381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3705__A (.DIODE(_0381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3457__B (.DIODE(_0381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__B (.DIODE(_0382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5352__B (.DIODE(_0382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3455__A2 (.DIODE(_0382_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout95_A (.DIODE(_0385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5620__A0 (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4739__B (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__B (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__A1 (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3468__A1 (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5620__A1 (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4732__B (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4731__B (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3711__A1 (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3469__A0 (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5805__A2 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5804__B2 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5622__A2 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3898__B (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3712__A0 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3486__A1 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5735__A1 (.DIODE(_0415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__A1 (.DIODE(_0415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3487__A2 (.DIODE(_0415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__A1 (.DIODE(_0422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3495__B (.DIODE(_0422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5633__A0 (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4811__A2 (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4787__B (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3720__A1 (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3509__A2 (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5633__A1 (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__B (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__B (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3721__A1 (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3512__A2 (.DIODE(_0439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5807__A2 (.DIODE(_0458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5805__B2 (.DIODE(_0458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5635__A2 (.DIODE(_0458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3898__C (.DIODE(_0458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3722__A1 (.DIODE(_0458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3531__A2 (.DIODE(_0458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5736__A1 (.DIODE(_0459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5719__A1 (.DIODE(_0459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3532__A2 (.DIODE(_0459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5646__A0 (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__A2 (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__B (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__B (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__A1 (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3548__A1 (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5646__A1 (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__B (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4805__B (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4804__B (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3730__A1 (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3551__A1 (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5807__B1 (.DIODE(_0494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5806__A (.DIODE(_0494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5797__A (.DIODE(_0494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5648__A2 (.DIODE(_0494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__B (.DIODE(_0494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3731__A0 (.DIODE(_0494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3568__A1 (.DIODE(_0494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5738__A1 (.DIODE(_0495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__A1 (.DIODE(_0495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3569__A2 (.DIODE(_0495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4414__S (.DIODE(_0498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4412__S (.DIODE(_0498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4410__S (.DIODE(_0498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4408__S (.DIODE(_0498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__S (.DIODE(_0498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4404__S (.DIODE(_0498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4402__S (.DIODE(_0498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4400__S (.DIODE(_0498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__A (.DIODE(_0498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3581__S (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3580__S (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3579__S (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3578__S (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3577__S (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3576__S (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3575__S (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3597__S (.DIODE(_0501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3595__S (.DIODE(_0501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__S (.DIODE(_0501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3591__S (.DIODE(_0501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3589__S (.DIODE(_0501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3587__S (.DIODE(_0501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3585__S (.DIODE(_0501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3608__S (.DIODE(_0512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3607__S (.DIODE(_0512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3606__S (.DIODE(_0512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3605__S (.DIODE(_0512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3604__S (.DIODE(_0512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3603__S (.DIODE(_0512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3602__S (.DIODE(_0512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4025__B (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3654__B (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3653__B (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3652__B (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3648__B1 (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3611__B (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3650__A2 (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3624__B (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4246__A1 (.DIODE(_0547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4026__A1 (.DIODE(_0547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3657__A2 (.DIODE(_0547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4244__B (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4022__B (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3723__B2 (.DIODE(_0553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3714__B2 (.DIODE(_0553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3704__B2 (.DIODE(_0553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3692__B2 (.DIODE(_0553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3681__B2 (.DIODE(_0553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4024__B1 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3732__A3 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3715__A3 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3713__A3 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3694__A2 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3683__A2 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3671__A2 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3658__B1 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3655__C1 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4280__A1 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4031__A1 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3668__A2 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4313__A1 (.DIODE(_0582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4043__A1 (.DIODE(_0582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3681__B1 (.DIODE(_0582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4343__A1 (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4061__A1 (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3692__B1 (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__A1 (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4086__A1 (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3704__B1 (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4382__A1 (.DIODE(_0611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4115__A1 (.DIODE(_0611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3714__B1 (.DIODE(_0611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4392__A1 (.DIODE(_0620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4150__A1 (.DIODE(_0620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3723__B1 (.DIODE(_0620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4396__A1 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4192__A1 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3732__B1 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5792__A2 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5640__A1 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5639__B (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__A2 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5547__A2 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3981__A2_N (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3736__B (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5791__B1 (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__B2 (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5625__C1 (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5545__B1 (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__C1 (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__B2 (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3738__C (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3737__B (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5809__A2 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__A2 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5613__B1 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5601__A1 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__A1 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5577__A1 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5069__B (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3765__A (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__B1 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5762__A1 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5761__B (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5169__A2 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5071__A (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3837__B (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3830__B (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3763__B (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_A (.DIODE(_0638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__C (.DIODE(_0638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__C1 (.DIODE(_0638_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_A (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout151_A (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__A2 (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__D (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3928__A3 (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3927__C (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3778__B (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3748__B (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3746__A2 (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5836__A3 (.DIODE(_0644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3978__A3 (.DIODE(_0644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3750__A2 (.DIODE(_0644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4431__S (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4429__S (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4427__S (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4425__S (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4423__S (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4421__S (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4419__S (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4417__S (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3786__B1 (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3793__S (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__S (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__S (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__S (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3789__S (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3788__S (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__S (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__A1 (.DIODE(_0683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__A1 (.DIODE(_0683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__B (.DIODE(_0683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__B1 (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__B2 (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4850__A1 (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__B1 (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4659__C1 (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__A1 (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__C1 (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__A1 (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__A1 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4792__A1 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4744__A1 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__A1 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__B (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__A1 (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4721__B2 (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4636__A1 (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__A1 (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4568__B1 (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3815__B (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__B (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__A (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4745__A1 (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__A1 (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3832__B (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__D (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5019__B1 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__A1 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4862__B1 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4823__B1 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__C1 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4674__C1 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__B1 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4569__B2 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__C (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__B (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5559__B (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__A (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5169__A4 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5093__C1 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__B (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__B1 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5031__A1 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4534__A3 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__A1 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4519__A1 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4513__C (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__A1 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout88_A (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5111__A2 (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__A2 (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout87_A (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout86_A (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5749__C (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__B1 (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__C (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4516__A (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__B1 (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4007__A2 (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4000__B (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3826__A (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__A1 (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4496__B (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__A (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3998__A2 (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3843__B (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__B1 (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__A2_N (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__A3 (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__A3 (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4492__B2 (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3918__B (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__B1 (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__A2 (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5444__A2_N (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__A2_N (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5393__B2 (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__A1_N (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3833__C (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout63_A (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5786__B1 (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4499__B (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout62_A (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__B1 (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5603__A2 (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5778__A2 (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__A3 (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__B1 (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__A1_N (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5393__A1 (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3920__B (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3908__C (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__A1 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3870__S (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3867__S (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3864__S (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3861__S (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__S (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3855__S (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3852__S (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__S (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3852__A1 (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3855__A1 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__A1 (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3861__A1 (.DIODE(_0744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3864__A1 (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3867__A1 (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3870__A1 (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4448__S (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4446__S (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4444__S (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4442__S (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__S (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4438__S (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__S (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__S (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3874__A (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__S (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__S (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3879__S (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3878__S (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3877__S (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3876__S (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3875__S (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__B1 (.DIODE(_0793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5775__A2 (.DIODE(_0793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5755__B (.DIODE(_0793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4533__C (.DIODE(_0793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__B1 (.DIODE(_0793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3921__A (.DIODE(_0793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5778__B1 (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5766__A2 (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5754__A2 (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4534__A4 (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5786__C1 (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__A3 (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4492__A2 (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3937__A (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__D (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4991__A (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4541__A_N (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__B (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5061__B (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3937__B (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__S (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4484__S (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4482__S (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4480__S (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4478__S (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4476__S (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4474__S (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4472__S (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__B1 (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3996__S (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3995__S (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3994__S (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3993__S (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3992__S (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3991__S (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3990__S (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5692__S (.DIODE(_0869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5690__S (.DIODE(_0869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__S (.DIODE(_0869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__S (.DIODE(_0869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5684__S (.DIODE(_0869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__S (.DIODE(_0869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5680__S (.DIODE(_0869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5678__S (.DIODE(_0869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4012__B1 (.DIODE(_0869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4019__S (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4018__S (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__S (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4016__S (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4015__S (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4014__S (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4013__S (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4396__A2 (.DIODE(_1079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4392__A2 (.DIODE(_1079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4382__A2 (.DIODE(_1079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__A2 (.DIODE(_1079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4343__A2 (.DIODE(_1079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4313__A2 (.DIODE(_1079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4280__A2 (.DIODE(_1079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4246__A2 (.DIODE(_1079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4245__B (.DIODE(_1079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4413__S (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__S (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__S (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4407__S (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4405__S (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4403__S (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4401__S (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__S (.DIODE(_1234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4428__S (.DIODE(_1234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4426__S (.DIODE(_1234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4424__S (.DIODE(_1234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4422__S (.DIODE(_1234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4420__S (.DIODE(_1234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4418__S (.DIODE(_1234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__S (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__S (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4443__S (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4441__S (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4439__S (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__S (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4435__S (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__S (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5491__B1_N (.DIODE(_1255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__B1 (.DIODE(_1255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5454__A1 (.DIODE(_1255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__A1 (.DIODE(_1255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4455__B2 (.DIODE(_1255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4469__S (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__S (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4467__S (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__S (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4465__S (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4464__S (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4463__S (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__S (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4485__S (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4483__S (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4481__S (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4479__S (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4477__S (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4475__S (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4473__S (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4471__S (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__A2 (.DIODE(_1279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4493__C1 (.DIODE(_1279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4505__A2 (.DIODE(_1288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__B (.DIODE(_1288_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout57_A (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5505__A1 (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__A1 (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5214__A1 (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__A1 (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4938__A1 (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__A1 (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__A1 (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4764__A1 (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__A1 (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4687__A1 (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__A1 (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__A1 (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__A (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5151__S (.DIODE(_1322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__C (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5063__B (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__C (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__C1 (.DIODE(_1324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__A1 (.DIODE(_1324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4541__B (.DIODE(_1324_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout50_A (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5388__B2 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__A1 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__A (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__A1 (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__B2 (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__B2 (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5148__A2 (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4553__B (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4568__B2 (.DIODE(_1350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5561__B1 (.DIODE(_1362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__A2_N (.DIODE(_1362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__A2 (.DIODE(_1362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__B1 (.DIODE(_1362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4588__A2 (.DIODE(_1362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__A2 (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5175__A2 (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__A2 (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4933__A2 (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__B1 (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4769__B1 (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__B1 (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4688__B1 (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__A2 (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4603__A2 (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4636__A2 (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__A2 (.DIODE(_1448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4721__B1 (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4745__A2 (.DIODE(_1523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__A2 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__B1 (.DIODE(_1595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__A (.DIODE(_1617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4906__B (.DIODE(_1617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__B (.DIODE(_1617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__B (.DIODE(_1617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5490__C (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5489__A2 (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5464__A1 (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4964__B (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4940__B (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4908__B (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5465__A2 (.DIODE(_1736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4967__C1 (.DIODE(_1736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__B (.DIODE(_1736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__B1 (.DIODE(_1768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__A2 (.DIODE(_1768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__S (.DIODE(_1805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__S (.DIODE(_1805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5056__S (.DIODE(_1805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5054__S (.DIODE(_1805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5051__S (.DIODE(_1805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__S (.DIODE(_1805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5045__A2 (.DIODE(_1805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__B (.DIODE(_1805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5041__S (.DIODE(_1805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__B (.DIODE(_1822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5349__A1 (.DIODE(_1822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5268__A1 (.DIODE(_1822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__A1 (.DIODE(_1822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5512__A2 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5185__B (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5087__A2 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5067__B1 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__B1 (.DIODE(_1870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5120__B1 (.DIODE(_1870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__A2 (.DIODE(_1905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5546__A2 (.DIODE(_1915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__A2_N (.DIODE(_1915_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout46_A (.DIODE(_1929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5539__A1 (.DIODE(_1930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__A1 (.DIODE(_1930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5247__C1 (.DIODE(_1930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5182__C1 (.DIODE(_1930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__A1 (.DIODE(_1933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5477__A1 (.DIODE(_1933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5457__A1 (.DIODE(_1933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5386__B2 (.DIODE(_1933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5326__B2 (.DIODE(_1933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__B1 (.DIODE(_1933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__A2 (.DIODE(_1933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5528__A (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5499__C1 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5476__C1 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5456__A2 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5350__A1 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5296__A2 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5268__B2 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__B2 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__B1 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__A2 (.DIODE(_1957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__B1 (.DIODE(_1958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5211__A (.DIODE(_1958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__B2 (.DIODE(_1991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__B1 (.DIODE(_1991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__A2 (.DIODE(_2021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__B1 (.DIODE(_2022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__A (.DIODE(_2022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__A2 (.DIODE(_2036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5610__B (.DIODE(_2048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5304__A2 (.DIODE(_2048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5334__A2 (.DIODE(_2077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5624__B (.DIODE(_2078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__B1 (.DIODE(_2078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__B (.DIODE(_2108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__B1 (.DIODE(_2108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__A2 (.DIODE(_2131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5651__A2 (.DIODE(_2134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5393__B1 (.DIODE(_2134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__B1 (.DIODE(_2308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__B1 (.DIODE(_2319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5601__B1 (.DIODE(_2330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5693__B1 (.DIODE(_2383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5676__B (.DIODE(_2383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5658__B (.DIODE(_2383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5675__S (.DIODE(_2384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5673__S (.DIODE(_2384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5671__S (.DIODE(_2384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5669__S (.DIODE(_2384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5667__S (.DIODE(_2384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5665__S (.DIODE(_2384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5663__S (.DIODE(_2384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5661__S (.DIODE(_2384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5674__S (.DIODE(_2385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5672__S (.DIODE(_2385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5670__S (.DIODE(_2385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5668__S (.DIODE(_2385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__S (.DIODE(_2385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5664__S (.DIODE(_2385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5662__S (.DIODE(_2385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5660__S (.DIODE(_2385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5691__S (.DIODE(_2394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5689__S (.DIODE(_2394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5687__S (.DIODE(_2394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5685__S (.DIODE(_2394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5683__S (.DIODE(_2394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5681__S (.DIODE(_2394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5679__S (.DIODE(_2394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5677__S (.DIODE(_2394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__S (.DIODE(_2403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__S (.DIODE(_2403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5698__S (.DIODE(_2403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5697__S (.DIODE(_2403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5696__S (.DIODE(_2403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__S (.DIODE(_2403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5694__S (.DIODE(_2403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__A2 (.DIODE(_2405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5719__A2 (.DIODE(_2405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__A2 (.DIODE(_2405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5715__A2 (.DIODE(_2405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5713__A2 (.DIODE(_2405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5710__A2 (.DIODE(_2405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__A2 (.DIODE(_2405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5706__B1 (.DIODE(_2405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__A2 (.DIODE(_2405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5703__B (.DIODE(_2405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5738__A2 (.DIODE(_2418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5736__A2 (.DIODE(_2418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5735__A2 (.DIODE(_2418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5733__A2 (.DIODE(_2418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5731__A2 (.DIODE(_2418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5729__A2 (.DIODE(_2418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5727__A2 (.DIODE(_2418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5725__A2 (.DIODE(_2418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5724__B (.DIODE(_2418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3647__C1 (.DIODE(_2525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3644__A1 (.DIODE(_2525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3641__A (.DIODE(_2525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3621__A (.DIODE(_2525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3084__A (.DIODE(_2525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__A2 (.DIODE(_2535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5139__A1 (.DIODE(_2535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__A1 (.DIODE(_2535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__A (.DIODE(_2535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5125__A1 (.DIODE(_2535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__A1 (.DIODE(_2535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5111__A1 (.DIODE(_2535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5095__A1 (.DIODE(_2535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__A (.DIODE(_2535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4496__A (.DIODE(_2535_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_A (.DIODE(_2544_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_A (.DIODE(_2544_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout321_A (.DIODE(_2547_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout312_A (.DIODE(_2548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5766__A1 (.DIODE(_2550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__A (.DIODE(_2550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__A (.DIODE(_2550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3971__A2 (.DIODE(_2550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3965__A2 (.DIODE(_2550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3957__A1 (.DIODE(_2550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__B2 (.DIODE(_2552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__A (.DIODE(_2552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4660__A (.DIODE(_2552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3970__B1 (.DIODE(_2552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3962__A2 (.DIODE(_2552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3959__A1 (.DIODE(_2552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5615__A1 (.DIODE(_2553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__A (.DIODE(_2553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3972__B1 (.DIODE(_2553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3962__B1 (.DIODE(_2553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__A1 (.DIODE(_2553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__B2 (.DIODE(_2554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3969__B1 (.DIODE(_2554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3964__B1 (.DIODE(_2554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3959__B2 (.DIODE(_2554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5841__B2 (.DIODE(_2556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4787__A (.DIODE(_2556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4786__A0 (.DIODE(_2556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3971__B1 (.DIODE(_2556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3963__B1 (.DIODE(_2556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__B2 (.DIODE(_2556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3944__D (.DIODE(_2556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__A1 (.DIODE(_2557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__A (.DIODE(_2557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__A (.DIODE(_2557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3997__B (.DIODE(_2560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3609__B (.DIODE(_2560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3094__A (.DIODE(_2560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3091__B (.DIODE(_2560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3064__A (.DIODE(_2560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3041__B1 (.DIODE(_2560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3033__B1 (.DIODE(_2560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3028__B1 (.DIODE(_2560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2991__A (.DIODE(_2560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4459__A (.DIODE(_2561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3621__B (.DIODE(_2561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3228__B (.DIODE(_2561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3199__A (.DIODE(_2561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3164__B (.DIODE(_2561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3127__A (.DIODE(_2561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3108__A1 (.DIODE(_2561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3100__A (.DIODE(_2561_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout165_A (.DIODE(_2564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__B (.DIODE(_2564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__B (.DIODE(_2564_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout163_A (.DIODE(_2566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__C (.DIODE(_2566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__C (.DIODE(_2566_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_A (.DIODE(_2568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5745__B (.DIODE(_2568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__B1 (.DIODE(_2568_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_A (.DIODE(_2570_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_A (.DIODE(_2570_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_A (.DIODE(_2570_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_A (.DIODE(_2570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3911__A (.DIODE(_2571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3186__B (.DIODE(_2571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2982__B (.DIODE(_2571_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_A (.DIODE(_2576_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_A (.DIODE(_2576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5768__S (.DIODE(_2579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5759__S (.DIODE(_2579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3760__A (.DIODE(_2579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3759__A (.DIODE(_2579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3752__A (.DIODE(_2579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3751__A (.DIODE(_2579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2990__B (.DIODE(_2579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5783__A_N (.DIODE(_2580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5563__A (.DIODE(_2580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5015__A (.DIODE(_2580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4534__B1 (.DIODE(_2580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2991__B (.DIODE(_2580_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout49_A (.DIODE(_2581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3598__S (.DIODE(_2582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3596__S (.DIODE(_2582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3594__S (.DIODE(_2582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3592__S (.DIODE(_2582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3590__S (.DIODE(_2582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3588__S (.DIODE(_2582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3586__S (.DIODE(_2582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3584__S (.DIODE(_2582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3029__B1 (.DIODE(_2582_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_A (.DIODE(_2583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3341__B2 (.DIODE(_2583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3398__B2 (.DIODE(_2583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3455__A1 (.DIODE(_2583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5723__A (.DIODE(_2584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4244__A (.DIODE(_2584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__C (.DIODE(_2584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3771__A (.DIODE(_2584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3000__A (.DIODE(_2584_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_A (.DIODE(_2585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3563__B2 (.DIODE(_2585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4528__A2 (.DIODE(_2586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3483__A1 (.DIODE(_2586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3375__A1 (.DIODE(_2586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3177__B (.DIODE(_2586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3176__B (.DIODE(_2586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3000__B (.DIODE(_2586_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout162_A (.DIODE(_2587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5643__A1 (.DIODE(_2587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5654__A1 (.DIODE(_2587_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_A (.DIODE(_2588_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_A (.DIODE(_2588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__A (.DIODE(_2590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5118__A2 (.DIODE(_2590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__C1 (.DIODE(_2590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4529__B (.DIODE(_2590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4458__B1 (.DIODE(_2590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3012__B (.DIODE(_2590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3011__B (.DIODE(_2590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3002__B (.DIODE(_2590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3001__B (.DIODE(_2590_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(_2596_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(_2596_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_A (.DIODE(_2596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5561__A1 (.DIODE(_2596_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_A (.DIODE(_2597_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_A (.DIODE(_2597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3166__B (.DIODE(_2597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5747__A3 (.DIODE(_2599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3238__A (.DIODE(_2599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3069__B (.DIODE(_2599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3068__B (.DIODE(_2599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3067__B (.DIODE(_2599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3015__C_N (.DIODE(_2599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3917__B (.DIODE(_2600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__A (.DIODE(_2600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3238__B (.DIODE(_2600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3096__B (.DIODE(_2600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3015__A (.DIODE(_2600_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(_2601_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_A (.DIODE(_2601_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_A (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5433__C1 (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3998__A1 (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__B (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5023__B (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5745__C (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__C1 (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5388__C1 (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__C1 (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5270__C1 (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__B2 (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5007__C (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5004__B (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4933__B1 (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__C (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5122__A2 (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5116__A2 (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5090__C_N (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5021__A3 (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__B (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5019__A3 (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__B1 (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__B (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3038__B1 (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3024__B2 (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire161_A (.DIODE(_2609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__A1 (.DIODE(_2609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__A1 (.DIODE(_2609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3750__B1 (.DIODE(_2609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5755__A (.DIODE(_2610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__B1 (.DIODE(_2610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__B (.DIODE(_2610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4493__A2 (.DIODE(_2610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3928__A2 (.DIODE(_2610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__B (.DIODE(_2610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3100__B (.DIODE(_2610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3036__B (.DIODE(_2610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3021__B (.DIODE(_2610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__A (.DIODE(_2612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5347__B1 (.DIODE(_2612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__A1 (.DIODE(_2612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__B2 (.DIODE(_2612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5191__B1 (.DIODE(_2612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5174__C (.DIODE(_2612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5101__A1 (.DIODE(_2612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4501__A2 (.DIODE(_2612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__B (.DIODE(_2612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__C (.DIODE(_2612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__A2 (.DIODE(_2615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4951__A2 (.DIODE(_2615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__A2 (.DIODE(_2615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4891__A2 (.DIODE(_2615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__A2 (.DIODE(_2615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4677__A2 (.DIODE(_2615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4557__A1 (.DIODE(_2615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__A2 (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4769__A2 (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__A2 (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4688__A2 (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__B1 (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4602__A2 (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4556__A1 (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3039__A1 (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3027__A2 (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5693__A2 (.DIODE(_2618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4012__A2 (.DIODE(_2618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__A2 (.DIODE(_2618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3029__A2 (.DIODE(_2618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3060__S (.DIODE(_2619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3057__S (.DIODE(_2619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3054__S (.DIODE(_2619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3051__S (.DIODE(_2619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3048__S (.DIODE(_2619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3045__S (.DIODE(_2619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3042__S (.DIODE(_2619_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap47_A (.DIODE(_2623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4398__A (.DIODE(_2623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5694__A0 (.DIODE(_2625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4013__A1 (.DIODE(_2625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3990__A1 (.DIODE(_2625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3875__A1 (.DIODE(_2625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__A0 (.DIODE(_2625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3602__A0 (.DIODE(_2625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3575__A0 (.DIODE(_2625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3042__A1 (.DIODE(_2625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5453__A1 (.DIODE(_2627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5383__A1 (.DIODE(_2627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5348__B2 (.DIODE(_2627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5321__A (.DIODE(_2627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__A1 (.DIODE(_2627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5256__A1 (.DIODE(_2627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__A1 (.DIODE(_2627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__A1 (.DIODE(_2627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__A3 (.DIODE(_2627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3038__A2 (.DIODE(_2627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3873__C (.DIODE(_2631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3786__A1 (.DIODE(_2631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3600__A (.DIODE(_2631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3573__A (.DIODE(_2631_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_A (.DIODE(_2632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5574__A1 (.DIODE(_2632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3044__A0 (.DIODE(_2632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__A0 (.DIODE(_2633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4014__A1 (.DIODE(_2633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3991__A1 (.DIODE(_2633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3876__A1 (.DIODE(_2633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3788__A0 (.DIODE(_2633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3603__A0 (.DIODE(_2633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3576__A0 (.DIODE(_2633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3045__A1 (.DIODE(_2633_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_A (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__A1 (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3047__A0 (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_A (.DIODE(_2636_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_A (.DIODE(_2636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__A1 (.DIODE(_2636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3050__A0 (.DIODE(_2636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5697__A0 (.DIODE(_2637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4016__A1 (.DIODE(_2637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3993__A1 (.DIODE(_2637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3878__A1 (.DIODE(_2637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__A0 (.DIODE(_2637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3605__A0 (.DIODE(_2637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3578__A0 (.DIODE(_2637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3051__A1 (.DIODE(_2637_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_A (.DIODE(_2638_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_A (.DIODE(_2638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5613__A1 (.DIODE(_2638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3053__A0 (.DIODE(_2638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5698__A0 (.DIODE(_2639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__A1 (.DIODE(_2639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3994__A1 (.DIODE(_2639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3879__A1 (.DIODE(_2639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__A0 (.DIODE(_2639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3606__A0 (.DIODE(_2639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3579__A0 (.DIODE(_2639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3054__A1 (.DIODE(_2639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__A0 (.DIODE(_2641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4018__A1 (.DIODE(_2641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3995__A1 (.DIODE(_2641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__A1 (.DIODE(_2641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__A0 (.DIODE(_2641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3607__A0 (.DIODE(_2641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3580__A0 (.DIODE(_2641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3057__A1 (.DIODE(_2641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__A0 (.DIODE(_2643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4019__A1 (.DIODE(_2643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3996__A1 (.DIODE(_2643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__A1 (.DIODE(_2643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3793__A0 (.DIODE(_2643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3608__A0 (.DIODE(_2643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3581__A0 (.DIODE(_2643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3060__A1 (.DIODE(_2643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5705__A (.DIODE(_2647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3226__A (.DIODE(_2647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3065__B (.DIODE(_2647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5153__S (.DIODE(_2649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4539__A (.DIODE(_2649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3199__B (.DIODE(_2649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3108__A2 (.DIODE(_2649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3735__B (.DIODE(_2653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3449__A (.DIODE(_2653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3390__B2 (.DIODE(_2653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3288__A (.DIODE(_2653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3286__A1 (.DIODE(_2653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3239__A0 (.DIODE(_2653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3072__B (.DIODE(_2653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__B2 (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3648__A1 (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3620__A (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3619__A (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3074__B (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3073__B (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3375__B1 (.DIODE(_2660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3320__A (.DIODE(_2660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3079__C (.DIODE(_2660_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_A (.DIODE(_2661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3187__A1 (.DIODE(_2661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3929__B (.DIODE(_2661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3080__C (.DIODE(_2661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5641__A1 (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5547__C1 (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4513__A (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3948__A1 (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3736__A (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3081__B (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3916__B (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3648__A2 (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3613__A (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3612__A (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3083__B (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3082__B (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3202__A1 (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3156__A (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3154__A (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3148__A (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3147__A (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3128__A (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3117__A (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3116__A (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3095__A (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout74_A (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5608__A1 (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5607__A (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__A1 (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__A (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__A (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3633__A (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3632__A (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3618__A (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3617__A (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3156__B (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3154__B (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3095__B (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3869__S (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3866__S (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__S (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3860__S (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3857__S (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3854__S (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3851__S (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3842__S (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3094__B (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3633__B (.DIODE(_2677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3632__B (.DIODE(_2677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3618__B (.DIODE(_2677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3617__B (.DIODE(_2677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3156__C (.DIODE(_2677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3154__C (.DIODE(_2677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3095__C (.DIODE(_2677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3626__A (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3625__A (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3200__A (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3117__B (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3116__B (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3108__C1 (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__A1 (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__A2 (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__B (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3158__B (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3105__B (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4658__B (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3105__C (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3158__C (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__A2 (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4786__S (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__A2 (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__A2 (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4561__A (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3115__C (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5750__B1 (.DIODE(_2689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__B2 (.DIODE(_2689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5388__A1 (.DIODE(_2689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__A1 (.DIODE(_2689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5270__B2 (.DIODE(_2689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5134__A2 (.DIODE(_2689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__A (.DIODE(_2690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__B (.DIODE(_2690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3199__C (.DIODE(_2690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3108__A3 (.DIODE(_2690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5786__A2 (.DIODE(_2696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__B2 (.DIODE(_2696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5172__B1 (.DIODE(_2696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4531__C (.DIODE(_2696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3847__C (.DIODE(_2696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3841__A (.DIODE(_2696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3639__A (.DIODE(_2696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3621__C (.DIODE(_2696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3164__C (.DIODE(_2696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5561__A2 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__A (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__A1 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3115__D (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5825__A_N (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3757__C (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__C (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3396__A1 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3339__A1 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5189__B (.DIODE(_2703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5188__A2 (.DIODE(_2703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__B (.DIODE(_2703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3123__A2 (.DIODE(_2703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3455__B2 (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3292__B1 (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3243__B2 (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3141__B2 (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3134__B1 (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3123__B1 (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3248__A2_N (.DIODE(_2706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3171__A3 (.DIODE(_2706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3168__A3 (.DIODE(_2706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3125__B (.DIODE(_2706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3124__B (.DIODE(_2706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3255__A1 (.DIODE(_2707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3251__A1 (.DIODE(_2707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3239__S (.DIODE(_2707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3163__A (.DIODE(_2707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3153__A (.DIODE(_2707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3126__B (.DIODE(_2707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3647__A2 (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3627__A (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3128__B (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5187__B (.DIODE(_2715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5186__B (.DIODE(_2715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3133__B (.DIODE(_2715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3248__B1 (.DIODE(_2716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3135__A (.DIODE(_2716_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout112_A (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3136__A2 (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3629__A1 (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3540__B1 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3539__B1 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3183__A1 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3180__A (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3144__B1 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__B (.DIODE(_2721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__B (.DIODE(_2721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3141__A2 (.DIODE(_2721_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_A (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5650__A1 (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5540__A0 (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__B (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__A (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3636__A (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3157__B2 (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5540__A1 (.DIODE(_2746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__B (.DIODE(_2746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4561__B (.DIODE(_2746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__A1 (.DIODE(_2746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3165__A1 (.DIODE(_2746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3909__D (.DIODE(_2759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3757__D (.DIODE(_2759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3478__B (.DIODE(_2759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3191__D (.DIODE(_2759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3190__B (.DIODE(_2759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__B (.DIODE(_2764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3482__A1 (.DIODE(_2764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3265__B1 (.DIODE(_2764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3966__C (.DIODE(_2765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3564__A1 (.DIODE(_2765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3522__B1 (.DIODE(_2765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3419__A (.DIODE(_2765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3368__B (.DIODE(_2765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3319__A1 (.DIODE(_2765_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout159_A (.DIODE(_2769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3322__S (.DIODE(_2769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3484__B1 (.DIODE(_2769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5798__C1 (.DIODE(_2771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5542__A2 (.DIODE(_2771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3897__A (.DIODE(_2771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3643__A1 (.DIODE(_2771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3189__A1 (.DIODE(_2771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5725__A1 (.DIODE(_2772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5706__B2 (.DIODE(_2772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3230__A1 (.DIODE(_2772_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout67_A (.DIODE(_2778_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout66_A (.DIODE(_2778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5723__B (.DIODE(_2785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5702__B (.DIODE(_2785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3203__B (.DIODE(_2785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3570__A2 (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3533__A2 (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3488__A2 (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3434__A2 (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3381__A2 (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3325__A2 (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3277__A2 (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3231__A2 (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_A (.DIODE(_2800_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout107_A (.DIODE(_2800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__C1 (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__C1 (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__C1 (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3441__A1 (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3329__C1 (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3236__S (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__A1_N (.DIODE(_2804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3655__B1 (.DIODE(_2804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3228__C (.DIODE(_2804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4515__A (.DIODE(_2805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4514__A (.DIODE(_2805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4020__B (.DIODE(_2805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3912__A (.DIODE(_2806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3225__B (.DIODE(_2806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3224__B (.DIODE(_2806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5761__A (.DIODE(_2810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5012__B (.DIODE(_2810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__B1 (.DIODE(_2810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4511__B1 (.DIODE(_2810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3228__D_N (.DIODE(_2810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5444__A1_N (.DIODE(_2818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3658__A1 (.DIODE(_2818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3237__A2 (.DIODE(_2818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5229__B (.DIODE(_2823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5228__B (.DIODE(_2823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5227__B (.DIODE(_2823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3243__A2 (.DIODE(_2823_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout106_A (.DIODE(_2826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__C (.DIODE(_2826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3854__A0 (.DIODE(_2826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3957__B1 (.DIODE(_2826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3349__A2 (.DIODE(_2830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3348__B (.DIODE(_2830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3297__B (.DIODE(_2830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3288__C (.DIODE(_2830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3286__A2 (.DIODE(_2830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5570__A0 (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__B (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__B (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__B (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3664__A (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3254__A2 (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5570__A1 (.DIODE(_2838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4573__B (.DIODE(_2838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__B (.DIODE(_2838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3666__A1 (.DIODE(_2838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3257__A1 (.DIODE(_2838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3745__B (.DIODE(_2851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__B (.DIODE(_2851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3563__C1 (.DIODE(_2851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3321__A1 (.DIODE(_2851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3270__B1 (.DIODE(_2851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5799__A2 (.DIODE(_2856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5572__A2 (.DIODE(_2856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3897__B (.DIODE(_2856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3667__A1 (.DIODE(_2856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3275__A1 (.DIODE(_2856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5727__A1 (.DIODE(_2857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__A1 (.DIODE(_2857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3276__A2 (.DIODE(_2857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__B1 (.DIODE(_2865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3670__A (.DIODE(_2865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3285__A2 (.DIODE(_2865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__B (.DIODE(_2871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5258__B (.DIODE(_2871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__B (.DIODE(_2871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3293__A2 (.DIODE(_2871_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout103_A (.DIODE(_2874_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout102_A (.DIODE(_2874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3295__A2 (.DIODE(_2874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3374__A1 (.DIODE(_2874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5582__A0 (.DIODE(_2882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__A2 (.DIODE(_2882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4621__B (.DIODE(_2882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4620__B (.DIODE(_2882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3677__A (.DIODE(_2882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3303__A2 (.DIODE(_2882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5582__A1 (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4655__A2 (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__B (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__B (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3679__A1 (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3306__A1 (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5801__B2 (.DIODE(_2903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5800__A (.DIODE(_2903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5584__A2 (.DIODE(_2903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3897__C (.DIODE(_2903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3680__A0 (.DIODE(_2903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3323__A1 (.DIODE(_2903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5729__A1 (.DIODE(_2904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5710__A1 (.DIODE(_2904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3324__A2 (.DIODE(_2904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__A1 (.DIODE(_2910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3682__A (.DIODE(_2910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3331__B (.DIODE(_2910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__B (.DIODE(_2920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__B (.DIODE(_2920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3341__B1 (.DIODE(_2920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4661__B (.DIODE(_2932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3689__A1 (.DIODE(_2932_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout296_A (.DIODE(\as2650.addr_buff[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4907__A (.DIODE(\as2650.addr_buff[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout295_A (.DIODE(\as2650.addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5436__A1 (.DIODE(\as2650.addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5451__A1 (.DIODE(\as2650.addr_buff[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__A (.DIODE(\as2650.addr_buff[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__A1 (.DIODE(\as2650.addr_buff[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4933__A1 (.DIODE(\as2650.addr_buff[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4912__B1 (.DIODE(\as2650.addr_buff[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4907__C (.DIODE(\as2650.addr_buff[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4464__A1 (.DIODE(\as2650.addr_buff[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5490__A (.DIODE(\as2650.addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5489__A1 (.DIODE(\as2650.addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__A1 (.DIODE(\as2650.addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5464__B1 (.DIODE(\as2650.addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__A1 (.DIODE(\as2650.addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4964__A (.DIODE(\as2650.addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4951__B2 (.DIODE(\as2650.addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4941__C1 (.DIODE(\as2650.addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4939__B1 (.DIODE(\as2650.addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4465__A1 (.DIODE(\as2650.addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__A1 (.DIODE(\as2650.addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5490__B (.DIODE(\as2650.addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5489__B1 (.DIODE(\as2650.addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__A1 (.DIODE(\as2650.addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__B2 (.DIODE(\as2650.addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__A (.DIODE(\as2650.addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4968__A (.DIODE(\as2650.addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__A (.DIODE(\as2650.addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__A1 (.DIODE(\as2650.addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5515__A1 (.DIODE(\as2650.addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__A (.DIODE(\as2650.addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5032__A1 (.DIODE(\as2650.addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4467__A1 (.DIODE(\as2650.addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3151__A_N (.DIODE(\as2650.addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3150__B (.DIODE(\as2650.addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3149__B (.DIODE(\as2650.addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3092__B (.DIODE(\as2650.addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5530__A1 (.DIODE(\as2650.addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5346__A (.DIODE(\as2650.addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__A1 (.DIODE(\as2650.addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__A1 (.DIODE(\as2650.addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3151__B (.DIODE(\as2650.addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3150__A_N (.DIODE(\as2650.addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3149__A_N (.DIODE(\as2650.addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3092__A (.DIODE(\as2650.addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout291_A (.DIODE(\as2650.cycle[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__A (.DIODE(\as2650.cycle[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__A_N (.DIODE(\as2650.cycle[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5098__A1 (.DIODE(\as2650.cycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__B (.DIODE(\as2650.cycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__A (.DIODE(\as2650.cycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__B (.DIODE(\as2650.cycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3087__B (.DIODE(\as2650.cycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3018__A (.DIODE(\as2650.cycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3003__A (.DIODE(\as2650.cycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2978__A (.DIODE(\as2650.cycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2946__A (.DIODE(\as2650.cycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout293_A (.DIODE(\as2650.halted ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2944__A (.DIODE(\as2650.halted ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3774__A (.DIODE(\as2650.halted ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5051__A1 (.DIODE(\as2650.holding_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3374__A0 (.DIODE(\as2650.holding_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3372__A (.DIODE(\as2650.holding_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3361__A (.DIODE(\as2650.holding_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3360__A (.DIODE(\as2650.holding_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3359__A (.DIODE(\as2650.holding_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout308_A (.DIODE(\as2650.ins_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout307_A (.DIODE(\as2650.ins_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout301_A (.DIODE(\as2650.ins_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3183__D1 (.DIODE(\as2650.ins_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3186__A (.DIODE(\as2650.ins_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3269__A (.DIODE(\as2650.ins_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3481__A1 (.DIODE(\as2650.ins_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout299_A (.DIODE(\as2650.ins_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3114__B (.DIODE(\as2650.ins_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2995__A_N (.DIODE(\as2650.ins_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5835__B1 (.DIODE(\as2650.psl[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5573__A0 (.DIODE(\as2650.psl[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3971__A1 (.DIODE(\as2650.psl[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__A (.DIODE(\as2650.psl[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__A1 (.DIODE(\as2650.psl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5784__A1 (.DIODE(\as2650.psl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__A0 (.DIODE(\as2650.psl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3970__B2 (.DIODE(\as2650.psl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3540__A1 (.DIODE(\as2650.psl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3539__A1 (.DIODE(\as2650.psl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3144__A1 (.DIODE(\as2650.psl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3143__A (.DIODE(\as2650.psl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3137__A (.DIODE(\as2650.psl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout258_A (.DIODE(\as2650.r0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout255_A (.DIODE(\as2650.r0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout254_A (.DIODE(\as2650.r0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout253_A (.DIODE(\as2650.r0[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout251_A (.DIODE(\as2650.r0[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_A (.DIODE(\as2650.r0[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout245_A (.DIODE(\as2650.r0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout244_A (.DIODE(\as2650.r0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_A (.DIODE(\as2650.r0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4096__A1 (.DIODE(\as2650.r0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout242_A (.DIODE(\as2650.r0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout240_A (.DIODE(\as2650.r0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__A1 (.DIODE(\as2650.r0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3904__B (.DIODE(\as2650.r0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5710__B2 (.DIODE(\as2650.r123[1][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3242__A0 (.DIODE(\as2650.r123[1][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(io_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(io_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(io_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(io_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(io_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(io_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(io_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(io_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(io_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(rst));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout350_A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout349_A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__5809__A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__5777__B2 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout346_A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout340_A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout337_A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout334_A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout331_A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout330_A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__5642__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__5057__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout327_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__5143__B2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout348_A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout347_A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__2957__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_output11_A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_output14_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__4677__A1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__4649__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__4648__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__2951__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_output15_A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__4728__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__4727__B (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__4725__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__4700__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__4689__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__4688__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_output16_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__4763__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__4728__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__4727__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__2950__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_output17_A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__4799__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__4778__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__4769__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__4766__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_output18_A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__4838__B (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__4837__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__4833__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__4802__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_output19_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__4877__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__4838__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_output20_A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__4891__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__4878__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_output21_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__4937__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__4932__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__4903__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__2949__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_output22_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__4951__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__2948__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_output24_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__4988__A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__4983__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_output26_A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__5028__A0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__5019__A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_output30_A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__5636__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__3963__B2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__2933__A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__5720__B (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__5716__B (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__5712__B (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__5709__A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__5711__A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__5730__B (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__5734__B (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__5728__B (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__5732__A2_N (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__5726__B (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__4764__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__4687__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__B (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__4191__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__4114__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__4060__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__4032__A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__4042__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__4365__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__4381__B2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__4342__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__4312__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__4279__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout44_A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__5181__A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__A2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__B (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__5538__B (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__5524__A2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__5523__C1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__A2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__5463__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__5461__B1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout45_A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__5306__B1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__5183__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__5338__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__B1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__3053__S (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__3050__S (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__3047__S (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__3044__S (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__3035__S (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__4011__B (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__5693__A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__3988__B (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__3872__C (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__3785__A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__3056__S (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__3059__S (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout48_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__3599__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__5658__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__3572__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__2992__B (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__B2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__5203__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__5270__A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__4872__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__A1_N (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__5025__C_N (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__4893__A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__A2_N (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__A2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__B (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__A2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__4762__A2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__A2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__4685__A2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__4646__A2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__A2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__4610__A2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__4960__A2_N (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__3841__B (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__4987__A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout51_A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__4936__A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__B1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__5584__B1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__5572__B1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__5542__B1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__4986__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__4924__B1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__C1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__4751__B1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__B1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__4451__A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__4461__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__5648__B1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__5635__B1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__5622__B1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__C1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__5574__B1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__5812__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__3980__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__3912__B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__5817__A2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__5784__A3 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__3739__B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__3948__B2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__5650__C1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout55_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__5101__A2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__5395__A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__5522__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__5445__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__5482__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__5422__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__5336__A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__5305__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__5247__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__5182__A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__5461__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__5213__A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__5462__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__5483__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__5523__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__5537__S (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__S (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__5423__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__B1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5446__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout58_A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__C1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__4935__C1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5506__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__5306__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__5444__B1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__4487__A3 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout60_A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__B1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__5579__B1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__5567__A2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__A1_N (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__B2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__5655__A2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__A2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__B1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__3836__B (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__5644__A2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5504__A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5304__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__3755__B (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout64_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__A2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__5743__A2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__3237__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__3224__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__5651__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__5599__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__5575__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__5546__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__3227__B (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__3225__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__3197__B (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout68_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout69_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__5624__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__5610__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__5611__A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__5594__A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5582__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5540__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5633__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5570__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3090__B (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__B2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__4744__B2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5646__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5620__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5595__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout72_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5136__A2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__4911__B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__4906__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__4451__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__B2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__B2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4941__B2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4850__B2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3798__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__5517__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__5477__C1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__5237__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__B2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__B2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__4893__B2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__B2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__5501__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__5297__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__5154__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__4760__B2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__B2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__4553__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__4549__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__B1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5065__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5441__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5743__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5418__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5496__B1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout76_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__B1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__5481__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__5533__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__5521__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__2990__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__5840__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__5776__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout77_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__B2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__C1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5742__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3764__A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__4495__A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__4992__B (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5090__A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__A2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__C1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3916__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__B (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__5036__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3983__C1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4507__A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3756__A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3933__A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__5827__A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4021__A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__5843__A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__5847__A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3947__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3895__A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout81_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout79_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout80_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__B (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__B2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5437__A1_N (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5512__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5382__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5348__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__B2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5256__B2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5194__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5453__B2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout83_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4554__B (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4979__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4952__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4892__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__A3 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__C (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__5088__B1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__C1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4923__B1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4888__B1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4795__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4750__B1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4567__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4885__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__B1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4925__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4862__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4824__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4823__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4721__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4674__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4949__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__5077__B1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__4457__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__B (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__5032__A2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3938__D (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3847__B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__4960__B2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__4924__C1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__B2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__4834__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__4526__B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3836__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4525__B (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__B2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__B2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4762__B2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__B2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4685__B2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4646__B2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4610__B2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__B2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4987__B2 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__4457__C1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3812__B (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__4945__B2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__4884__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__4651__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__B2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__4568__A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__4851__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__5742__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__B (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3938__B (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3746__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4489__B (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4495__B (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__D (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3839__B (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__C (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3511__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3508__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3505__B (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3504__B (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3503__B (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3506__B (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5644__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3535__S (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3498__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3727__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3707__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3542__A2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3459__A2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__A0 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3981__A1_N (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__5793__A0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3524__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3514__B (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3513__B (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3866__A0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout94_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout93_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3697__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3718__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3501__A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__A0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3467__A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3465__A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3450__B1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3448__C (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3444__B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3400__A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3399__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__A0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3959__B1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3480__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3471__B (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__B (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3450__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3448__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3444__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3409__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3407__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3405__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3404__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3391__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3403__A_N (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__B2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3708__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3686__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3342__A2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3460__A2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__5600__A0 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout98_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout99_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3860__A0 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__A2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5792__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3425__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3424__A2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3414__B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3413__B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout100_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3401__A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3356__B (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3351__B (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3349__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3348__C (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3346__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3345__D (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3334__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5603__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3857__A0 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3373__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3361__B (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3698__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3360__B (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__A0 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3359__B (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3959__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__D (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3289__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout104_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3246__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3343__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__B2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5600__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__A0 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3687__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3661__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3364__B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3318__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3308__B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3307__B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout105_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3221__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__5762__B2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__5303__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__5334__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__5166__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3387__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3438__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3494__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3284__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3330__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3883__A2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3561__A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3553__B (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3552__B (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3717__A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__B (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3144__A2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__A2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3903__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__5641__A2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3960__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout109_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5810__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5655__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3869__A0 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3550__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3547__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3546__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3536__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3544__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3296__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3272__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3266__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3675__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3258__B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3259__B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3957__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout111_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3851__A0 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5579__B2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3346__A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3345__B (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3299__A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3287__B (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3250__B (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3249__B (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3240__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3173__B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5567__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3842__A0 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3250__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3346__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3345__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3299__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3287__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3249__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3247__A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3540__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3960__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__5810__A0 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3539__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3662__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__C1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5577__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5549__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3982__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__4502__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__B (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3099__B (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5106__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5004__C (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5467__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5529__C (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5514__A3 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5495__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__B2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5148__B2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3127__B (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__C (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__B2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__A1_N (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__5452__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__5437__B2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__A1_N (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__5019__A4 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__5036__B2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3935__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3927__B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__5108__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5481__C1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5501__C1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5521__C1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5533__C1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5419__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__B2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5297__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__C1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__4550__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3013__B (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5456__B1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__C1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__C1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5327__C1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5271__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__B (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3014__B (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5192__S (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__B2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__A1_N (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3025__B (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__5019__A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__A1_N (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3031__A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__4455__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5116__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5021__A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5235__A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5346__B (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__B (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5291__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__3641__B (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__5635__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__5648__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__5622__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__5584__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__5572__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__4500__A2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__5542__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__5451__S (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__4754__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__4602__B2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__4556__A0 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__4675__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__A2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__4676__A3 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__B (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__B (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5067__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__B (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__4890__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__4950__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__S (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__B (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5402__B (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__S (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5515__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5347__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5530__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__4753__B (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5385__S (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5319__S (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5232__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5190__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5436__S (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__A2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3008__C (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__C (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__5606__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__5595__C1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__5541__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__5571__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__5634__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__B (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__4487__A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3113__B (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__5647__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__5608__C1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__5583__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__5476__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__5454__B2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__5296__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__C1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__C1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__5269__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__B (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__5499__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__5067__C1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5021__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__B1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5456__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__B1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__4452__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5514__B1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__B (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__C1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5417__B1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5386__A1_N (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5326__A1_N (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5013__B (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5224__B1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__4454__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__B (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__5106__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__C (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__5010__A3 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__3008__B (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__3039__B2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__5517__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__5174__B (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__5116__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__5087__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__5530__D1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__5443__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__5349__C1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__4547__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__5149__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__3806__B (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__5159__A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4547__C1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__B2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__B2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4643__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4554__A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4607__A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__B (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5169__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__4530__A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__4487__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__4458__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5136__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__3834__B (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5760__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__3920__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__5532__C (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__3227__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__3107__B (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__5349__B2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__5358__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__5057__S (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__5059__S (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__5053__A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__5047__A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__5828__A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__3063__B (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__3644__A3 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__3780__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__5832__A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__3922__B (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__3907__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__3979__S (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__3946__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__5826__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__5838__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5769__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__B (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5841__A2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5770__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__4502__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__3774__B (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__3908__A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2979__B (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__5430__A1_N (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__5426__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__4933__C1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__C1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__4951__C1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__4891__C1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__C1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5417__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5517__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__A2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5013__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5066__B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__4487__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3935__B2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__C (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5093__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__4502__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__4644__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__4609__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5615__B1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3966__D (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3936__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3911__B (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3745__C (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5169__A3 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4513__B (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__C (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__3839__C (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__B1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__B1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5567__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5654__B1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5642__B1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5602__B1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__3280__B1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__A3 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5163__B1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3491__B1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5273__B1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3384__B1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3439__B1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3437__B1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__B1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__B1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout155_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout156_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__B1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__4432__C (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__B1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__B1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__B1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5242__B1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3571__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3385__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3281__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3219__A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5332__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5274__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5164__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3218__A_N (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3217__A_N (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3485__A1_N (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__3530__S (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__3429__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__3378__S (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__3430__A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__3566__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__3273__A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__3188__A2_N (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__3187__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__3567__A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5604__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5579__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5568__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4488__B (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4958__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__2999__C (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__C (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5039__C (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3777__C (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3772__B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__2980__B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5106__A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4521__A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4500__A1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3998__D1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5007__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3811__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3810__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3023__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3022__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__2977__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__B (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3777__B (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5039__B (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3772__A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3809__B (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__2980__A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__2978__B (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3234__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__3872__B (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5163__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__3491__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5273__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__3384__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__3439__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__3437__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__2969__B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__4415__B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__3492__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3440__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3385__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3436__B1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5164__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3281__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3328__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__3282__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5274__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5657__B (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5363__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5301__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5332__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__3440__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__3328__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__3283__B1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__3235__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__4011__C (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__4012__A3 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5363__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5301__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5242__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__3490__C (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__3383__C (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__3209__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5272__C (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__C (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__C (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__C (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__C (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__4470__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__3210__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__3215__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__3279__C (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__3211__C (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4211__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4177__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4176__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4353__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4354__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__3244__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__3142__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__A3 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5553__A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__3193__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__3115__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__3647__B1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__3065__A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__3648__C1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__3611__A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__3134__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__3118__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__3398__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__3456__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__3341__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__3292__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4255__D (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__D (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4161__B1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4221__D (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4222__B1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4284__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4285__D (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4367__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4286__B1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4344__B1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4256__B1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4122__D (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__B1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__A1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__3059__A0 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4345__D (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4087__B1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4314__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4286__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4256__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4255__C (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4222__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4221__C (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__C (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4161__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4285__C (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4122__C (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4088__D (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3396__B1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4344__A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4345__C (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__5625__A1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3056__A0 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4261__A2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__A2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4164__B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4220__B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4348__A2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4318__B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4289__B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4288__B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4088__C (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__3339__B1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4087__A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4062__B (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4124__B (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4123__A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4064__D (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__B1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__B1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__D (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__4253__D (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__4252__B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__4215__B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__4214__B1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__4129__B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__4128__B1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__4092__C (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__4064__C (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__D (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__4046__C (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__4065__C (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__4063__A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__4035__B1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__C (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4128__A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4090__B (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4253__C (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4251__B (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4214__A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4153__B (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__B (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4095__B (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4096__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4157__A2_N (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4156__D (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__B (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4247__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4218__B (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4117__C1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4119__A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4103__A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4102__C1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4072__B (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4106__A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4044__B (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4036__B (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4173__B (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4174__B (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4028__A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__4029__C (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__4027__A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__5545__A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3035__A0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__5706__A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__A1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__4984__C1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__C1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__4833__B1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__C1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__B2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__C1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__B2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__4639__B1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__4606__C1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__4000__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__3938__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__3000__C (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__3527__B2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__3427__B2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__3319__B2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__3267__B2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__3184__B2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__3183__C1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__3182__B (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__3181__B (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__5786__A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__2999__B (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__3293__A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__3243__A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__3123__A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__3133__A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__3141__A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__3967__A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__3909__C (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__3753__C (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__3746__A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__2999__A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__3364__A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__3271__B (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__3168__A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__3167__B (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__3924__A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__3917__A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__3110__A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__3223__B (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__3192__A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__3882__B (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__3523__B (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__3479__S (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__3423__B (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__3372__B (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__3425__S (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__3424__A1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__3373__A1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__3318__S (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__3374__S (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__3363__B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__3266__S (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__3272__A1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__3170__B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__3171__A1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__3480__S (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__3524__A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__S (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__3561__S (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__3883__A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__3191__B (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__3115__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__3072__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5036__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__3909__B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__3757__B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__3753__B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__3193__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__2989__B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5551__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__3109__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__2997__B (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__4985__A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__4954__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__4898__A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__4829__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__4525__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__3806__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__5026__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__B1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__3907__C1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__3091__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__3080__B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5785__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__3067__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__3070__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4992__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4533__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4528__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__B2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__3099__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4549__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__3106__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__3014__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__3013__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5161__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4555__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__2997__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5747__C1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__3830__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__3081__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__5762__C1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__5174__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__5753__A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__5079__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__4490__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__3740__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__4547__B1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__3037__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__3024__A1_N (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__3002__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__3001__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__3741__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__3966__B (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__3944__B (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__3745__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__3735__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__3079__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__3242__S1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__3052__S (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__3228__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__3063__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__4021__A1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__3046__S (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5829__A1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__3972__B2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__3616__A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__3609__A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__3166__A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__3164__A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__2934__A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__5609__A0 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__3034__S (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__3122__S1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__3207__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__2936__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__3214__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__3208__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__3212__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__3233__S0 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__3327__S0 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__3386__S0 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__3493__S0 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__3220__S0 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__A1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__5778__C1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__S0 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__S0 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__S0 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__S0 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__S0 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__S0 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__S0 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__5767__A1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__3208__B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__3214__B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__2937__A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__2968__B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__3493__S1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__3386__S1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__3327__S1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__3233__S1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__3220__S1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__5573__A1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__3207__B (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__S1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__S1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__S1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__S1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__S1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__S1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__S1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout219_A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__3210__A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__2938__A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__4432__A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5272__A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__4415__A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__3965__B2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5585__A1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5765__A1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__3279__A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout220_A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__3066__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__3010__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__3071__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__5562__A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout222_A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout223_A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout224_A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__4534__A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__5747__A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__4526__A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__2998__B (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__5007__A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__4874__A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__4569__A1_N (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__5794__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__3901__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__2982__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__3929__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__3757__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__3909__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__3190__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__3922__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__3914__A1_N (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__A1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5808__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5821__A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5819__C1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__3191__A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5813__A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__3079__B (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5741__A0 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__B (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout227_A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout226_A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__A1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__A1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout225_A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5534__C1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5740__A0 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__2955__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__C1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__2998__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__4932__D1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5419__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__3932__A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__3918__A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__4518__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__4490__B (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__B2 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5118__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__4529__A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__2985__B (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5817__A1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5784__A2 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__3944__C (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__A (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__A (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__2986__B (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__5105__A (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout230_A (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__3983__A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__3869__A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5692__A0 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5675__A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__A0 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__4448__A0 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__4431__A0 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__4414__A0 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__3598__A0 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__4209__A0 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__4345__A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__4384__A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__4251__A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__4252__A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__4247__A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__4218__A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__4253__A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__4367__A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__4348__A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__4318__A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__3979__A0 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__4173__A (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5059__A0 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__3732__A1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__3534__A1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__3142__A1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__4174__A (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__3728__A1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout233_A (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__4344__A1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout234_A (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__3543__A0 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__2939__A (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5143__A1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5656__A1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout232_A (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__4157__A1_N (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__4345__B (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__4344__B2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__4369__A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__4370__A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__4288__A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__4289__A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__4253__B (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__4215__A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__4314__A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout236_A (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__3489__A (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5690__A0 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5673__A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__4484__A0 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__4446__A0 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__4412__A0 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__3596__A0 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__4429__A0 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__4207__A0 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5057__A0 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__4119__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__5841__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__4117__B1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3904__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3502__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3719__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3945__A0 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__5645__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3866__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3456__A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout238_A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__4214__A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__4156__C (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__3461__A1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__5632__A1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__A0 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__5671__A1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__4427__A0 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__4410__A0 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__3594__A0 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__4205__A0 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__4482__A0 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__4444__A0 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__4153__A (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__A (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__4285__A (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__4286__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__A (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__4353__A (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__4354__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__4284__A (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__3709__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__3777__A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__3398__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__4102__B1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__4103__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__3435__A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout241_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__4214__B2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__3382__A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3860__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__A0 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__5669__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__4480__A0 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__4442__A0 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__4408__A0 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3592__A0 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__4425__A0 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__4203__A0 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__4256__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__4255__A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__4261__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__4220__A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__4286__B2 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__4285__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__4128__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__4129__A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__4326__A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__4095__A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__3341__A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__4106__A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__4072__A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__3904__C (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__3402__A0 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__3699__A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__5619__A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__3688__A1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__5605__A1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__3344__A1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__3857__A1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__5684__A0 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__5667__A1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__A0 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__3590__A0 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__4423__A0 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__4201__A0 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__4128__B2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__4282__A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__4090__A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__4164__A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__4281__A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__3292__A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__3326__A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__4478__A0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__A0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__4068__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__4067__A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__4044__A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__4066__A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__4222__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__4221__A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__4255__B (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__4256__B2 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__4092__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout248_A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__3904__D (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout246_A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__5759__A0 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__A0 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__5665__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__4404__A0 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__3588__A0 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__4421__A0 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__4199__A0 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__4476__A0 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__4438__A0 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__3854__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__3278__A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__3244__A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__4222__B2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__4221__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__4249__A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__4248__A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__4161__A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__A1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4064__A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4050__A1_N (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4036__A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4049__C (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__B2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4092__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4124__A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4123__A1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4063__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__4065__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout252_A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__3302__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__A0 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__3232__A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__4474__A0 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__A0 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5680__A0 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5663__A1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__4419__A0 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__4402__A0 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__4197__A0 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__3586__A0 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5768__A0 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__4065__B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__4046__A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__4063__B2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__4035__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__4029__A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__4028__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__4088__A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__4064__B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__4087__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__3134__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout257_A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__3253__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__3663__A0 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__5581__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__3851__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__4176__A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__4177__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5678__A0 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5661__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__4400__A0 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__3584__A0 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__4195__A0 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__4417__A0 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__4472__A0 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__A0 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__4062__A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__4029__B (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__4046__B (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__4028__B2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__B2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__B2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__3229__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5039__A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__4027__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5706__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__3118__A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__4035__B2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__4087__B2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__4088__B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout260_A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout261_A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__3842__A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5569__A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__3631__A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__A3 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__3155__A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout262_A (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__3655__A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__B2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__4122__B (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout259_A (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5486__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5485__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__3053__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__A0 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__4987__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__4979__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__4972__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__A (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__3050__A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5475__B1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5484__A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5466__A0 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__4960__A1_N (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__4952__A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__4946__A (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5463__A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__3047__A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5455__A (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5450__A (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__4936__A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__2940__A (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__4915__A (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__4916__A (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5434__A (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__A (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5427__A (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__A0 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__A3 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__4919__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__4893__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__A (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__4892__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__B1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5400__A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5399__A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__A4 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__4919__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__A1_N (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__2941__A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__4852__A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__A0 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__A1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__A1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__4856__A1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__4820__A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5691__A1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5674__A1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__4413__A1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__3597__A1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__A1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__B (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5370__A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5371__B1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__4485__A1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__A1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__A1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__4208__A1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5372__A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__4856__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__A1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__A1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__A1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__4770__A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__5689__A1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__5672__A1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__A1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__3595__A1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__5341__A (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5340__A (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5370__B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5371__A1 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__4483__A1 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__A1 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__4206__A1 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__4428__A1 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__A (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout271_A (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5320__A0 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__4760__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__4762__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5670__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5687__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__A1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__B (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__5313__A1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__B (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__4479__A1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__4441__A1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__4424__A1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__4202__A1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__A1 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__4693__A (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__5668__A1 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__5685__A1 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__4407__A1 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__3591__A1 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__A1 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__A1 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__A (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__2942__A (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__A1 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__3589__A1 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__5683__A1 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__4405__A1 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__A1 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__A1 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__4685__A1 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__4670__A (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__4669__A (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__4695__A1 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__4477__A1 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__4439__A1 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__4422__A1 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__4200__A1 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__5252__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__5265__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__5266__B1 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__5249__A0 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout277_A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__5266__A1 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__A1 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5219__A0 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__4672__A1 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__4646__A1 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__4644__A1 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__4639__A1 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__B1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__4475__A1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__A1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__4420__A1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__4198__A1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout280_A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__B1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__4591__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__4589__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__A1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__5662__A1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__3585__A1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__5679__A1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__4401__A1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__4473__A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__4435__A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__4418__A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__4196__A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout282_A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout283_A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout285_A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5660__A1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__4544__A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5677__A1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__3583__A0 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__4399__A0 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__A2 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__C (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5183__A1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__4194__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__4416__A0 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__4471__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__B (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout286_A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__A1 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__C (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__C (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__3087__C_N (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__3003__B (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__5098__A2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__3018__B (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__2976__B (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__3085__B (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__3763__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__3997__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__A1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2979__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5010__A2 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5077__A1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__3017__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5066__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__5082__A2_N (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout290_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__3833__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__C1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__C1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__5082__A1_N (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__5122__B1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__C1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__5031__C1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__C1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__5134__C1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__B1 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__3644__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__3198__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__2970__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__4020__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__C1 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__4488__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__2971__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5012__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout292_A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__3090__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__3031__A1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__A0 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__4676__A1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__3026__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__3025__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5426__A1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5425__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5192__A1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__4907__B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__4891__B2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__4463__A1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__4911__A2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__A2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__5416__A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5415__A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5402__A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__A1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__4911__A1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__A1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__4847__A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__2967__A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__B2 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__3097__A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__3009__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__3098__A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__3114__C (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__2995__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5600__S (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__S (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__S (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__4010__A1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__4501__A1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__3076__A_N (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__3075__A_N (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__2996__B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__2981__B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__5810__S (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__S (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__C_N (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__3901__D (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout297_A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__3901__C (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__4009__A1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__3076__B (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__3075__B (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__2981__A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__A1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__2996__A_N (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__3009__A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__4497__A1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__3066__B (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__3935__A1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__3069__A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__3068__A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__3030__A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__3008__A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__5747__A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__4008__A1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__3773__A1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__2984__A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__2983__A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__3182__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3181__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3177__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3176__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3078__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3077__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3901__B (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3114__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3010__B (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout300_A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3080__A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__4006__A1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__5150__B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3036__A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3011__A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__C (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3012__A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__2954__A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__2986__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3734__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__B (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3096__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__5134__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__4458__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__2985__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__2993__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__2987__A_N (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__4004__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3944__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__B (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3768__B (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3223__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__2953__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3649__B1 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3062__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__5702__A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__4022__A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout306_A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3140__S0 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3242__S0 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3291__S0 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3454__S0 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3767__B (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__3766__B (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__3999__A (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__3927__A (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__2988__B (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__3946__D1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__3062__B (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__5839__A_N (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__5750__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__3928__A1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__S (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__5193__S (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__5249__S (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__S (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__5320__S (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__S (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__5146__S (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__5219__S (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__4833__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__5401__S (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__A (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__3964__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout309_A (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout310_A (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__A1_N (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__A (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__3978__A2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__3970__A2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__3960__B2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__3537__A (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout311_A (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__C1 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__5183__C1 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__3865__A (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__A (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__3868__A (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__A (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__3859__A (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__3856__A (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__3853__A (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__3850__A (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__C1 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__C1 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__4877__C1 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__4837__C1 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__C1 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__4687__C1 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__C1 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__4764__C1 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__C1 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout313_A (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__5338__C1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__C1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__C1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__C1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5539__C1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5524__C1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__C1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5424__C1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__C1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout314_A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5581__C1 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__5035__C1 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__5033__C1 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__B1 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__5139__B1 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__C1 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__A (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__4498__A (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__C1 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__A (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout316_A (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout317_A (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__C1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__A (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__4938__C1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__C1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__5484__C1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5463__C1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5447__C1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__3782__B1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5846__A (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__B1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__C1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5767__B1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__3644__B1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5850__A (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__C1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5830__A (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5834__A (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5796__C1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__3987__C1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__3955__C1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout318_A (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout320_A (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout319_A (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__B1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout315_A (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__4932__A2 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__B2 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__3038__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__3021__A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout323_A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__B (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5345__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5385__A0 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__A (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__A (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__4010__B2 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__2958__A (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__4957__A (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__4958__A2 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__4984__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5004__A (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout324_A (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5653__A0 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__A (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__A (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4810__A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__A (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4805__A (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4804__A (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4469__A0 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__A (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__3724__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5059__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout326_A (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5514__A2 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__A2 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5529__B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5532__B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout325_A (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__4916__B (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4915__B (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__B (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__B (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4852__B (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4856__B1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4820__B (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__B (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4770__B (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4769__B2 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__5840__A1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__A (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__5352__A (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__A (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__5347__A1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__4009__B2 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout328_A (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout329_A (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__C (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__3946__A2 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__3716__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__3499__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__4811__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__A1_N (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__A (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__A (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__A0 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__2966__A (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__3779__A (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__3706__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__3458__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__A0 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__4739__A (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__A (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__4732__A (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__4731__A (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__4467__A0 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__5628__A (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__B (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__3780__A2 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout332_A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout333_A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5319__A0 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__4753__A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__B (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__B (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__4007__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__2964__A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__3696__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__3393__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__4710__A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__A0 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__2963__A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout335_A (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout336_A (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__5741__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__A (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__A (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__A (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__A0 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__4693__B (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__B (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__4688__B2 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__A (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__5258__A (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__A (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__A0 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__4695__A2 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__4676__A2 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__4670__B (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__4669__B (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__4465__A0 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__5602__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__D (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__3685__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__4661__A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__4658__A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__4653__A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__4652__A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__3336__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__2962__A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5832__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5847__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5848__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout339_A (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__A0 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5740__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout338_A (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5227__A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__4006__B2 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__2961__A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5451__A0 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__A0 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__4672__A2 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__B (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__B (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__4464__A0 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__3673__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__3294__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__4655__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__4624__A0 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__4621__A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__4620__A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__C (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__5047__A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__5817__B2 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout342_A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__5228__A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__5229__A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__5235__A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout341_A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__5191__A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__5187__A (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__5186__A (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__4005__A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__5192__A0 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__4603__A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__4591__B (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__B (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__4589__B (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__4463__A0 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__B (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__3660__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__3245__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__4588__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__A (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__A (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__A (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__4573__A (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__A (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__2960__A (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__5836__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout345_A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__5436__A0 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout344_A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__3205__C1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__2970__B (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__5128__B1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__5127__A (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__A (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__A (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__5061__A (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__A (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__4505__C1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__2971__B (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__5842__C1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__5837__C1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__5822__A (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__5814__B1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__B1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__5701__B1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__4021__B1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__3206__C1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__5775__A1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__5189__A (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__5188__A1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__A (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__4003__A1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__5155__A (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__A (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__4544__B (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__B (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__A0 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__5549__A1 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__A1 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__A (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__3628__A1 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__3129__A0 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__2959__A (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__A (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__A (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__A (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__4562__A (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6067__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6132__CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_729 ();
endmodule

