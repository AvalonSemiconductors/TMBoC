// This is the unpowered netlist.
module tt2_tholin_namebadge (clk,
    rst,
    io_in,
    io_oeb,
    io_out);
 input clk;
 input rst;
 input [2:0] io_in;
 output [26:0] io_oeb;
 output [7:0] io_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire net14;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net15;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire clknet_0_clk;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire \lcd.num_state[0] ;
 wire \lcd.num_state[1] ;
 wire \lcd.rom_addr[0] ;
 wire \lcd.rom_addr[1] ;
 wire \lcd.rom_addr[3] ;
 wire \lcd.rom_addr[4] ;
 wire \lcd.rom_addr[5] ;
 wire \lcd.rom_addr[6] ;
 wire \lcd.round[0] ;
 wire \lcd.round[1] ;
 wire \lcd.s_ROM[0] ;
 wire \lcd.s_ROM[1] ;
 wire \lcd.s_ROM[2] ;
 wire \lcd.s_ROM[3] ;
 wire \lcd.s_ROM[4] ;
 wire \lcd.s_ROM[5] ;
 wire \lcd.s_ROM[6] ;
 wire \lcd.seq[0] ;
 wire \lcd.seq[1] ;
 wire \lcd.seq[2] ;
 wire \lcd.seq[3] ;
 wire \lcd.seq[4] ;
 wire \lcd.seq[5] ;
 wire \lcd.seq[6] ;
 wire \lcd.seq[7] ;
 wire \lcd.toggle ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 sky130_fd_sc_hd__nor2_4 _404_ (.A(\lcd.toggle ),
    .B(net4),
    .Y(_007_));
 sky130_fd_sc_hd__inv_2 _405_ (.A(\lcd.toggle ),
    .Y(_375_));
 sky130_fd_sc_hd__buf_2 _406_ (.A(\lcd.seq[3] ),
    .X(_376_));
 sky130_fd_sc_hd__a211o_1 _407_ (.A1(\lcd.seq[2] ),
    .A2(\lcd.seq[1] ),
    .B1(\lcd.seq[4] ),
    .C1(_376_),
    .X(_377_));
 sky130_fd_sc_hd__buf_2 _408_ (.A(\lcd.seq[5] ),
    .X(_378_));
 sky130_fd_sc_hd__inv_2 _409_ (.A(_378_),
    .Y(_379_));
 sky130_fd_sc_hd__clkbuf_2 _410_ (.A(\lcd.seq[7] ),
    .X(_380_));
 sky130_fd_sc_hd__clkbuf_4 _411_ (.A(\lcd.seq[6] ),
    .X(_381_));
 sky130_fd_sc_hd__nor2_1 _412_ (.A(_380_),
    .B(_381_),
    .Y(_382_));
 sky130_fd_sc_hd__and3b_1 _413_ (.A_N(_377_),
    .B(_379_),
    .C(_382_),
    .X(_383_));
 sky130_fd_sc_hd__or4_1 _414_ (.A(\lcd.seq[5] ),
    .B(\lcd.seq[4] ),
    .C(\lcd.seq[3] ),
    .D(\lcd.seq[2] ),
    .X(_384_));
 sky130_fd_sc_hd__and2_1 _415_ (.A(_380_),
    .B(\lcd.seq[6] ),
    .X(_385_));
 sky130_fd_sc_hd__nor2b_4 _416_ (.A(\lcd.round[0] ),
    .B_N(\lcd.round[1] ),
    .Y(_386_));
 sky130_fd_sc_hd__nor2_1 _417_ (.A(\lcd.seq[1] ),
    .B(\lcd.seq[0] ),
    .Y(_387_));
 sky130_fd_sc_hd__nand4b_4 _418_ (.A_N(_384_),
    .B(_385_),
    .C(_386_),
    .D(_387_),
    .Y(_388_));
 sky130_fd_sc_hd__nor3_1 _419_ (.A(_375_),
    .B(_383_),
    .C(_388_),
    .Y(_389_));
 sky130_fd_sc_hd__nor2_2 _420_ (.A(_007_),
    .B(_389_),
    .Y(_390_));
 sky130_fd_sc_hd__or2b_1 _421_ (.A(\lcd.seq[1] ),
    .B_N(\lcd.seq[4] ),
    .X(_391_));
 sky130_fd_sc_hd__nand2_1 _422_ (.A(_376_),
    .B(\lcd.seq[2] ),
    .Y(_392_));
 sky130_fd_sc_hd__or2b_1 _423_ (.A(\lcd.seq[4] ),
    .B_N(\lcd.seq[1] ),
    .X(_393_));
 sky130_fd_sc_hd__or2_1 _424_ (.A(\lcd.seq[3] ),
    .B(\lcd.seq[2] ),
    .X(_394_));
 sky130_fd_sc_hd__or3b_1 _425_ (.A(_380_),
    .B(\lcd.seq[6] ),
    .C_N(\lcd.seq[5] ),
    .X(_395_));
 sky130_fd_sc_hd__a221o_1 _426_ (.A1(_391_),
    .A2(_392_),
    .B1(_393_),
    .B2(_394_),
    .C1(_395_),
    .X(_396_));
 sky130_fd_sc_hd__buf_2 _427_ (.A(\lcd.seq[4] ),
    .X(_397_));
 sky130_fd_sc_hd__and3_2 _428_ (.A(_397_),
    .B(_376_),
    .C(\lcd.seq[2] ),
    .X(_398_));
 sky130_fd_sc_hd__or3b_2 _429_ (.A(\lcd.seq[5] ),
    .B(\lcd.seq[6] ),
    .C_N(_380_),
    .X(_399_));
 sky130_fd_sc_hd__or2_1 _430_ (.A(_398_),
    .B(_399_),
    .X(_400_));
 sky130_fd_sc_hd__or2b_2 _431_ (.A(\lcd.round[0] ),
    .B_N(\lcd.round[1] ),
    .X(_401_));
 sky130_fd_sc_hd__mux2_1 _432_ (.A0(_396_),
    .A1(_400_),
    .S(_401_),
    .X(_402_));
 sky130_fd_sc_hd__and2_2 _433_ (.A(_378_),
    .B(\lcd.seq[6] ),
    .X(_403_));
 sky130_fd_sc_hd__clkbuf_4 _434_ (.A(_380_),
    .X(_033_));
 sky130_fd_sc_hd__a211oi_4 _435_ (.A1(_381_),
    .A2(_398_),
    .B1(_403_),
    .C1(_033_),
    .Y(_034_));
 sky130_fd_sc_hd__xor2_1 _436_ (.A(\lcd.round[0] ),
    .B(\lcd.round[1] ),
    .X(_035_));
 sky130_fd_sc_hd__or2_1 _437_ (.A(\lcd.seq[7] ),
    .B(\lcd.seq[6] ),
    .X(_036_));
 sky130_fd_sc_hd__clkbuf_2 _438_ (.A(_036_),
    .X(_037_));
 sky130_fd_sc_hd__o21ai_1 _439_ (.A1(_397_),
    .A2(_376_),
    .B1(_378_),
    .Y(_038_));
 sky130_fd_sc_hd__or3_1 _440_ (.A(\lcd.seq[4] ),
    .B(\lcd.seq[2] ),
    .C(\lcd.seq[1] ),
    .X(_039_));
 sky130_fd_sc_hd__or4b_1 _441_ (.A(_037_),
    .B(_035_),
    .C(_038_),
    .D_N(_039_),
    .X(_040_));
 sky130_fd_sc_hd__buf_2 _442_ (.A(_378_),
    .X(_041_));
 sky130_fd_sc_hd__or3_2 _443_ (.A(_041_),
    .B(_037_),
    .C(_377_),
    .X(_042_));
 sky130_fd_sc_hd__o211a_1 _444_ (.A1(_034_),
    .A2(_035_),
    .B1(_040_),
    .C1(_042_),
    .X(_043_));
 sky130_fd_sc_hd__inv_2 _445_ (.A(\lcd.seq[6] ),
    .Y(_044_));
 sky130_fd_sc_hd__and4_2 _446_ (.A(_033_),
    .B(_379_),
    .C(_044_),
    .D(_398_),
    .X(_045_));
 sky130_fd_sc_hd__nand3b_1 _447_ (.A_N(\lcd.seq[6] ),
    .B(_378_),
    .C(_380_),
    .Y(_046_));
 sky130_fd_sc_hd__o21a_1 _448_ (.A1(_378_),
    .A2(_381_),
    .B1(_380_),
    .X(_047_));
 sky130_fd_sc_hd__o221a_1 _449_ (.A1(_385_),
    .A2(_398_),
    .B1(_046_),
    .B2(_391_),
    .C1(_047_),
    .X(_048_));
 sky130_fd_sc_hd__or2_2 _450_ (.A(_397_),
    .B(_376_),
    .X(_049_));
 sky130_fd_sc_hd__and4bb_1 _451_ (.A_N(_049_),
    .B_N(_033_),
    .C(\lcd.seq[2] ),
    .D(_403_),
    .X(_050_));
 sky130_fd_sc_hd__nor2b_4 _452_ (.A(\lcd.round[1] ),
    .B_N(\lcd.round[0] ),
    .Y(_051_));
 sky130_fd_sc_hd__buf_2 _453_ (.A(\lcd.seq[2] ),
    .X(_052_));
 sky130_fd_sc_hd__a211o_2 _454_ (.A1(_378_),
    .A2(_397_),
    .B1(\lcd.seq[6] ),
    .C1(_380_),
    .X(_053_));
 sky130_fd_sc_hd__a31o_1 _455_ (.A1(_041_),
    .A2(_376_),
    .A3(_052_),
    .B1(_053_),
    .X(_054_));
 sky130_fd_sc_hd__o311ai_4 _456_ (.A1(_045_),
    .A2(_048_),
    .A3(_050_),
    .B1(_051_),
    .C1(_054_),
    .Y(_055_));
 sky130_fd_sc_hd__o311a_1 _457_ (.A1(\lcd.seq[4] ),
    .A2(\lcd.seq[3] ),
    .A3(\lcd.seq[2] ),
    .B1(\lcd.seq[6] ),
    .C1(_378_),
    .X(_056_));
 sky130_fd_sc_hd__o31a_1 _458_ (.A1(_378_),
    .A2(\lcd.seq[4] ),
    .A3(_376_),
    .B1(_381_),
    .X(_057_));
 sky130_fd_sc_hd__or3b_1 _459_ (.A(_380_),
    .B(_056_),
    .C_N(_057_),
    .X(_058_));
 sky130_fd_sc_hd__or2_1 _460_ (.A(_386_),
    .B(_053_),
    .X(_059_));
 sky130_fd_sc_hd__or4_1 _461_ (.A(_380_),
    .B(_378_),
    .C(_381_),
    .D(_397_),
    .X(_060_));
 sky130_fd_sc_hd__nand2_1 _462_ (.A(_051_),
    .B(_060_),
    .Y(_061_));
 sky130_fd_sc_hd__a21o_1 _463_ (.A1(_058_),
    .A2(_059_),
    .B1(_061_),
    .X(_062_));
 sky130_fd_sc_hd__a41o_1 _464_ (.A1(_402_),
    .A2(_043_),
    .A3(_055_),
    .A4(_062_),
    .B1(_375_),
    .X(_063_));
 sky130_fd_sc_hd__a31o_1 _465_ (.A1(_049_),
    .A2(_403_),
    .A3(_039_),
    .B1(_033_),
    .X(_064_));
 sky130_fd_sc_hd__a21o_1 _466_ (.A1(_386_),
    .A2(_064_),
    .B1(_375_),
    .X(_065_));
 sky130_fd_sc_hd__and3_1 _467_ (.A(_390_),
    .B(_063_),
    .C(_065_),
    .X(_066_));
 sky130_fd_sc_hd__clkbuf_4 _468_ (.A(_066_),
    .X(_067_));
 sky130_fd_sc_hd__or2_1 _469_ (.A(_007_),
    .B(_389_),
    .X(_068_));
 sky130_fd_sc_hd__a41oi_4 _470_ (.A1(_402_),
    .A2(_043_),
    .A3(_055_),
    .A4(_062_),
    .B1(_375_),
    .Y(_069_));
 sky130_fd_sc_hd__clkbuf_4 _471_ (.A(\lcd.seq[0] ),
    .X(_070_));
 sky130_fd_sc_hd__inv_2 _472_ (.A(\lcd.rom_addr[0] ),
    .Y(_071_));
 sky130_fd_sc_hd__nand2_1 _473_ (.A(_070_),
    .B(_071_),
    .Y(_072_));
 sky130_fd_sc_hd__nor2_1 _474_ (.A(\lcd.rom_addr[1] ),
    .B(_072_),
    .Y(_073_));
 sky130_fd_sc_hd__or4b_1 _475_ (.A(net11),
    .B(_068_),
    .C(_069_),
    .D_N(_073_),
    .X(_074_));
 sky130_fd_sc_hd__buf_4 _476_ (.A(_074_),
    .X(_075_));
 sky130_fd_sc_hd__xnor2_4 _477_ (.A(\lcd.rom_addr[3] ),
    .B(_075_),
    .Y(_076_));
 sky130_fd_sc_hd__nor2_2 _478_ (.A(_067_),
    .B(_076_),
    .Y(_077_));
 sky130_fd_sc_hd__inv_2 _479_ (.A(_077_),
    .Y(_078_));
 sky130_fd_sc_hd__clkbuf_4 _480_ (.A(_078_),
    .X(_019_));
 sky130_fd_sc_hd__clkinv_2 _481_ (.A(_070_),
    .Y(_079_));
 sky130_fd_sc_hd__buf_2 _482_ (.A(_068_),
    .X(_080_));
 sky130_fd_sc_hd__o31a_2 _483_ (.A1(_079_),
    .A2(_080_),
    .A3(_069_),
    .B1(\lcd.rom_addr[0] ),
    .X(_081_));
 sky130_fd_sc_hd__nor2_1 _484_ (.A(_079_),
    .B(\lcd.rom_addr[0] ),
    .Y(_082_));
 sky130_fd_sc_hd__o211a_1 _485_ (.A1(_082_),
    .A2(_065_),
    .B1(_390_),
    .C1(_063_),
    .X(_083_));
 sky130_fd_sc_hd__or3_2 _486_ (.A(\lcd.rom_addr[1] ),
    .B(_081_),
    .C(_083_),
    .X(_084_));
 sky130_fd_sc_hd__inv_2 _487_ (.A(net11),
    .Y(_085_));
 sky130_fd_sc_hd__a31o_1 _488_ (.A1(_390_),
    .A2(_063_),
    .A3(_073_),
    .B1(_085_),
    .X(_086_));
 sky130_fd_sc_hd__a21o_2 _489_ (.A1(_075_),
    .A2(_086_),
    .B1(_066_),
    .X(_087_));
 sky130_fd_sc_hd__nand2_2 _490_ (.A(_084_),
    .B(_087_),
    .Y(_088_));
 sky130_fd_sc_hd__and3_1 _491_ (.A(_390_),
    .B(_063_),
    .C(_082_),
    .X(_089_));
 sky130_fd_sc_hd__or4_4 _492_ (.A(_085_),
    .B(_089_),
    .C(_066_),
    .D(_081_),
    .X(_090_));
 sky130_fd_sc_hd__or2_2 _493_ (.A(\lcd.rom_addr[1] ),
    .B(_090_),
    .X(_091_));
 sky130_fd_sc_hd__inv_2 _494_ (.A(\lcd.rom_addr[1] ),
    .Y(_092_));
 sky130_fd_sc_hd__a31o_1 _495_ (.A1(_070_),
    .A2(_390_),
    .A3(_063_),
    .B1(_071_),
    .X(_093_));
 sky130_fd_sc_hd__a21oi_1 _496_ (.A1(_386_),
    .A2(_064_),
    .B1(_375_),
    .Y(_094_));
 sky130_fd_sc_hd__a211o_1 _497_ (.A1(_072_),
    .A2(_094_),
    .B1(_080_),
    .C1(_069_),
    .X(_095_));
 sky130_fd_sc_hd__and3_1 _498_ (.A(_092_),
    .B(_093_),
    .C(_095_),
    .X(_096_));
 sky130_fd_sc_hd__o31a_1 _499_ (.A1(_080_),
    .A2(_069_),
    .A3(_072_),
    .B1(\lcd.rom_addr[1] ),
    .X(_097_));
 sky130_fd_sc_hd__o211a_1 _500_ (.A1(_073_),
    .A2(_065_),
    .B1(_390_),
    .C1(_063_),
    .X(_098_));
 sky130_fd_sc_hd__o22a_2 _501_ (.A1(_081_),
    .A2(_083_),
    .B1(_097_),
    .B2(_098_),
    .X(_099_));
 sky130_fd_sc_hd__nor2_1 _502_ (.A(_096_),
    .B(_099_),
    .Y(_100_));
 sky130_fd_sc_hd__a31o_1 _503_ (.A1(\lcd.rom_addr[3] ),
    .A2(_075_),
    .A3(_086_),
    .B1(_067_),
    .X(_101_));
 sky130_fd_sc_hd__nor3_1 _504_ (.A(\lcd.rom_addr[3] ),
    .B(\lcd.rom_addr[4] ),
    .C(_075_),
    .Y(_102_));
 sky130_fd_sc_hd__o21a_1 _505_ (.A1(\lcd.rom_addr[3] ),
    .A2(_075_),
    .B1(\lcd.rom_addr[4] ),
    .X(_103_));
 sky130_fd_sc_hd__nor3_2 _506_ (.A(_102_),
    .B(_067_),
    .C(_103_),
    .Y(_104_));
 sky130_fd_sc_hd__buf_2 _507_ (.A(_104_),
    .X(_105_));
 sky130_fd_sc_hd__a21oi_1 _508_ (.A1(_100_),
    .A2(_101_),
    .B1(_105_),
    .Y(_106_));
 sky130_fd_sc_hd__o211ai_1 _509_ (.A1(_019_),
    .A2(_088_),
    .B1(_091_),
    .C1(_106_),
    .Y(_107_));
 sky130_fd_sc_hd__or3_2 _510_ (.A(_080_),
    .B(_069_),
    .C(_094_),
    .X(_108_));
 sky130_fd_sc_hd__or4_1 _511_ (.A(\lcd.rom_addr[3] ),
    .B(\lcd.rom_addr[4] ),
    .C(\lcd.rom_addr[5] ),
    .D(_075_),
    .X(_109_));
 sky130_fd_sc_hd__or2b_1 _512_ (.A(_102_),
    .B_N(\lcd.rom_addr[5] ),
    .X(_110_));
 sky130_fd_sc_hd__and3_2 _513_ (.A(_108_),
    .B(_109_),
    .C(_110_),
    .X(_111_));
 sky130_fd_sc_hd__inv_2 _514_ (.A(_111_),
    .Y(_112_));
 sky130_fd_sc_hd__clkbuf_4 _515_ (.A(_112_),
    .X(_021_));
 sky130_fd_sc_hd__nor2_2 _516_ (.A(_097_),
    .B(_098_),
    .Y(_113_));
 sky130_fd_sc_hd__inv_2 _517_ (.A(_087_),
    .Y(_114_));
 sky130_fd_sc_hd__clkbuf_4 _518_ (.A(_114_),
    .X(_018_));
 sky130_fd_sc_hd__o22a_1 _519_ (.A1(_113_),
    .A2(_018_),
    .B1(_076_),
    .B2(_067_),
    .X(_115_));
 sky130_fd_sc_hd__or3_1 _520_ (.A(_092_),
    .B(_081_),
    .C(_083_),
    .X(_116_));
 sky130_fd_sc_hd__buf_2 _521_ (.A(_116_),
    .X(_117_));
 sky130_fd_sc_hd__or2_1 _522_ (.A(net11),
    .B(_117_),
    .X(_118_));
 sky130_fd_sc_hd__clkbuf_2 _523_ (.A(_118_),
    .X(_119_));
 sky130_fd_sc_hd__or3_2 _524_ (.A(_085_),
    .B(_097_),
    .C(_098_),
    .X(_120_));
 sky130_fd_sc_hd__inv_2 _525_ (.A(_104_),
    .Y(_121_));
 sky130_fd_sc_hd__a31o_1 _526_ (.A1(_077_),
    .A2(_119_),
    .A3(_120_),
    .B1(_121_),
    .X(_122_));
 sky130_fd_sc_hd__a21o_1 _527_ (.A1(_100_),
    .A2(_115_),
    .B1(_122_),
    .X(_123_));
 sky130_fd_sc_hd__nor2_1 _528_ (.A(_077_),
    .B(_119_),
    .Y(_124_));
 sky130_fd_sc_hd__a2bb2o_2 _529_ (.A1_N(_098_),
    .A2_N(_097_),
    .B1(_095_),
    .B2(_093_),
    .X(_125_));
 sky130_fd_sc_hd__or4_4 _530_ (.A(net11),
    .B(_089_),
    .C(_067_),
    .D(_081_),
    .X(_126_));
 sky130_fd_sc_hd__and4_1 _531_ (.A(_125_),
    .B(_077_),
    .C(_126_),
    .D(_120_),
    .X(_127_));
 sky130_fd_sc_hd__nand2_1 _532_ (.A(_117_),
    .B(_114_),
    .Y(_128_));
 sky130_fd_sc_hd__xor2_4 _533_ (.A(\lcd.rom_addr[3] ),
    .B(_075_),
    .X(_129_));
 sky130_fd_sc_hd__o311a_1 _534_ (.A1(_096_),
    .A2(_099_),
    .A3(_114_),
    .B1(_129_),
    .C1(_108_),
    .X(_130_));
 sky130_fd_sc_hd__o211a_1 _535_ (.A1(_067_),
    .A2(_076_),
    .B1(_090_),
    .C1(_084_),
    .X(_131_));
 sky130_fd_sc_hd__buf_2 _536_ (.A(_121_),
    .X(_132_));
 sky130_fd_sc_hd__a211o_1 _537_ (.A1(_128_),
    .A2(_130_),
    .B1(_131_),
    .C1(_132_),
    .X(_133_));
 sky130_fd_sc_hd__o311a_1 _538_ (.A1(_105_),
    .A2(_124_),
    .A3(_127_),
    .B1(_111_),
    .C1(_133_),
    .X(_134_));
 sky130_fd_sc_hd__a31o_1 _539_ (.A1(_107_),
    .A2(_021_),
    .A3(_123_),
    .B1(_134_),
    .X(_135_));
 sky130_fd_sc_hd__buf_2 _540_ (.A(_078_),
    .X(_136_));
 sky130_fd_sc_hd__nor2_1 _541_ (.A(_099_),
    .B(_136_),
    .Y(_137_));
 sky130_fd_sc_hd__a221o_1 _542_ (.A1(_126_),
    .A2(_115_),
    .B1(_137_),
    .B2(_088_),
    .C1(_105_),
    .X(_138_));
 sky130_fd_sc_hd__o21a_1 _543_ (.A1(_067_),
    .A2(_076_),
    .B1(_120_),
    .X(_139_));
 sky130_fd_sc_hd__nor2_2 _544_ (.A(_081_),
    .B(_083_),
    .Y(_140_));
 sky130_fd_sc_hd__clkinv_2 _545_ (.A(_140_),
    .Y(_016_));
 sky130_fd_sc_hd__and4_1 _546_ (.A(_108_),
    .B(_016_),
    .C(_129_),
    .D(_120_),
    .X(_141_));
 sky130_fd_sc_hd__a211o_1 _547_ (.A1(_125_),
    .A2(_139_),
    .B1(_141_),
    .C1(_121_),
    .X(_142_));
 sky130_fd_sc_hd__and2_1 _548_ (.A(_112_),
    .B(_142_),
    .X(_143_));
 sky130_fd_sc_hd__or3_1 _549_ (.A(_080_),
    .B(_069_),
    .C(_072_),
    .X(_144_));
 sky130_fd_sc_hd__and3_1 _550_ (.A(_390_),
    .B(_063_),
    .C(_073_),
    .X(_145_));
 sky130_fd_sc_hd__a2111o_1 _551_ (.A1(_144_),
    .A2(_093_),
    .B1(_097_),
    .C1(_145_),
    .D1(_066_),
    .X(_146_));
 sky130_fd_sc_hd__nor2_1 _552_ (.A(_146_),
    .B(_114_),
    .Y(_147_));
 sky130_fd_sc_hd__and2_1 _553_ (.A(_146_),
    .B(_114_),
    .X(_148_));
 sky130_fd_sc_hd__o211a_1 _554_ (.A1(_147_),
    .A2(_148_),
    .B1(_117_),
    .C1(_076_),
    .X(_149_));
 sky130_fd_sc_hd__a21o_1 _555_ (.A1(_084_),
    .A2(_125_),
    .B1(_087_),
    .X(_150_));
 sky130_fd_sc_hd__a21o_1 _556_ (.A1(_150_),
    .A2(_130_),
    .B1(_121_),
    .X(_151_));
 sky130_fd_sc_hd__o211a_1 _557_ (.A1(_125_),
    .A2(_018_),
    .B1(_077_),
    .C1(_084_),
    .X(_152_));
 sky130_fd_sc_hd__nand2_1 _558_ (.A(_146_),
    .B(_018_),
    .Y(_153_));
 sky130_fd_sc_hd__a31o_1 _559_ (.A1(_078_),
    .A2(_126_),
    .A3(_153_),
    .B1(_105_),
    .X(_154_));
 sky130_fd_sc_hd__o22a_1 _560_ (.A1(_149_),
    .A2(_151_),
    .B1(_152_),
    .B2(_154_),
    .X(_155_));
 sky130_fd_sc_hd__a22o_1 _561_ (.A1(_138_),
    .A2(_143_),
    .B1(_155_),
    .B2(_111_),
    .X(_156_));
 sky130_fd_sc_hd__nor2_1 _562_ (.A(\lcd.rom_addr[6] ),
    .B(_109_),
    .Y(_157_));
 sky130_fd_sc_hd__a211o_1 _563_ (.A1(\lcd.rom_addr[6] ),
    .A2(_109_),
    .B1(_157_),
    .C1(_067_),
    .X(_158_));
 sky130_fd_sc_hd__clkbuf_4 _564_ (.A(_158_),
    .X(_022_));
 sky130_fd_sc_hd__mux2_1 _565_ (.A0(_135_),
    .A1(_156_),
    .S(_022_),
    .X(_159_));
 sky130_fd_sc_hd__clkbuf_1 _566_ (.A(_159_),
    .X(_000_));
 sky130_fd_sc_hd__buf_2 _567_ (.A(_111_),
    .X(_160_));
 sky130_fd_sc_hd__clkinv_2 _568_ (.A(_022_),
    .Y(_161_));
 sky130_fd_sc_hd__buf_2 _569_ (.A(_077_),
    .X(_162_));
 sky130_fd_sc_hd__and3_1 _570_ (.A(_162_),
    .B(_088_),
    .C(_153_),
    .X(_163_));
 sky130_fd_sc_hd__and2_1 _571_ (.A(_117_),
    .B(_087_),
    .X(_164_));
 sky130_fd_sc_hd__clkbuf_4 _572_ (.A(_105_),
    .X(_165_));
 sky130_fd_sc_hd__a21o_1 _573_ (.A1(_136_),
    .A2(_164_),
    .B1(_165_),
    .X(_166_));
 sky130_fd_sc_hd__buf_2 _574_ (.A(_132_),
    .X(_167_));
 sky130_fd_sc_hd__a21o_1 _575_ (.A1(_128_),
    .A2(_130_),
    .B1(_167_),
    .X(_168_));
 sky130_fd_sc_hd__o21ai_1 _576_ (.A1(_163_),
    .A2(_166_),
    .B1(_168_),
    .Y(_169_));
 sky130_fd_sc_hd__or3_1 _577_ (.A(_132_),
    .B(_129_),
    .C(_119_),
    .X(_170_));
 sky130_fd_sc_hd__o32a_1 _578_ (.A1(_100_),
    .A2(_018_),
    .A3(_162_),
    .B1(_090_),
    .B2(_076_),
    .X(_171_));
 sky130_fd_sc_hd__a311o_1 _579_ (.A1(_136_),
    .A2(_119_),
    .A3(_150_),
    .B1(_141_),
    .C1(_105_),
    .X(_172_));
 sky130_fd_sc_hd__o211a_1 _580_ (.A1(_167_),
    .A2(_171_),
    .B1(_172_),
    .C1(_022_),
    .X(_173_));
 sky130_fd_sc_hd__a31o_1 _581_ (.A1(_161_),
    .A2(_169_),
    .A3(_170_),
    .B1(_173_),
    .X(_174_));
 sky130_fd_sc_hd__buf_2 _582_ (.A(_132_),
    .X(_020_));
 sky130_fd_sc_hd__nand2_1 _583_ (.A(_020_),
    .B(_126_),
    .Y(_175_));
 sky130_fd_sc_hd__inv_2 _584_ (.A(_113_),
    .Y(_017_));
 sky130_fd_sc_hd__a31o_1 _585_ (.A1(_019_),
    .A2(_090_),
    .A3(_088_),
    .B1(_167_),
    .X(_176_));
 sky130_fd_sc_hd__a31o_1 _586_ (.A1(_017_),
    .A2(_162_),
    .A3(_126_),
    .B1(_176_),
    .X(_177_));
 sky130_fd_sc_hd__o211ai_1 _587_ (.A1(_115_),
    .A2(_175_),
    .B1(_177_),
    .C1(_161_),
    .Y(_178_));
 sky130_fd_sc_hd__nor2_1 _588_ (.A(_087_),
    .B(_129_),
    .Y(_179_));
 sky130_fd_sc_hd__or2_1 _589_ (.A(_105_),
    .B(_179_),
    .X(_180_));
 sky130_fd_sc_hd__a221o_1 _590_ (.A1(_120_),
    .A2(_130_),
    .B1(_153_),
    .B2(_136_),
    .C1(_167_),
    .X(_181_));
 sky130_fd_sc_hd__o211a_1 _591_ (.A1(_163_),
    .A2(_180_),
    .B1(_181_),
    .C1(_022_),
    .X(_182_));
 sky130_fd_sc_hd__nor2_1 _592_ (.A(_160_),
    .B(_182_),
    .Y(_183_));
 sky130_fd_sc_hd__a22oi_1 _593_ (.A1(_160_),
    .A2(_174_),
    .B1(_178_),
    .B2(_183_),
    .Y(_001_));
 sky130_fd_sc_hd__o211a_1 _594_ (.A1(_146_),
    .A2(_018_),
    .B1(_129_),
    .C1(_108_),
    .X(_184_));
 sky130_fd_sc_hd__a221o_1 _595_ (.A1(_090_),
    .A2(_115_),
    .B1(_184_),
    .B2(_091_),
    .C1(_020_),
    .X(_185_));
 sky130_fd_sc_hd__a211oi_1 _596_ (.A1(_126_),
    .A2(_120_),
    .B1(_067_),
    .C1(_076_),
    .Y(_186_));
 sky130_fd_sc_hd__a211o_1 _597_ (.A1(_019_),
    .A2(_088_),
    .B1(_186_),
    .C1(_165_),
    .X(_187_));
 sky130_fd_sc_hd__nand2_1 _598_ (.A(_085_),
    .B(_113_),
    .Y(_188_));
 sky130_fd_sc_hd__and3_1 _599_ (.A(_117_),
    .B(_136_),
    .C(_188_),
    .X(_189_));
 sky130_fd_sc_hd__xnor2_1 _600_ (.A(_113_),
    .B(_018_),
    .Y(_190_));
 sky130_fd_sc_hd__o22a_1 _601_ (.A1(_140_),
    .A2(_018_),
    .B1(_076_),
    .B2(_067_),
    .X(_191_));
 sky130_fd_sc_hd__a211o_1 _602_ (.A1(_162_),
    .A2(_190_),
    .B1(_191_),
    .C1(_165_),
    .X(_192_));
 sky130_fd_sc_hd__o211a_1 _603_ (.A1(_122_),
    .A2(_189_),
    .B1(_192_),
    .C1(_160_),
    .X(_193_));
 sky130_fd_sc_hd__a31o_1 _604_ (.A1(_021_),
    .A2(_185_),
    .A3(_187_),
    .B1(_193_),
    .X(_194_));
 sky130_fd_sc_hd__o21a_1 _605_ (.A1(_100_),
    .A2(_018_),
    .B1(_139_),
    .X(_195_));
 sky130_fd_sc_hd__o21a_1 _606_ (.A1(_147_),
    .A2(_148_),
    .B1(_162_),
    .X(_196_));
 sky130_fd_sc_hd__nor2_1 _607_ (.A(_092_),
    .B(_016_),
    .Y(_197_));
 sky130_fd_sc_hd__nor4_1 _608_ (.A(_197_),
    .B(_162_),
    .C(_147_),
    .D(_148_),
    .Y(_198_));
 sky130_fd_sc_hd__nand2_1 _609_ (.A(_084_),
    .B(_018_),
    .Y(_199_));
 sky130_fd_sc_hd__a31o_1 _610_ (.A1(_162_),
    .A2(_126_),
    .A3(_199_),
    .B1(_132_),
    .X(_200_));
 sky130_fd_sc_hd__o32a_1 _611_ (.A1(_165_),
    .A2(_195_),
    .A3(_196_),
    .B1(_198_),
    .B2(_200_),
    .X(_201_));
 sky130_fd_sc_hd__o211a_1 _612_ (.A1(_147_),
    .A2(_148_),
    .B1(_117_),
    .C1(_162_),
    .X(_202_));
 sky130_fd_sc_hd__a21o_1 _613_ (.A1(_136_),
    .A2(_128_),
    .B1(_132_),
    .X(_203_));
 sky130_fd_sc_hd__or3_1 _614_ (.A(_105_),
    .B(_139_),
    .C(_186_),
    .X(_204_));
 sky130_fd_sc_hd__o211a_1 _615_ (.A1(_202_),
    .A2(_203_),
    .B1(_204_),
    .C1(_160_),
    .X(_205_));
 sky130_fd_sc_hd__a211o_1 _616_ (.A1(_021_),
    .A2(_201_),
    .B1(_205_),
    .C1(_022_),
    .X(_206_));
 sky130_fd_sc_hd__o21a_1 _617_ (.A1(_161_),
    .A2(_194_),
    .B1(_206_),
    .X(_002_));
 sky130_fd_sc_hd__and3_1 _618_ (.A(_016_),
    .B(_114_),
    .C(_129_),
    .X(_207_));
 sky130_fd_sc_hd__a31o_1 _619_ (.A1(_117_),
    .A2(_120_),
    .A3(_191_),
    .B1(_207_),
    .X(_208_));
 sky130_fd_sc_hd__a21boi_1 _620_ (.A1(_020_),
    .A2(_208_),
    .B1_N(_170_),
    .Y(_209_));
 sky130_fd_sc_hd__a31o_1 _621_ (.A1(_125_),
    .A2(_019_),
    .A3(_199_),
    .B1(_207_),
    .X(_210_));
 sky130_fd_sc_hd__a22o_1 _622_ (.A1(_016_),
    .A2(_087_),
    .B1(_129_),
    .B2(_108_),
    .X(_211_));
 sky130_fd_sc_hd__and4_1 _623_ (.A(_132_),
    .B(_090_),
    .C(_188_),
    .D(_211_),
    .X(_212_));
 sky130_fd_sc_hd__a211o_1 _624_ (.A1(_165_),
    .A2(_210_),
    .B1(_212_),
    .C1(_160_),
    .X(_213_));
 sky130_fd_sc_hd__o21ai_1 _625_ (.A1(_021_),
    .A2(_209_),
    .B1(_213_),
    .Y(_214_));
 sky130_fd_sc_hd__a21oi_1 _626_ (.A1(_119_),
    .A2(_150_),
    .B1(_019_),
    .Y(_215_));
 sky130_fd_sc_hd__a211o_1 _627_ (.A1(_019_),
    .A2(_147_),
    .B1(_215_),
    .C1(_165_),
    .X(_216_));
 sky130_fd_sc_hd__a211o_1 _628_ (.A1(_140_),
    .A2(_139_),
    .B1(_141_),
    .C1(_167_),
    .X(_217_));
 sky130_fd_sc_hd__and3_1 _629_ (.A(_021_),
    .B(_216_),
    .C(_217_),
    .X(_218_));
 sky130_fd_sc_hd__nand2_1 _630_ (.A(_113_),
    .B(_207_),
    .Y(_219_));
 sky130_fd_sc_hd__nand3_1 _631_ (.A(_020_),
    .B(_188_),
    .C(_219_),
    .Y(_220_));
 sky130_fd_sc_hd__a2111o_1 _632_ (.A1(_099_),
    .A2(_179_),
    .B1(_202_),
    .C1(_124_),
    .D1(_167_),
    .X(_221_));
 sky130_fd_sc_hd__a31o_1 _633_ (.A1(_160_),
    .A2(_220_),
    .A3(_221_),
    .B1(_022_),
    .X(_222_));
 sky130_fd_sc_hd__o22a_1 _634_ (.A1(_161_),
    .A2(_214_),
    .B1(_218_),
    .B2(_222_),
    .X(_003_));
 sky130_fd_sc_hd__o21ai_1 _635_ (.A1(_096_),
    .A2(_191_),
    .B1(_091_),
    .Y(_223_));
 sky130_fd_sc_hd__nand2_1 _636_ (.A(_020_),
    .B(_223_),
    .Y(_224_));
 sky130_fd_sc_hd__nor2_1 _637_ (.A(_016_),
    .B(_087_),
    .Y(_225_));
 sky130_fd_sc_hd__and2_1 _638_ (.A(_099_),
    .B(_101_),
    .X(_226_));
 sky130_fd_sc_hd__a211o_1 _639_ (.A1(_129_),
    .A2(_225_),
    .B1(_226_),
    .C1(_020_),
    .X(_227_));
 sky130_fd_sc_hd__a221o_1 _640_ (.A1(_140_),
    .A2(_087_),
    .B1(_129_),
    .B2(_108_),
    .C1(_113_),
    .X(_228_));
 sky130_fd_sc_hd__o211a_1 _641_ (.A1(_019_),
    .A2(_119_),
    .B1(_228_),
    .C1(_167_),
    .X(_229_));
 sky130_fd_sc_hd__o2111a_1 _642_ (.A1(_125_),
    .A2(_101_),
    .B1(_090_),
    .C1(_188_),
    .D1(_165_),
    .X(_230_));
 sky130_fd_sc_hd__nor3_1 _643_ (.A(_021_),
    .B(_229_),
    .C(_230_),
    .Y(_231_));
 sky130_fd_sc_hd__a31o_1 _644_ (.A1(_021_),
    .A2(_224_),
    .A3(_227_),
    .B1(_231_),
    .X(_232_));
 sky130_fd_sc_hd__nand2_1 _645_ (.A(_117_),
    .B(_087_),
    .Y(_233_));
 sky130_fd_sc_hd__a32o_1 _646_ (.A1(_019_),
    .A2(_233_),
    .A3(_199_),
    .B1(_184_),
    .B2(_128_),
    .X(_234_));
 sky130_fd_sc_hd__nor2_1 _647_ (.A(_020_),
    .B(_171_),
    .Y(_235_));
 sky130_fd_sc_hd__a211o_1 _648_ (.A1(_020_),
    .A2(_234_),
    .B1(_235_),
    .C1(_021_),
    .X(_236_));
 sky130_fd_sc_hd__nor2_1 _649_ (.A(_136_),
    .B(_119_),
    .Y(_237_));
 sky130_fd_sc_hd__o32a_1 _650_ (.A1(_167_),
    .A2(_101_),
    .A3(_207_),
    .B1(_237_),
    .B2(_180_),
    .X(_238_));
 sky130_fd_sc_hd__o21a_1 _651_ (.A1(_160_),
    .A2(_238_),
    .B1(_022_),
    .X(_239_));
 sky130_fd_sc_hd__a22o_1 _652_ (.A1(_161_),
    .A2(_232_),
    .B1(_236_),
    .B2(_239_),
    .X(_004_));
 sky130_fd_sc_hd__a211o_1 _653_ (.A1(_019_),
    .A2(_164_),
    .B1(_148_),
    .C1(_167_),
    .X(_240_));
 sky130_fd_sc_hd__a31o_1 _654_ (.A1(_017_),
    .A2(_162_),
    .A3(_225_),
    .B1(_226_),
    .X(_241_));
 sky130_fd_sc_hd__a2bb2o_1 _655_ (.A1_N(_184_),
    .A2_N(_240_),
    .B1(_241_),
    .B2(_020_),
    .X(_242_));
 sky130_fd_sc_hd__nand2_1 _656_ (.A(_160_),
    .B(_242_),
    .Y(_243_));
 sky130_fd_sc_hd__or3_1 _657_ (.A(_117_),
    .B(_160_),
    .C(_180_),
    .X(_244_));
 sky130_fd_sc_hd__a21o_1 _658_ (.A1(_197_),
    .A2(_179_),
    .B1(_132_),
    .X(_245_));
 sky130_fd_sc_hd__o311a_1 _659_ (.A1(_165_),
    .A2(_237_),
    .A3(_226_),
    .B1(_245_),
    .C1(_160_),
    .X(_246_));
 sky130_fd_sc_hd__a2111o_1 _660_ (.A1(_125_),
    .A2(_136_),
    .B1(_101_),
    .C1(_184_),
    .D1(_132_),
    .X(_247_));
 sky130_fd_sc_hd__a221o_1 _661_ (.A1(_162_),
    .A2(_091_),
    .B1(_139_),
    .B2(_117_),
    .C1(_105_),
    .X(_248_));
 sky130_fd_sc_hd__a21o_1 _662_ (.A1(_247_),
    .A2(_248_),
    .B1(_111_),
    .X(_249_));
 sky130_fd_sc_hd__and3b_1 _663_ (.A_N(_246_),
    .B(_161_),
    .C(_249_),
    .X(_250_));
 sky130_fd_sc_hd__a31o_1 _664_ (.A1(_022_),
    .A2(_243_),
    .A3(_244_),
    .B1(_250_),
    .X(_005_));
 sky130_fd_sc_hd__inv_2 _665_ (.A(_226_),
    .Y(_251_));
 sky130_fd_sc_hd__or3_1 _666_ (.A(_078_),
    .B(_148_),
    .C(_164_),
    .X(_252_));
 sky130_fd_sc_hd__o21a_1 _667_ (.A1(_077_),
    .A2(_091_),
    .B1(_104_),
    .X(_253_));
 sky130_fd_sc_hd__a32o_1 _668_ (.A1(_132_),
    .A2(_219_),
    .A3(_251_),
    .B1(_252_),
    .B2(_253_),
    .X(_254_));
 sky130_fd_sc_hd__o21a_1 _669_ (.A1(_137_),
    .A2(_139_),
    .B1(_167_),
    .X(_255_));
 sky130_fd_sc_hd__a21o_1 _670_ (.A1(_165_),
    .A2(_076_),
    .B1(_112_),
    .X(_256_));
 sky130_fd_sc_hd__o22a_1 _671_ (.A1(_111_),
    .A2(_254_),
    .B1(_255_),
    .B2(_256_),
    .X(_257_));
 sky130_fd_sc_hd__a21o_1 _672_ (.A1(_017_),
    .A2(_225_),
    .B1(_136_),
    .X(_258_));
 sky130_fd_sc_hd__nand2_1 _673_ (.A(_091_),
    .B(_115_),
    .Y(_259_));
 sky130_fd_sc_hd__a21o_1 _674_ (.A1(_016_),
    .A2(_188_),
    .B1(_136_),
    .X(_260_));
 sky130_fd_sc_hd__a32o_1 _675_ (.A1(_165_),
    .A2(_258_),
    .A3(_259_),
    .B1(_260_),
    .B2(_106_),
    .X(_261_));
 sky130_fd_sc_hd__a21o_1 _676_ (.A1(_099_),
    .A2(_179_),
    .B1(_105_),
    .X(_262_));
 sky130_fd_sc_hd__o211a_1 _677_ (.A1(_237_),
    .A2(_245_),
    .B1(_262_),
    .C1(_111_),
    .X(_263_));
 sky130_fd_sc_hd__a21oi_1 _678_ (.A1(_021_),
    .A2(_261_),
    .B1(_263_),
    .Y(_264_));
 sky130_fd_sc_hd__mux2_1 _679_ (.A0(_257_),
    .A1(_264_),
    .S(_022_),
    .X(_265_));
 sky130_fd_sc_hd__clkbuf_1 _680_ (.A(_265_),
    .X(_006_));
 sky130_fd_sc_hd__or2_1 _681_ (.A(net1),
    .B(net3),
    .X(_266_));
 sky130_fd_sc_hd__nand2_1 _682_ (.A(net1),
    .B(net3),
    .Y(_267_));
 sky130_fd_sc_hd__nand2_1 _683_ (.A(_266_),
    .B(_267_),
    .Y(_268_));
 sky130_fd_sc_hd__xnor2_1 _684_ (.A(net2),
    .B(_268_),
    .Y(_009_));
 sky130_fd_sc_hd__a21bo_1 _685_ (.A1(net2),
    .A2(_266_),
    .B1_N(_267_),
    .X(_008_));
 sky130_fd_sc_hd__nor3_2 _686_ (.A(_041_),
    .B(_397_),
    .C(_037_),
    .Y(_269_));
 sky130_fd_sc_hd__mux2_2 _687_ (.A0(\lcd.s_ROM[4] ),
    .A1(\lcd.s_ROM[0] ),
    .S(_070_),
    .X(_270_));
 sky130_fd_sc_hd__buf_2 _688_ (.A(_070_),
    .X(_271_));
 sky130_fd_sc_hd__a22o_1 _689_ (.A1(_079_),
    .A2(_045_),
    .B1(_053_),
    .B2(_399_),
    .X(_272_));
 sky130_fd_sc_hd__nor2_1 _690_ (.A(_045_),
    .B(_048_),
    .Y(_273_));
 sky130_fd_sc_hd__nand2_1 _691_ (.A(_399_),
    .B(_273_),
    .Y(_274_));
 sky130_fd_sc_hd__a21oi_2 _692_ (.A1(_049_),
    .A2(_403_),
    .B1(_033_),
    .Y(_275_));
 sky130_fd_sc_hd__nand2_1 _693_ (.A(_275_),
    .B(_057_),
    .Y(_276_));
 sky130_fd_sc_hd__o21a_1 _694_ (.A1(_270_),
    .A2(_274_),
    .B1(_276_),
    .X(_277_));
 sky130_fd_sc_hd__a2bb2o_1 _695_ (.A1_N(_271_),
    .A2_N(_053_),
    .B1(_272_),
    .B2(_277_),
    .X(_278_));
 sky130_fd_sc_hd__or2b_2 _696_ (.A(\lcd.round[1] ),
    .B_N(\lcd.round[0] ),
    .X(_279_));
 sky130_fd_sc_hd__a221o_1 _697_ (.A1(_269_),
    .A2(_270_),
    .B1(_278_),
    .B2(_054_),
    .C1(_279_),
    .X(_280_));
 sky130_fd_sc_hd__and3_1 _698_ (.A(_041_),
    .B(_049_),
    .C(_039_),
    .X(_281_));
 sky130_fd_sc_hd__nor2_1 _699_ (.A(_037_),
    .B(_281_),
    .Y(_282_));
 sky130_fd_sc_hd__a31o_1 _700_ (.A1(_079_),
    .A2(_382_),
    .A3(_281_),
    .B1(_051_),
    .X(_283_));
 sky130_fd_sc_hd__buf_2 _701_ (.A(\lcd.seq[1] ),
    .X(_284_));
 sky130_fd_sc_hd__o22a_1 _702_ (.A1(\lcd.seq[1] ),
    .A2(\lcd.num_state[1] ),
    .B1(\lcd.num_state[0] ),
    .B2(_052_),
    .X(_285_));
 sky130_fd_sc_hd__o221a_1 _703_ (.A1(_052_),
    .A2(_284_),
    .B1(_079_),
    .B2(_285_),
    .C1(_403_),
    .X(_286_));
 sky130_fd_sc_hd__o21ai_1 _704_ (.A1(_041_),
    .A2(_398_),
    .B1(_381_),
    .Y(_287_));
 sky130_fd_sc_hd__a21bo_1 _705_ (.A1(_287_),
    .A2(_270_),
    .B1_N(_275_),
    .X(_288_));
 sky130_fd_sc_hd__o21a_1 _706_ (.A1(_286_),
    .A2(_288_),
    .B1(_037_),
    .X(_289_));
 sky130_fd_sc_hd__a211o_1 _707_ (.A1(_270_),
    .A2(_282_),
    .B1(_283_),
    .C1(_289_),
    .X(_290_));
 sky130_fd_sc_hd__and2_1 _708_ (.A(_386_),
    .B(_396_),
    .X(_291_));
 sky130_fd_sc_hd__o21a_1 _709_ (.A1(_064_),
    .A2(_270_),
    .B1(_291_),
    .X(_292_));
 sky130_fd_sc_hd__a31o_1 _710_ (.A1(_401_),
    .A2(_280_),
    .A3(_290_),
    .B1(_292_),
    .X(_293_));
 sky130_fd_sc_hd__or2_1 _711_ (.A(_383_),
    .B(_293_),
    .X(_294_));
 sky130_fd_sc_hd__nor2_1 _712_ (.A(_052_),
    .B(_284_),
    .Y(_295_));
 sky130_fd_sc_hd__a21o_1 _713_ (.A1(_052_),
    .A2(_284_),
    .B1(_271_),
    .X(_296_));
 sky130_fd_sc_hd__or4_1 _714_ (.A(_376_),
    .B(_295_),
    .C(_060_),
    .D(_296_),
    .X(_297_));
 sky130_fd_sc_hd__nor3_1 _715_ (.A(_041_),
    .B(_052_),
    .C(_049_),
    .Y(_298_));
 sky130_fd_sc_hd__and3_1 _716_ (.A(_271_),
    .B(_382_),
    .C(_298_),
    .X(_299_));
 sky130_fd_sc_hd__mux2_1 _717_ (.A0(_297_),
    .A1(_284_),
    .S(_299_),
    .X(_300_));
 sky130_fd_sc_hd__nor2_1 _718_ (.A(_375_),
    .B(_389_),
    .Y(_301_));
 sky130_fd_sc_hd__a32o_1 _719_ (.A1(_294_),
    .A2(_300_),
    .A3(_301_),
    .B1(_080_),
    .B2(net12),
    .X(_010_));
 sky130_fd_sc_hd__inv_2 _720_ (.A(_034_),
    .Y(_302_));
 sky130_fd_sc_hd__mux2_2 _721_ (.A0(\lcd.s_ROM[5] ),
    .A1(\lcd.s_ROM[1] ),
    .S(_070_),
    .X(_303_));
 sky130_fd_sc_hd__a21o_1 _722_ (.A1(_377_),
    .A2(_403_),
    .B1(_033_),
    .X(_304_));
 sky130_fd_sc_hd__or3_1 _723_ (.A(_079_),
    .B(_034_),
    .C(_304_),
    .X(_305_));
 sky130_fd_sc_hd__a22o_1 _724_ (.A1(_282_),
    .A2(_303_),
    .B1(_305_),
    .B2(_037_),
    .X(_306_));
 sky130_fd_sc_hd__o2111a_1 _725_ (.A1(_302_),
    .A2(_303_),
    .B1(_306_),
    .C1(_279_),
    .D1(_401_),
    .X(_307_));
 sky130_fd_sc_hd__a21o_1 _726_ (.A1(_271_),
    .A2(_398_),
    .B1(_399_),
    .X(_308_));
 sky130_fd_sc_hd__a32o_1 _727_ (.A1(_053_),
    .A2(_276_),
    .A3(_308_),
    .B1(_303_),
    .B2(_269_),
    .X(_309_));
 sky130_fd_sc_hd__o211a_1 _728_ (.A1(_274_),
    .A2(_303_),
    .B1(_309_),
    .C1(_051_),
    .X(_310_));
 sky130_fd_sc_hd__o21a_1 _729_ (.A1(_064_),
    .A2(_303_),
    .B1(_291_),
    .X(_311_));
 sky130_fd_sc_hd__or4_1 _730_ (.A(_383_),
    .B(_307_),
    .C(_310_),
    .D(_311_),
    .X(_312_));
 sky130_fd_sc_hd__or4b_1 _731_ (.A(_041_),
    .B(_284_),
    .C(_049_),
    .D_N(_052_),
    .X(_313_));
 sky130_fd_sc_hd__or3_1 _732_ (.A(_079_),
    .B(_037_),
    .C(_313_),
    .X(_314_));
 sky130_fd_sc_hd__o211a_1 _733_ (.A1(_051_),
    .A2(_314_),
    .B1(_301_),
    .C1(_297_),
    .X(_315_));
 sky130_fd_sc_hd__a22o_1 _734_ (.A1(net8),
    .A2(_080_),
    .B1(_312_),
    .B2(_315_),
    .X(_011_));
 sky130_fd_sc_hd__a21oi_1 _735_ (.A1(_381_),
    .A2(_281_),
    .B1(_033_),
    .Y(_316_));
 sky130_fd_sc_hd__mux2_1 _736_ (.A0(\lcd.s_ROM[6] ),
    .A1(\lcd.s_ROM[2] ),
    .S(_070_),
    .X(_317_));
 sky130_fd_sc_hd__nor2_1 _737_ (.A(_271_),
    .B(_396_),
    .Y(_318_));
 sky130_fd_sc_hd__a31o_1 _738_ (.A1(_396_),
    .A2(_316_),
    .A3(_317_),
    .B1(_318_),
    .X(_319_));
 sky130_fd_sc_hd__and2_1 _739_ (.A(_386_),
    .B(_319_),
    .X(_320_));
 sky130_fd_sc_hd__nor2_1 _740_ (.A(_033_),
    .B(_056_),
    .Y(_321_));
 sky130_fd_sc_hd__a21boi_1 _741_ (.A1(_271_),
    .A2(_045_),
    .B1_N(_276_),
    .Y(_322_));
 sky130_fd_sc_hd__a41o_1 _742_ (.A1(_399_),
    .A2(_053_),
    .A3(_058_),
    .A4(_273_),
    .B1(_269_),
    .X(_323_));
 sky130_fd_sc_hd__a2bb2o_1 _743_ (.A1_N(_321_),
    .A2_N(_322_),
    .B1(_317_),
    .B2(_323_),
    .X(_324_));
 sky130_fd_sc_hd__a221o_1 _744_ (.A1(_382_),
    .A2(_281_),
    .B1(_317_),
    .B2(_034_),
    .C1(_051_),
    .X(_325_));
 sky130_fd_sc_hd__o211a_1 _745_ (.A1(_279_),
    .A2(_324_),
    .B1(_325_),
    .C1(_401_),
    .X(_326_));
 sky130_fd_sc_hd__or3_1 _746_ (.A(_383_),
    .B(_320_),
    .C(_326_),
    .X(_327_));
 sky130_fd_sc_hd__nand3b_1 _747_ (.A_N(_299_),
    .B(_297_),
    .C(_314_),
    .Y(_328_));
 sky130_fd_sc_hd__nand2_1 _748_ (.A(_284_),
    .B(_070_),
    .Y(_329_));
 sky130_fd_sc_hd__xnor2_1 _749_ (.A(_052_),
    .B(_329_),
    .Y(_330_));
 sky130_fd_sc_hd__a31o_1 _750_ (.A1(_284_),
    .A2(_279_),
    .A3(_299_),
    .B1(_042_),
    .X(_331_));
 sky130_fd_sc_hd__a31o_1 _751_ (.A1(_051_),
    .A2(_328_),
    .A3(_330_),
    .B1(_331_),
    .X(_332_));
 sky130_fd_sc_hd__a32o_1 _752_ (.A1(_301_),
    .A2(_327_),
    .A3(_332_),
    .B1(_080_),
    .B2(net9),
    .X(_012_));
 sky130_fd_sc_hd__nand2_1 _753_ (.A(_070_),
    .B(\lcd.s_ROM[3] ),
    .Y(_333_));
 sky130_fd_sc_hd__inv_2 _754_ (.A(_333_),
    .Y(_334_));
 sky130_fd_sc_hd__a31o_1 _755_ (.A1(_396_),
    .A2(_316_),
    .A3(_334_),
    .B1(_318_),
    .X(_335_));
 sky130_fd_sc_hd__nor2_1 _756_ (.A(_033_),
    .B(_057_),
    .Y(_336_));
 sky130_fd_sc_hd__o21bai_1 _757_ (.A1(_275_),
    .A2(_274_),
    .B1_N(_336_),
    .Y(_337_));
 sky130_fd_sc_hd__and2_1 _758_ (.A(_058_),
    .B(_334_),
    .X(_338_));
 sky130_fd_sc_hd__nor2_1 _759_ (.A(_045_),
    .B(_275_),
    .Y(_339_));
 sky130_fd_sc_hd__o41a_1 _760_ (.A1(_070_),
    .A2(_339_),
    .A3(_321_),
    .A4(_336_),
    .B1(_053_),
    .X(_340_));
 sky130_fd_sc_hd__a21bo_1 _761_ (.A1(_337_),
    .A2(_338_),
    .B1_N(_340_),
    .X(_341_));
 sky130_fd_sc_hd__a22o_1 _762_ (.A1(_269_),
    .A2(_334_),
    .B1(_341_),
    .B2(_054_),
    .X(_342_));
 sky130_fd_sc_hd__a21o_1 _763_ (.A1(_381_),
    .A2(_034_),
    .B1(_282_),
    .X(_343_));
 sky130_fd_sc_hd__a21o_1 _764_ (.A1(_334_),
    .A2(_343_),
    .B1(_283_),
    .X(_344_));
 sky130_fd_sc_hd__o211a_1 _765_ (.A1(_279_),
    .A2(_342_),
    .B1(_344_),
    .C1(_401_),
    .X(_345_));
 sky130_fd_sc_hd__a211o_1 _766_ (.A1(_386_),
    .A2(_335_),
    .B1(_345_),
    .C1(_383_),
    .X(_346_));
 sky130_fd_sc_hd__or2b_1 _767_ (.A(_387_),
    .B_N(_329_),
    .X(_347_));
 sky130_fd_sc_hd__a31o_1 _768_ (.A1(_051_),
    .A2(_328_),
    .A3(_347_),
    .B1(_331_),
    .X(_348_));
 sky130_fd_sc_hd__a32o_1 _769_ (.A1(_301_),
    .A2(_346_),
    .A3(_348_),
    .B1(_080_),
    .B2(net10),
    .X(_013_));
 sky130_fd_sc_hd__buf_2 _770_ (.A(\lcd.toggle ),
    .X(_349_));
 sky130_fd_sc_hd__nor2_1 _771_ (.A(_392_),
    .B(_329_),
    .Y(_350_));
 sky130_fd_sc_hd__and3_1 _772_ (.A(_041_),
    .B(_397_),
    .C(_350_),
    .X(_351_));
 sky130_fd_sc_hd__and3_1 _773_ (.A(_349_),
    .B(_385_),
    .C(_351_),
    .X(_352_));
 sky130_fd_sc_hd__a21oi_1 _774_ (.A1(\lcd.round[0] ),
    .A2(\lcd.round[1] ),
    .B1(_375_),
    .Y(_353_));
 sky130_fd_sc_hd__a211o_1 _775_ (.A1(_349_),
    .A2(_042_),
    .B1(_353_),
    .C1(_007_),
    .X(_354_));
 sky130_fd_sc_hd__and2b_1 _776_ (.A_N(_352_),
    .B(_354_),
    .X(_355_));
 sky130_fd_sc_hd__mux2_1 _777_ (.A0(_352_),
    .A1(_355_),
    .S(\lcd.round[0] ),
    .X(_356_));
 sky130_fd_sc_hd__clkbuf_1 _778_ (.A(_356_),
    .X(_014_));
 sky130_fd_sc_hd__a22o_1 _779_ (.A1(_035_),
    .A2(_352_),
    .B1(_355_),
    .B2(\lcd.round[1] ),
    .X(_015_));
 sky130_fd_sc_hd__nor2_1 _780_ (.A(_349_),
    .B(net4),
    .Y(_023_));
 sky130_fd_sc_hd__nor2_1 _781_ (.A(_375_),
    .B(_271_),
    .Y(_357_));
 sky130_fd_sc_hd__a22o_1 _782_ (.A1(_271_),
    .A2(_007_),
    .B1(_388_),
    .B2(_357_),
    .X(_024_));
 sky130_fd_sc_hd__nand2_1 _783_ (.A(_388_),
    .B(_347_),
    .Y(_358_));
 sky130_fd_sc_hd__a22o_1 _784_ (.A1(_284_),
    .A2(_007_),
    .B1(_358_),
    .B2(_349_),
    .X(_025_));
 sky130_fd_sc_hd__a41o_1 _785_ (.A1(_298_),
    .A2(_385_),
    .A3(_386_),
    .A4(_387_),
    .B1(_330_),
    .X(_359_));
 sky130_fd_sc_hd__a22o_1 _786_ (.A1(_052_),
    .A2(_007_),
    .B1(_359_),
    .B2(_349_),
    .X(_026_));
 sky130_fd_sc_hd__a31oi_1 _787_ (.A1(_052_),
    .A2(_284_),
    .A3(_271_),
    .B1(_376_),
    .Y(_360_));
 sky130_fd_sc_hd__o21ai_1 _788_ (.A1(_350_),
    .A2(_360_),
    .B1(_388_),
    .Y(_361_));
 sky130_fd_sc_hd__a22o_1 _789_ (.A1(_376_),
    .A2(_007_),
    .B1(_361_),
    .B2(_349_),
    .X(_027_));
 sky130_fd_sc_hd__nor2_1 _790_ (.A(_397_),
    .B(_350_),
    .Y(_362_));
 sky130_fd_sc_hd__a31o_1 _791_ (.A1(_284_),
    .A2(_271_),
    .A3(_398_),
    .B1(_362_),
    .X(_363_));
 sky130_fd_sc_hd__nand2_1 _792_ (.A(_388_),
    .B(_363_),
    .Y(_364_));
 sky130_fd_sc_hd__a22o_1 _793_ (.A1(_397_),
    .A2(_007_),
    .B1(_364_),
    .B2(_349_),
    .X(_028_));
 sky130_fd_sc_hd__a21oi_1 _794_ (.A1(_397_),
    .A2(_350_),
    .B1(_041_),
    .Y(_365_));
 sky130_fd_sc_hd__o21ai_1 _795_ (.A1(_351_),
    .A2(_365_),
    .B1(_388_),
    .Y(_366_));
 sky130_fd_sc_hd__a22o_1 _796_ (.A1(_041_),
    .A2(_007_),
    .B1(_366_),
    .B2(_349_),
    .X(_029_));
 sky130_fd_sc_hd__and3_1 _797_ (.A(_349_),
    .B(_381_),
    .C(_351_),
    .X(_367_));
 sky130_fd_sc_hd__a21oi_1 _798_ (.A1(_375_),
    .A2(net4),
    .B1(_367_),
    .Y(_368_));
 sky130_fd_sc_hd__a21o_1 _799_ (.A1(_349_),
    .A2(_351_),
    .B1(_381_),
    .X(_369_));
 sky130_fd_sc_hd__and2_1 _800_ (.A(_368_),
    .B(_369_),
    .X(_370_));
 sky130_fd_sc_hd__clkbuf_1 _801_ (.A(_370_),
    .X(_030_));
 sky130_fd_sc_hd__mux2_1 _802_ (.A0(_367_),
    .A1(_368_),
    .S(_033_),
    .X(_371_));
 sky130_fd_sc_hd__clkbuf_1 _803_ (.A(_371_),
    .X(_031_));
 sky130_fd_sc_hd__a21o_1 _804_ (.A1(_053_),
    .A2(_337_),
    .B1(_061_),
    .X(_372_));
 sky130_fd_sc_hd__o221ai_1 _805_ (.A1(_037_),
    .A2(_281_),
    .B1(_304_),
    .B2(_044_),
    .C1(_279_),
    .Y(_373_));
 sky130_fd_sc_hd__a32o_1 _806_ (.A1(_401_),
    .A2(_372_),
    .A3(_373_),
    .B1(_291_),
    .B2(_316_),
    .X(_374_));
 sky130_fd_sc_hd__a32o_1 _807_ (.A1(_042_),
    .A2(_301_),
    .A3(_374_),
    .B1(_080_),
    .B2(net5),
    .X(_032_));
 sky130_fd_sc_hd__dfxtp_1 _808_ (.CLK(clknet_2_1__leaf_clk),
    .D(_010_),
    .Q(net12));
 sky130_fd_sc_hd__dfxtp_1 _809_ (.CLK(clknet_2_2__leaf_clk),
    .D(_011_),
    .Q(net8));
 sky130_fd_sc_hd__dfxtp_1 _810_ (.CLK(clknet_2_2__leaf_clk),
    .D(_012_),
    .Q(net9));
 sky130_fd_sc_hd__dfxtp_1 _811_ (.CLK(clknet_2_2__leaf_clk),
    .D(_013_),
    .Q(net10));
 sky130_fd_sc_hd__dfxtp_1 _812_ (.CLK(clknet_2_3__leaf_clk),
    .D(_009_),
    .Q(\lcd.num_state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _813_ (.CLK(clknet_2_3__leaf_clk),
    .D(_008_),
    .Q(\lcd.num_state[1] ));
 sky130_fd_sc_hd__dfxtp_2 _814_ (.CLK(clknet_2_1__leaf_clk),
    .D(_014_),
    .Q(\lcd.round[0] ));
 sky130_fd_sc_hd__dfxtp_2 _815_ (.CLK(clknet_2_0__leaf_clk),
    .D(_015_),
    .Q(\lcd.round[1] ));
 sky130_fd_sc_hd__dfxtp_1 _816_ (.CLK(clknet_2_2__leaf_clk),
    .D(_016_),
    .Q(\lcd.rom_addr[0] ));
 sky130_fd_sc_hd__dfxtp_2 _817_ (.CLK(clknet_2_2__leaf_clk),
    .D(_017_),
    .Q(\lcd.rom_addr[1] ));
 sky130_fd_sc_hd__dfxtp_2 _818_ (.CLK(clknet_2_2__leaf_clk),
    .D(_018_),
    .Q(net11));
 sky130_fd_sc_hd__dfxtp_4 _819_ (.CLK(clknet_2_3__leaf_clk),
    .D(_019_),
    .Q(\lcd.rom_addr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _820_ (.CLK(clknet_2_3__leaf_clk),
    .D(_020_),
    .Q(\lcd.rom_addr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _821_ (.CLK(clknet_2_3__leaf_clk),
    .D(_021_),
    .Q(\lcd.rom_addr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _822_ (.CLK(clknet_2_2__leaf_clk),
    .D(_022_),
    .Q(\lcd.rom_addr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _823_ (.CLK(clknet_2_1__leaf_clk),
    .D(_023_),
    .Q(net6));
 sky130_fd_sc_hd__dfxtp_1 _824_ (.CLK(clknet_2_0__leaf_clk),
    .D(_007_),
    .Q(\lcd.toggle ));
 sky130_fd_sc_hd__dfxtp_1 _825_ (.CLK(clknet_2_3__leaf_clk),
    .D(_000_),
    .Q(\lcd.s_ROM[0] ));
 sky130_fd_sc_hd__dfxtp_1 _826_ (.CLK(clknet_2_3__leaf_clk),
    .D(_001_),
    .Q(\lcd.s_ROM[1] ));
 sky130_fd_sc_hd__dfxtp_1 _827_ (.CLK(clknet_2_3__leaf_clk),
    .D(_002_),
    .Q(\lcd.s_ROM[2] ));
 sky130_fd_sc_hd__dfxtp_1 _828_ (.CLK(clknet_2_0__leaf_clk),
    .D(_003_),
    .Q(\lcd.s_ROM[3] ));
 sky130_fd_sc_hd__dfxtp_1 _829_ (.CLK(clknet_2_3__leaf_clk),
    .D(_004_),
    .Q(\lcd.s_ROM[4] ));
 sky130_fd_sc_hd__dfxtp_1 _830_ (.CLK(clknet_2_2__leaf_clk),
    .D(_005_),
    .Q(\lcd.s_ROM[5] ));
 sky130_fd_sc_hd__dfxtp_1 _831_ (.CLK(clknet_2_2__leaf_clk),
    .D(_006_),
    .Q(\lcd.s_ROM[6] ));
 sky130_fd_sc_hd__dfxtp_1 _832_ (.CLK(clknet_2_1__leaf_clk),
    .D(_024_),
    .Q(\lcd.seq[0] ));
 sky130_fd_sc_hd__dfxtp_1 _833_ (.CLK(clknet_2_1__leaf_clk),
    .D(_025_),
    .Q(\lcd.seq[1] ));
 sky130_fd_sc_hd__dfxtp_2 _834_ (.CLK(clknet_2_0__leaf_clk),
    .D(_026_),
    .Q(\lcd.seq[2] ));
 sky130_fd_sc_hd__dfxtp_1 _835_ (.CLK(clknet_2_0__leaf_clk),
    .D(_027_),
    .Q(\lcd.seq[3] ));
 sky130_fd_sc_hd__dfxtp_2 _836_ (.CLK(clknet_2_0__leaf_clk),
    .D(_028_),
    .Q(\lcd.seq[4] ));
 sky130_fd_sc_hd__dfxtp_1 _837_ (.CLK(clknet_2_0__leaf_clk),
    .D(_029_),
    .Q(\lcd.seq[5] ));
 sky130_fd_sc_hd__dfxtp_2 _838_ (.CLK(clknet_2_1__leaf_clk),
    .D(_030_),
    .Q(\lcd.seq[6] ));
 sky130_fd_sc_hd__dfxtp_1 _839_ (.CLK(clknet_2_0__leaf_clk),
    .D(_031_),
    .Q(\lcd.seq[7] ));
 sky130_fd_sc_hd__dfxtp_1 _840_ (.CLK(clknet_2_1__leaf_clk),
    .D(_032_),
    .Q(net5));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_14 (.LO(net14));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_15 (.LO(net15));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_16 (.LO(net16));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_17 (.LO(net17));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_18 (.LO(net18));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_19 (.LO(net19));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_20 (.LO(net20));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_21 (.LO(net21));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_22 (.LO(net22));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_23 (.LO(net23));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_24 (.LO(net24));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_25 (.LO(net25));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_26 (.LO(net26));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_27 (.LO(net27));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_28 (.LO(net28));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_29 (.LO(net29));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_30 (.LO(net30));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_31 (.LO(net31));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_32 (.LO(net32));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_33 (.LO(net33));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_34 (.LO(net34));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_35 (.LO(net35));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_36 (.LO(net36));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_37 (.LO(net37));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_38 (.LO(net38));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_39 (.LO(net39));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_1 _868_ (.A(net12),
    .X(net7));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(io_in[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(io_in[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(io_in[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(rst),
    .X(net4));
 sky130_fd_sc_hd__buf_2 output5 (.A(net5),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_2 output6 (.A(net6),
    .X(io_out[1]));
 sky130_fd_sc_hd__buf_2 output7 (.A(net7),
    .X(io_out[2]));
 sky130_fd_sc_hd__buf_2 output8 (.A(net8),
    .X(io_out[3]));
 sky130_fd_sc_hd__buf_2 output9 (.A(net9),
    .X(io_out[4]));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_2 output11 (.A(net11),
    .X(io_out[6]));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .X(io_out[7]));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_13 (.LO(net13));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__827__D (.DIODE(_002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__816__D (.DIODE(_016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__674__A1 (.DIODE(_016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__637__A (.DIODE(_016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__622__A1 (.DIODE(_016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__618__A (.DIODE(_016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__607__B (.DIODE(_016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__546__B (.DIODE(_016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__818__D (.DIODE(_018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__609__B (.DIODE(_018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__605__A2 (.DIODE(_018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__601__A2 (.DIODE(_018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__600__B (.DIODE(_018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__594__A2 (.DIODE(_018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__578__A2 (.DIODE(_018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__558__B (.DIODE(_018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__557__A2 (.DIODE(_018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__519__A2 (.DIODE(_018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__819__D (.DIODE(_019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__653__A1 (.DIODE(_019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__646__A1 (.DIODE(_019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__641__A1 (.DIODE(_019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__627__A1 (.DIODE(_019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__626__B1 (.DIODE(_019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__621__A2 (.DIODE(_019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__597__A1 (.DIODE(_019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__585__A1 (.DIODE(_019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__509__A1 (.DIODE(_019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__821__D (.DIODE(_021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__678__A1 (.DIODE(_021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__648__C1 (.DIODE(_021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__644__A1 (.DIODE(_021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__643__A (.DIODE(_021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__629__A (.DIODE(_021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__625__A1 (.DIODE(_021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__616__A1 (.DIODE(_021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__604__A1 (.DIODE(_021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__539__A2 (.DIODE(_021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__822__D (.DIODE(_022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__679__S (.DIODE(_022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__664__A1 (.DIODE(_022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__651__B1 (.DIODE(_022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__633__B1 (.DIODE(_022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__616__C1 (.DIODE(_022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__591__C1 (.DIODE(_022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__580__C1 (.DIODE(_022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__568__A (.DIODE(_022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__565__S (.DIODE(_022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__760__A1 (.DIODE(_070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__753__A (.DIODE(_070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__748__B (.DIODE(_070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__736__S (.DIODE(_070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__721__S (.DIODE(_070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__688__A (.DIODE(_070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__687__S (.DIODE(_070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__495__A1 (.DIODE(_070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__481__A (.DIODE(_070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__473__A (.DIODE(_070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__675__A1 (.DIODE(_165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__670__A1 (.DIODE(_165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__659__A1 (.DIODE(_165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__642__D1 (.DIODE(_165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__627__C1 (.DIODE(_165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__624__A1 (.DIODE(_165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__611__A1 (.DIODE(_165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__602__C1 (.DIODE(_165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__597__C1 (.DIODE(_165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__573__B1 (.DIODE(_165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__798__A1 (.DIODE(_375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__781__A (.DIODE(_375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__774__B1 (.DIODE(_375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__718__A (.DIODE(_375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__496__B1 (.DIODE(_375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__470__B1 (.DIODE(_375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__466__B1 (.DIODE(_375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__464__B1 (.DIODE(_375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__419__A (.DIODE(_375_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(io_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(io_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(io_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__499__B1 (.DIODE(\lcd.rom_addr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__494__A (.DIODE(\lcd.rom_addr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__493__A (.DIODE(\lcd.rom_addr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__486__A (.DIODE(\lcd.rom_addr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__474__A (.DIODE(\lcd.rom_addr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__702__A1 (.DIODE(\lcd.seq[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__701__A (.DIODE(\lcd.seq[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__440__C (.DIODE(\lcd.seq[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__423__B_N (.DIODE(\lcd.seq[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__421__A (.DIODE(\lcd.seq[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__417__A (.DIODE(\lcd.seq[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__407__A2 (.DIODE(\lcd.seq[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__457__B1 (.DIODE(\lcd.seq[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__454__B1 (.DIODE(\lcd.seq[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__447__A_N (.DIODE(\lcd.seq[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__445__A (.DIODE(\lcd.seq[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__437__B (.DIODE(\lcd.seq[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__433__B (.DIODE(\lcd.seq[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__429__B (.DIODE(\lcd.seq[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__425__B (.DIODE(\lcd.seq[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__415__B (.DIODE(\lcd.seq[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__411__A (.DIODE(\lcd.seq[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(rst));
 sky130_fd_sc_hd__diode_2 ANTENNA_output5_A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__807__B2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_output8_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__734__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_output9_A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__752__B2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_output10_A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__769__B2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_output11_A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__530__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__522__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__487__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__475__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_output12_A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__868__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__719__B2 (.DIODE(net12));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_241 ();
 assign io_oeb[0] = net13;
 assign io_oeb[10] = net23;
 assign io_oeb[11] = net24;
 assign io_oeb[12] = net25;
 assign io_oeb[13] = net26;
 assign io_oeb[14] = net27;
 assign io_oeb[15] = net28;
 assign io_oeb[16] = net29;
 assign io_oeb[17] = net30;
 assign io_oeb[18] = net31;
 assign io_oeb[19] = net32;
 assign io_oeb[1] = net14;
 assign io_oeb[20] = net33;
 assign io_oeb[21] = net34;
 assign io_oeb[22] = net35;
 assign io_oeb[23] = net36;
 assign io_oeb[24] = net37;
 assign io_oeb[25] = net38;
 assign io_oeb[26] = net39;
 assign io_oeb[2] = net15;
 assign io_oeb[3] = net16;
 assign io_oeb[4] = net17;
 assign io_oeb[5] = net18;
 assign io_oeb[6] = net19;
 assign io_oeb[7] = net20;
 assign io_oeb[8] = net21;
 assign io_oeb[9] = net22;
endmodule

