magic
tech sky130B
magscale 1 2
timestamp 1680002332
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 842 2128 39178 37584
<< metal2 >>
rect 1766 39200 1822 40000
rect 5078 39200 5134 40000
rect 8390 39200 8446 40000
rect 11702 39200 11758 40000
rect 15014 39200 15070 40000
rect 18326 39200 18382 40000
rect 21638 39200 21694 40000
rect 24950 39200 25006 40000
rect 28262 39200 28318 40000
rect 31574 39200 31630 40000
rect 34886 39200 34942 40000
rect 38198 39200 38254 40000
rect 846 0 902 800
rect 2318 0 2374 800
rect 3790 0 3846 800
rect 5262 0 5318 800
rect 6734 0 6790 800
rect 8206 0 8262 800
rect 9678 0 9734 800
rect 11150 0 11206 800
rect 12622 0 12678 800
rect 14094 0 14150 800
rect 15566 0 15622 800
rect 17038 0 17094 800
rect 18510 0 18566 800
rect 19982 0 20038 800
rect 21454 0 21510 800
rect 22926 0 22982 800
rect 24398 0 24454 800
rect 25870 0 25926 800
rect 27342 0 27398 800
rect 28814 0 28870 800
rect 30286 0 30342 800
rect 31758 0 31814 800
rect 33230 0 33286 800
rect 34702 0 34758 800
rect 36174 0 36230 800
rect 37646 0 37702 800
rect 39118 0 39174 800
<< obsm2 >>
rect 848 39144 1710 39250
rect 1878 39144 5022 39250
rect 5190 39144 8334 39250
rect 8502 39144 11646 39250
rect 11814 39144 14958 39250
rect 15126 39144 18270 39250
rect 18438 39144 21582 39250
rect 21750 39144 24894 39250
rect 25062 39144 28206 39250
rect 28374 39144 31518 39250
rect 31686 39144 34830 39250
rect 34998 39144 38142 39250
rect 38310 39144 39172 39250
rect 848 856 39172 39144
rect 958 800 2262 856
rect 2430 800 3734 856
rect 3902 800 5206 856
rect 5374 800 6678 856
rect 6846 800 8150 856
rect 8318 800 9622 856
rect 9790 800 11094 856
rect 11262 800 12566 856
rect 12734 800 14038 856
rect 14206 800 15510 856
rect 15678 800 16982 856
rect 17150 800 18454 856
rect 18622 800 19926 856
rect 20094 800 21398 856
rect 21566 800 22870 856
rect 23038 800 24342 856
rect 24510 800 25814 856
rect 25982 800 27286 856
rect 27454 800 28758 856
rect 28926 800 30230 856
rect 30398 800 31702 856
rect 31870 800 33174 856
rect 33342 800 34646 856
rect 34814 800 36118 856
rect 36286 800 37590 856
rect 37758 800 39062 856
<< metal3 >>
rect 39200 19864 40000 19984
<< obsm3 >>
rect 4210 20064 39200 37569
rect 4210 19784 39120 20064
rect 4210 2143 39200 19784
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< obsm4 >>
rect 28211 22611 28277 31789
<< labels >>
rlabel metal2 s 1766 39200 1822 40000 6 clk
port 1 nsew signal input
rlabel metal2 s 8390 39200 8446 40000 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 11702 39200 11758 40000 6 io_in[1]
port 3 nsew signal input
rlabel metal2 s 15014 39200 15070 40000 6 io_in[2]
port 4 nsew signal input
rlabel metal2 s 18326 39200 18382 40000 6 io_in[3]
port 5 nsew signal input
rlabel metal2 s 21638 39200 21694 40000 6 io_in[4]
port 6 nsew signal input
rlabel metal2 s 24950 39200 25006 40000 6 io_in[5]
port 7 nsew signal input
rlabel metal2 s 28262 39200 28318 40000 6 io_in[6]
port 8 nsew signal input
rlabel metal2 s 31574 39200 31630 40000 6 io_in[7]
port 9 nsew signal input
rlabel metal2 s 34886 39200 34942 40000 6 io_in[8]
port 10 nsew signal input
rlabel metal2 s 38198 39200 38254 40000 6 io_in[9]
port 11 nsew signal input
rlabel metal3 s 39200 19864 40000 19984 6 io_oeb
port 12 nsew signal output
rlabel metal2 s 846 0 902 800 6 io_out[0]
port 13 nsew signal output
rlabel metal2 s 15566 0 15622 800 6 io_out[10]
port 14 nsew signal output
rlabel metal2 s 17038 0 17094 800 6 io_out[11]
port 15 nsew signal output
rlabel metal2 s 18510 0 18566 800 6 io_out[12]
port 16 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 io_out[13]
port 17 nsew signal output
rlabel metal2 s 21454 0 21510 800 6 io_out[14]
port 18 nsew signal output
rlabel metal2 s 22926 0 22982 800 6 io_out[15]
port 19 nsew signal output
rlabel metal2 s 24398 0 24454 800 6 io_out[16]
port 20 nsew signal output
rlabel metal2 s 25870 0 25926 800 6 io_out[17]
port 21 nsew signal output
rlabel metal2 s 27342 0 27398 800 6 io_out[18]
port 22 nsew signal output
rlabel metal2 s 28814 0 28870 800 6 io_out[19]
port 23 nsew signal output
rlabel metal2 s 2318 0 2374 800 6 io_out[1]
port 24 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 io_out[20]
port 25 nsew signal output
rlabel metal2 s 31758 0 31814 800 6 io_out[21]
port 26 nsew signal output
rlabel metal2 s 33230 0 33286 800 6 io_out[22]
port 27 nsew signal output
rlabel metal2 s 34702 0 34758 800 6 io_out[23]
port 28 nsew signal output
rlabel metal2 s 36174 0 36230 800 6 io_out[24]
port 29 nsew signal output
rlabel metal2 s 37646 0 37702 800 6 io_out[25]
port 30 nsew signal output
rlabel metal2 s 39118 0 39174 800 6 io_out[26]
port 31 nsew signal output
rlabel metal2 s 3790 0 3846 800 6 io_out[2]
port 32 nsew signal output
rlabel metal2 s 5262 0 5318 800 6 io_out[3]
port 33 nsew signal output
rlabel metal2 s 6734 0 6790 800 6 io_out[4]
port 34 nsew signal output
rlabel metal2 s 8206 0 8262 800 6 io_out[5]
port 35 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 io_out[6]
port 36 nsew signal output
rlabel metal2 s 11150 0 11206 800 6 io_out[7]
port 37 nsew signal output
rlabel metal2 s 12622 0 12678 800 6 io_out[8]
port 38 nsew signal output
rlabel metal2 s 14094 0 14150 800 6 io_out[9]
port 39 nsew signal output
rlabel metal2 s 5078 39200 5134 40000 6 rst
port 40 nsew signal input
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 41 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 41 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 42 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2868738
string GDS_FILE /run/media/tholin/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/AS5401/runs/23_03_28_13_15/results/signoff/tholin_avalonsemi_5401.magic.gds
string GDS_START 908300
<< end >>

