magic
tech sky130B
magscale 1 2
timestamp 1680008812
<< viali >>
rect 6653 29189 6687 29223
rect 10793 29189 10827 29223
rect 18153 29189 18187 29223
rect 30113 29189 30147 29223
rect 3157 29121 3191 29155
rect 3341 29121 3375 29155
rect 10241 29121 10275 29155
rect 14381 29121 14415 29155
rect 22017 29121 22051 29155
rect 25973 29121 26007 29155
rect 29101 29121 29135 29155
rect 29837 29121 29871 29155
rect 14657 29053 14691 29087
rect 28549 29053 28583 29087
rect 3341 28985 3375 29019
rect 6929 28985 6963 29019
rect 22201 28985 22235 29019
rect 26157 28985 26191 29019
rect 18245 28917 18279 28951
rect 3157 28645 3191 28679
rect 3341 28509 3375 28543
rect 3433 28509 3467 28543
rect 4997 28509 5031 28543
rect 7757 28509 7791 28543
rect 8217 28509 8251 28543
rect 9597 28509 9631 28543
rect 10333 28509 10367 28543
rect 11069 28509 11103 28543
rect 12541 28509 12575 28543
rect 14657 28509 14691 28543
rect 15301 28509 15335 28543
rect 18337 28509 18371 28543
rect 20821 28509 20855 28543
rect 21741 28509 21775 28543
rect 22753 28509 22787 28543
rect 22937 28509 22971 28543
rect 27077 28509 27111 28543
rect 28181 28509 28215 28543
rect 28365 28509 28399 28543
rect 3157 28441 3191 28475
rect 4169 28441 4203 28475
rect 11805 28441 11839 28475
rect 7665 28373 7699 28407
rect 8309 28373 8343 28407
rect 9505 28373 9539 28407
rect 10425 28373 10459 28407
rect 12633 28373 12667 28407
rect 14749 28373 14783 28407
rect 15393 28373 15427 28407
rect 18521 28373 18555 28407
rect 20913 28373 20947 28407
rect 21649 28373 21683 28407
rect 23765 28373 23799 28407
rect 27169 28373 27203 28407
rect 29193 28373 29227 28407
rect 13829 28169 13863 28203
rect 18153 28169 18187 28203
rect 24225 28169 24259 28203
rect 4782 28101 4816 28135
rect 8585 28101 8619 28135
rect 15945 28101 15979 28135
rect 27445 28101 27479 28135
rect 2964 28033 2998 28067
rect 8309 28033 8343 28067
rect 11161 28033 11195 28067
rect 12081 28033 12115 28067
rect 16221 28033 16255 28067
rect 17601 28033 17635 28067
rect 20821 28033 20855 28067
rect 21097 28033 21131 28067
rect 29469 28033 29503 28067
rect 2697 27965 2731 27999
rect 4537 27965 4571 27999
rect 7021 27965 7055 27999
rect 7757 27965 7791 27999
rect 12357 27965 12391 27999
rect 17509 27965 17543 27999
rect 19625 27965 19659 27999
rect 19901 27965 19935 27999
rect 21373 27965 21407 27999
rect 22477 27965 22511 27999
rect 22753 27965 22787 27999
rect 27169 27965 27203 27999
rect 10057 27897 10091 27931
rect 14473 27897 14507 27931
rect 4077 27829 4111 27863
rect 5917 27829 5951 27863
rect 11069 27829 11103 27863
rect 28917 27829 28951 27863
rect 29561 27829 29595 27863
rect 2329 27625 2363 27659
rect 2973 27625 3007 27659
rect 3341 27625 3375 27659
rect 6916 27625 6950 27659
rect 11148 27625 11182 27659
rect 19533 27625 19567 27659
rect 22121 27625 22155 27659
rect 22937 27625 22971 27659
rect 26617 27625 26651 27659
rect 5825 27557 5859 27591
rect 13645 27557 13679 27591
rect 23581 27557 23615 27591
rect 3433 27489 3467 27523
rect 3985 27489 4019 27523
rect 9229 27489 9263 27523
rect 9965 27489 9999 27523
rect 15485 27489 15519 27523
rect 18889 27489 18923 27523
rect 22385 27489 22419 27523
rect 25789 27489 25823 27523
rect 26065 27489 26099 27523
rect 28181 27489 28215 27523
rect 3157 27421 3191 27455
rect 6009 27421 6043 27455
rect 6101 27421 6135 27455
rect 6653 27421 6687 27455
rect 10885 27421 10919 27455
rect 13737 27421 13771 27455
rect 14565 27421 14599 27455
rect 18245 27421 18279 27455
rect 18521 27421 18555 27455
rect 19625 27421 19659 27455
rect 23029 27421 23063 27455
rect 23673 27421 23707 27455
rect 25697 27421 25731 27455
rect 26525 27421 26559 27455
rect 27629 27421 27663 27455
rect 27905 27421 27939 27455
rect 28733 27421 28767 27455
rect 2145 27353 2179 27387
rect 4230 27353 4264 27387
rect 5825 27353 5859 27387
rect 2345 27285 2379 27319
rect 2513 27285 2547 27319
rect 5365 27285 5399 27319
rect 8401 27285 8435 27319
rect 12633 27285 12667 27319
rect 20637 27285 20671 27319
rect 28825 27285 28859 27319
rect 7389 27081 7423 27115
rect 19441 27081 19475 27115
rect 3148 27013 3182 27047
rect 5181 27013 5215 27047
rect 13369 27013 13403 27047
rect 29929 27013 29963 27047
rect 2881 26945 2915 26979
rect 4813 26945 4847 26979
rect 4997 26945 5031 26979
rect 6837 26945 6871 26979
rect 7481 26945 7515 26979
rect 11897 26945 11931 26979
rect 14105 26945 14139 26979
rect 16057 26945 16091 26979
rect 18328 26945 18362 26979
rect 23673 26945 23707 26979
rect 24952 26945 24986 26979
rect 30205 26945 30239 26979
rect 4721 26877 4755 26911
rect 11805 26877 11839 26911
rect 16313 26877 16347 26911
rect 18061 26877 18095 26911
rect 23581 26877 23615 26911
rect 24685 26877 24719 26911
rect 4261 26809 4295 26843
rect 26065 26809 26099 26843
rect 6745 26741 6779 26775
rect 12265 26741 12299 26775
rect 14933 26741 14967 26775
rect 24041 26741 24075 26775
rect 28457 26741 28491 26775
rect 3433 26537 3467 26571
rect 12541 26537 12575 26571
rect 16313 26537 16347 26571
rect 24869 26537 24903 26571
rect 26065 26537 26099 26571
rect 26525 26537 26559 26571
rect 3341 26469 3375 26503
rect 8309 26469 8343 26503
rect 23213 26469 23247 26503
rect 4629 26401 4663 26435
rect 6469 26401 6503 26435
rect 8033 26401 8067 26435
rect 9413 26401 9447 26435
rect 9689 26401 9723 26435
rect 14565 26401 14599 26435
rect 15025 26401 15059 26435
rect 15669 26401 15703 26435
rect 15853 26401 15887 26435
rect 25329 26401 25363 26435
rect 25421 26401 25455 26435
rect 26157 26401 26191 26435
rect 3433 26333 3467 26367
rect 4261 26333 4295 26367
rect 4353 26333 4387 26367
rect 7941 26333 7975 26367
rect 9321 26333 9355 26367
rect 11161 26333 11195 26367
rect 14933 26333 14967 26367
rect 18797 26333 18831 26367
rect 20269 26333 20303 26367
rect 20453 26333 20487 26367
rect 21833 26333 21867 26367
rect 26341 26333 26375 26367
rect 28181 26333 28215 26367
rect 28365 26333 28399 26367
rect 29929 26333 29963 26367
rect 3157 26265 3191 26299
rect 4077 26265 4111 26299
rect 4445 26265 4479 26299
rect 7297 26265 7331 26299
rect 11428 26265 11462 26299
rect 15945 26265 15979 26299
rect 22100 26265 22134 26299
rect 25237 26265 25271 26299
rect 26065 26265 26099 26299
rect 18705 26197 18739 26231
rect 19441 26197 19475 26231
rect 29193 26197 29227 26231
rect 29837 26197 29871 26231
rect 2881 25993 2915 26027
rect 8309 25993 8343 26027
rect 10241 25993 10275 26027
rect 11713 25993 11747 26027
rect 12173 25993 12207 26027
rect 21005 25993 21039 26027
rect 22293 25993 22327 26027
rect 22753 25993 22787 26027
rect 29929 25993 29963 26027
rect 6837 25925 6871 25959
rect 12909 25925 12943 25959
rect 18705 25925 18739 25959
rect 4353 25857 4387 25891
rect 9128 25857 9162 25891
rect 12081 25857 12115 25891
rect 13185 25857 13219 25891
rect 18429 25857 18463 25891
rect 20913 25857 20947 25891
rect 22661 25857 22695 25891
rect 24860 25857 24894 25891
rect 6561 25789 6595 25823
rect 8861 25789 8895 25823
rect 12265 25789 12299 25823
rect 13001 25789 13035 25823
rect 20453 25789 20487 25823
rect 22845 25789 22879 25823
rect 24593 25789 24627 25823
rect 28181 25789 28215 25823
rect 28457 25789 28491 25823
rect 13093 25653 13127 25687
rect 13369 25653 13403 25687
rect 25973 25653 26007 25687
rect 4169 25449 4203 25483
rect 8125 25449 8159 25483
rect 9505 25449 9539 25483
rect 24777 25449 24811 25483
rect 27997 25449 28031 25483
rect 19993 25381 20027 25415
rect 10149 25313 10183 25347
rect 19533 25313 19567 25347
rect 25329 25313 25363 25347
rect 26065 25313 26099 25347
rect 26525 25313 26559 25347
rect 30113 25313 30147 25347
rect 2973 25245 3007 25279
rect 3157 25245 3191 25279
rect 3249 25245 3283 25279
rect 3985 25245 4019 25279
rect 4169 25245 4203 25279
rect 6745 25245 6779 25279
rect 9965 25245 9999 25279
rect 19625 25245 19659 25279
rect 22753 25245 22787 25279
rect 22937 25245 22971 25279
rect 25237 25245 25271 25279
rect 26157 25245 26191 25279
rect 27905 25245 27939 25279
rect 28733 25245 28767 25279
rect 29837 25245 29871 25279
rect 7012 25177 7046 25211
rect 10793 25177 10827 25211
rect 12541 25177 12575 25211
rect 2789 25109 2823 25143
rect 9873 25109 9907 25143
rect 22937 25109 22971 25143
rect 25145 25109 25179 25143
rect 28641 25109 28675 25143
rect 5917 24905 5951 24939
rect 6929 24905 6963 24939
rect 7389 24905 7423 24939
rect 8493 24905 8527 24939
rect 7297 24837 7331 24871
rect 28457 24837 28491 24871
rect 2809 24769 2843 24803
rect 3065 24769 3099 24803
rect 3525 24769 3559 24803
rect 6009 24769 6043 24803
rect 8585 24769 8619 24803
rect 11989 24769 12023 24803
rect 12633 24769 12667 24803
rect 14105 24769 14139 24803
rect 15945 24769 15979 24803
rect 17592 24769 17626 24803
rect 19993 24769 20027 24803
rect 22109 24769 22143 24803
rect 23305 24769 23339 24803
rect 25697 24769 25731 24803
rect 7573 24701 7607 24735
rect 8677 24701 8711 24735
rect 15025 24701 15059 24735
rect 15577 24701 15611 24735
rect 16037 24701 16071 24735
rect 17325 24701 17359 24735
rect 19901 24701 19935 24735
rect 22293 24701 22327 24735
rect 25789 24701 25823 24735
rect 26065 24701 26099 24735
rect 28181 24701 28215 24735
rect 29929 24701 29963 24735
rect 12541 24633 12575 24667
rect 18705 24633 18739 24667
rect 1685 24565 1719 24599
rect 4813 24565 4847 24599
rect 8125 24565 8159 24599
rect 11897 24565 11931 24599
rect 20361 24565 20395 24599
rect 24593 24565 24627 24599
rect 2973 24361 3007 24395
rect 4169 24361 4203 24395
rect 16037 24361 16071 24395
rect 17877 24361 17911 24395
rect 22753 24361 22787 24395
rect 4353 24293 4387 24327
rect 2421 24225 2455 24259
rect 3433 24225 3467 24259
rect 4813 24225 4847 24259
rect 7389 24225 7423 24259
rect 11345 24225 11379 24259
rect 11621 24225 11655 24259
rect 13369 24225 13403 24259
rect 18429 24225 18463 24259
rect 19901 24225 19935 24259
rect 19993 24225 20027 24259
rect 21373 24225 21407 24259
rect 25145 24225 25179 24259
rect 25973 24225 26007 24259
rect 29193 24225 29227 24259
rect 2329 24157 2363 24191
rect 2513 24157 2547 24191
rect 3157 24157 3191 24191
rect 3341 24157 3375 24191
rect 4997 24157 5031 24191
rect 5089 24157 5123 24191
rect 14289 24157 14323 24191
rect 18245 24157 18279 24191
rect 18337 24157 18371 24191
rect 23397 24157 23431 24191
rect 26065 24157 26099 24191
rect 26341 24157 26375 24191
rect 28181 24157 28215 24191
rect 28365 24157 28399 24191
rect 3985 24089 4019 24123
rect 6837 24089 6871 24123
rect 14565 24089 14599 24123
rect 21640 24089 21674 24123
rect 23213 24089 23247 24123
rect 4185 24021 4219 24055
rect 19441 24021 19475 24055
rect 19809 24021 19843 24055
rect 23581 24021 23615 24055
rect 24593 24021 24627 24055
rect 24961 24021 24995 24055
rect 25053 24021 25087 24055
rect 26157 24021 26191 24055
rect 3985 23817 4019 23851
rect 5273 23817 5307 23851
rect 13461 23817 13495 23851
rect 14105 23817 14139 23851
rect 16313 23817 16347 23851
rect 19901 23817 19935 23851
rect 22017 23817 22051 23851
rect 22477 23817 22511 23851
rect 26065 23817 26099 23851
rect 28365 23817 28399 23851
rect 2872 23749 2906 23783
rect 7849 23749 7883 23783
rect 9597 23749 9631 23783
rect 12541 23749 12575 23783
rect 18788 23749 18822 23783
rect 23397 23749 23431 23783
rect 25145 23749 25179 23783
rect 2605 23681 2639 23715
rect 4721 23681 4755 23715
rect 5181 23681 5215 23715
rect 5365 23681 5399 23715
rect 10149 23681 10183 23715
rect 10425 23681 10459 23715
rect 11805 23681 11839 23715
rect 13369 23681 13403 23715
rect 14013 23681 14047 23715
rect 15200 23681 15234 23715
rect 18521 23681 18555 23715
rect 21005 23681 21039 23715
rect 22385 23681 22419 23715
rect 26249 23681 26283 23715
rect 26525 23681 26559 23715
rect 28457 23681 28491 23715
rect 10241 23613 10275 23647
rect 14933 23613 14967 23647
rect 20913 23613 20947 23647
rect 22661 23613 22695 23647
rect 26433 23613 26467 23647
rect 4537 23477 4571 23511
rect 10149 23477 10183 23511
rect 10609 23477 10643 23511
rect 21373 23477 21407 23511
rect 26249 23477 26283 23511
rect 4261 23273 4295 23307
rect 4997 23273 5031 23307
rect 7573 23273 7607 23307
rect 9689 23273 9723 23307
rect 11897 23273 11931 23307
rect 15485 23273 15519 23307
rect 21097 23273 21131 23307
rect 23673 23273 23707 23307
rect 25973 23273 26007 23307
rect 26433 23273 26467 23307
rect 3065 23205 3099 23239
rect 12633 23205 12667 23239
rect 9229 23137 9263 23171
rect 13093 23137 13127 23171
rect 16129 23137 16163 23171
rect 19993 23137 20027 23171
rect 24593 23137 24627 23171
rect 26709 23137 26743 23171
rect 1685 23069 1719 23103
rect 1869 23069 1903 23103
rect 2881 23069 2915 23103
rect 3157 23069 3191 23103
rect 4353 23069 4387 23103
rect 5181 23069 5215 23103
rect 5825 23069 5859 23103
rect 9321 23069 9355 23103
rect 10425 23069 10459 23103
rect 13001 23069 13035 23103
rect 15945 23069 15979 23103
rect 19901 23069 19935 23103
rect 22569 23069 22603 23103
rect 23029 23069 23063 23103
rect 23122 23069 23156 23103
rect 23397 23069 23431 23103
rect 23535 23069 23569 23103
rect 24860 23069 24894 23103
rect 26801 23069 26835 23103
rect 28549 23069 28583 23103
rect 29193 23069 29227 23103
rect 1777 23001 1811 23035
rect 6101 23001 6135 23035
rect 23305 23001 23339 23035
rect 2697 22933 2731 22967
rect 15853 22933 15887 22967
rect 19441 22933 19475 22967
rect 19809 22933 19843 22967
rect 28457 22933 28491 22967
rect 29101 22933 29135 22967
rect 2053 22729 2087 22763
rect 6653 22729 6687 22763
rect 8769 22729 8803 22763
rect 15853 22729 15887 22763
rect 20269 22729 20303 22763
rect 21465 22729 21499 22763
rect 22385 22729 22419 22763
rect 23213 22729 23247 22763
rect 25881 22729 25915 22763
rect 30113 22729 30147 22763
rect 5457 22661 5491 22695
rect 7656 22661 7690 22695
rect 12909 22661 12943 22695
rect 14749 22661 14783 22695
rect 17785 22661 17819 22695
rect 19156 22661 19190 22695
rect 23581 22661 23615 22695
rect 28641 22661 28675 22695
rect 1961 22593 1995 22627
rect 2237 22593 2271 22627
rect 2964 22593 2998 22627
rect 4537 22593 4571 22627
rect 5641 22593 5675 22627
rect 6745 22593 6779 22627
rect 7389 22593 7423 22627
rect 9413 22593 9447 22627
rect 12081 22593 12115 22627
rect 12265 22593 12299 22627
rect 13185 22593 13219 22627
rect 15945 22593 15979 22627
rect 16957 22593 16991 22627
rect 18889 22593 18923 22627
rect 21281 22593 21315 22627
rect 21465 22593 21499 22627
rect 23397 22593 23431 22627
rect 24501 22593 24535 22627
rect 24768 22593 24802 22627
rect 28365 22593 28399 22627
rect 2697 22525 2731 22559
rect 4813 22525 4847 22559
rect 5825 22525 5859 22559
rect 9505 22525 9539 22559
rect 9781 22525 9815 22559
rect 15761 22525 15795 22559
rect 22477 22525 22511 22559
rect 22569 22525 22603 22559
rect 13093 22457 13127 22491
rect 2237 22389 2271 22423
rect 4077 22389 4111 22423
rect 12449 22389 12483 22423
rect 13185 22389 13219 22423
rect 15025 22389 15059 22423
rect 16313 22389 16347 22423
rect 22017 22389 22051 22423
rect 3433 22185 3467 22219
rect 5641 22185 5675 22219
rect 15577 22185 15611 22219
rect 24777 22185 24811 22219
rect 10149 22049 10183 22083
rect 10425 22049 10459 22083
rect 11437 22049 11471 22083
rect 11621 22049 11655 22083
rect 14749 22049 14783 22083
rect 16957 22049 16991 22083
rect 21465 22049 21499 22083
rect 25329 22049 25363 22083
rect 25973 22049 26007 22083
rect 26249 22049 26283 22083
rect 29193 22049 29227 22083
rect 2053 21981 2087 22015
rect 4997 21981 5031 22015
rect 5733 21981 5767 22015
rect 6285 21981 6319 22015
rect 10057 21981 10091 22015
rect 12173 21981 12207 22015
rect 12357 21981 12391 22015
rect 13001 21981 13035 22015
rect 16690 21981 16724 22015
rect 17877 21981 17911 22015
rect 21189 21981 21223 22015
rect 25237 21981 25271 22015
rect 26341 21981 26375 22015
rect 27445 21981 27479 22015
rect 28181 21981 28215 22015
rect 28457 21981 28491 22015
rect 29837 21981 29871 22015
rect 2320 21913 2354 21947
rect 4169 21913 4203 21947
rect 7021 21913 7055 21947
rect 13185 21913 13219 21947
rect 15025 21913 15059 21947
rect 17601 21913 17635 21947
rect 22937 21913 22971 21947
rect 23305 21913 23339 21947
rect 25145 21913 25179 21947
rect 30113 21913 30147 21947
rect 10977 21845 11011 21879
rect 11345 21845 11379 21879
rect 12265 21845 12299 21879
rect 12817 21845 12851 21879
rect 27537 21845 27571 21879
rect 10425 21641 10459 21675
rect 12817 21641 12851 21675
rect 16865 21641 16899 21675
rect 23397 21641 23431 21675
rect 25053 21641 25087 21675
rect 29377 21641 29411 21675
rect 4353 21573 4387 21607
rect 12449 21573 12483 21607
rect 12541 21573 12575 21607
rect 16068 21573 16102 21607
rect 18429 21573 18463 21607
rect 22262 21573 22296 21607
rect 25145 21573 25179 21607
rect 27905 21573 27939 21607
rect 5825 21505 5859 21539
rect 6745 21505 6779 21539
rect 9312 21505 9346 21539
rect 12173 21505 12207 21539
rect 12266 21505 12300 21539
rect 12638 21505 12672 21539
rect 16313 21505 16347 21539
rect 17233 21505 17267 21539
rect 18061 21505 18095 21539
rect 18337 21505 18371 21539
rect 22017 21505 22051 21539
rect 25881 21505 25915 21539
rect 2697 21437 2731 21471
rect 7021 21437 7055 21471
rect 9045 21437 9079 21471
rect 17325 21437 17359 21471
rect 17417 21437 17451 21471
rect 25237 21437 25271 21471
rect 26065 21437 26099 21471
rect 27629 21437 27663 21471
rect 5917 21301 5951 21335
rect 14933 21301 14967 21335
rect 24685 21301 24719 21335
rect 2973 21097 3007 21131
rect 3341 21097 3375 21131
rect 14565 21097 14599 21131
rect 16497 21097 16531 21131
rect 17785 21097 17819 21131
rect 25973 21097 26007 21131
rect 26893 21097 26927 21131
rect 7757 21029 7791 21063
rect 9413 21029 9447 21063
rect 12541 21029 12575 21063
rect 18705 21029 18739 21063
rect 20177 21029 20211 21063
rect 4353 20961 4387 20995
rect 5457 20961 5491 20995
rect 6009 20961 6043 20995
rect 6285 20961 6319 20995
rect 9873 20961 9907 20995
rect 9965 20961 9999 20995
rect 15008 20961 15042 20995
rect 18245 20961 18279 20995
rect 28181 20961 28215 20995
rect 29009 20961 29043 20995
rect 3157 20893 3191 20927
rect 3433 20893 3467 20927
rect 3985 20893 4019 20927
rect 4169 20893 4203 20927
rect 5549 20893 5583 20927
rect 10609 20893 10643 20927
rect 10876 20893 10910 20927
rect 12455 20893 12489 20927
rect 12633 20893 12667 20927
rect 14749 20893 14783 20927
rect 15301 20893 15335 20927
rect 15853 20893 15887 20927
rect 16589 20893 16623 20927
rect 17509 20893 17543 20927
rect 17601 20893 17635 20927
rect 18429 20893 18463 20927
rect 18797 20893 18831 20927
rect 19533 20893 19567 20927
rect 19993 20893 20027 20927
rect 20913 20893 20947 20927
rect 24593 20893 24627 20927
rect 24849 20893 24883 20927
rect 26801 20893 26835 20927
rect 28457 20893 28491 20927
rect 9781 20825 9815 20859
rect 21180 20825 21214 20859
rect 11989 20757 12023 20791
rect 15117 20757 15151 20791
rect 15209 20757 15243 20791
rect 22293 20757 22327 20791
rect 8309 20553 8343 20587
rect 10425 20553 10459 20587
rect 15485 20553 15519 20587
rect 18613 20553 18647 20587
rect 19901 20553 19935 20587
rect 5917 20485 5951 20519
rect 6837 20485 6871 20519
rect 18429 20485 18463 20519
rect 4721 20417 4755 20451
rect 5825 20417 5859 20451
rect 9312 20417 9346 20451
rect 14289 20417 14323 20451
rect 14473 20417 14507 20451
rect 14657 20417 14691 20451
rect 15577 20417 15611 20451
rect 16865 20417 16899 20451
rect 17141 20417 17175 20451
rect 17233 20417 17267 20451
rect 19717 20417 19751 20451
rect 20821 20417 20855 20451
rect 21097 20417 21131 20451
rect 22201 20417 22235 20451
rect 24501 20417 24535 20451
rect 24685 20417 24719 20451
rect 2513 20349 2547 20383
rect 2789 20349 2823 20383
rect 4261 20349 4295 20383
rect 6561 20349 6595 20383
rect 9045 20349 9079 20383
rect 19533 20349 19567 20383
rect 21373 20349 21407 20383
rect 4813 20281 4847 20315
rect 18061 20281 18095 20315
rect 18429 20213 18463 20247
rect 22109 20213 22143 20247
rect 24593 20213 24627 20247
rect 3157 20009 3191 20043
rect 4077 20009 4111 20043
rect 9505 20009 9539 20043
rect 18889 20009 18923 20043
rect 22201 19941 22235 19975
rect 7113 19873 7147 19907
rect 10057 19873 10091 19907
rect 17509 19873 17543 19907
rect 19901 19873 19935 19907
rect 20729 19873 20763 19907
rect 25329 19873 25363 19907
rect 27261 19873 27295 19907
rect 2605 19805 2639 19839
rect 3249 19805 3283 19839
rect 4169 19805 4203 19839
rect 5273 19805 5307 19839
rect 6101 19805 6135 19839
rect 9873 19805 9907 19839
rect 9965 19805 9999 19839
rect 19533 19805 19567 19839
rect 19717 19805 19751 19839
rect 20453 19805 20487 19839
rect 17776 19737 17810 19771
rect 25053 19737 25087 19771
rect 27528 19737 27562 19771
rect 2513 19669 2547 19703
rect 5457 19669 5491 19703
rect 24685 19669 24719 19703
rect 25145 19669 25179 19703
rect 28641 19669 28675 19703
rect 18429 19465 18463 19499
rect 23673 19465 23707 19499
rect 25881 19465 25915 19499
rect 27813 19465 27847 19499
rect 27905 19465 27939 19499
rect 2145 19397 2179 19431
rect 3893 19397 3927 19431
rect 24409 19397 24443 19431
rect 27997 19397 28031 19431
rect 12909 19329 12943 19363
rect 13165 19329 13199 19363
rect 15117 19329 15151 19363
rect 15761 19329 15795 19363
rect 18521 19329 18555 19363
rect 23489 19329 23523 19363
rect 23673 19329 23707 19363
rect 24133 19329 24167 19363
rect 28917 19329 28951 19363
rect 29009 19329 29043 19363
rect 29193 19329 29227 19363
rect 1869 19261 1903 19295
rect 14841 19261 14875 19295
rect 15393 19261 15427 19295
rect 16129 19261 16163 19295
rect 29377 19261 29411 19295
rect 27629 19193 27663 19227
rect 14289 19125 14323 19159
rect 28181 19125 28215 19159
rect 2421 18921 2455 18955
rect 3341 18921 3375 18955
rect 13001 18921 13035 18955
rect 20085 18921 20119 18955
rect 28457 18921 28491 18955
rect 29193 18921 29227 18955
rect 13553 18785 13587 18819
rect 21281 18785 21315 18819
rect 24593 18785 24627 18819
rect 27721 18785 27755 18819
rect 29745 18785 29779 18819
rect 30021 18785 30055 18819
rect 2513 18717 2547 18751
rect 3433 18717 3467 18751
rect 7757 18717 7791 18751
rect 8217 18717 8251 18751
rect 9137 18717 9171 18751
rect 13369 18717 13403 18751
rect 15117 18717 15151 18751
rect 17877 18717 17911 18751
rect 17969 18717 18003 18751
rect 19441 18717 19475 18751
rect 19901 18717 19935 18751
rect 21097 18717 21131 18751
rect 27445 18717 27479 18751
rect 27629 18717 27663 18751
rect 27849 18717 27883 18751
rect 28549 18717 28583 18751
rect 29009 18717 29043 18751
rect 29193 18717 29227 18751
rect 30113 18717 30147 18751
rect 13461 18649 13495 18683
rect 17417 18649 17451 18683
rect 17509 18649 17543 18683
rect 18061 18649 18095 18683
rect 24869 18649 24903 18683
rect 27721 18649 27755 18683
rect 7665 18581 7699 18615
rect 8309 18581 8343 18615
rect 9229 18581 9263 18615
rect 16405 18581 16439 18615
rect 20637 18581 20671 18615
rect 21005 18581 21039 18615
rect 26341 18581 26375 18615
rect 12357 18377 12391 18411
rect 14565 18377 14599 18411
rect 17141 18377 17175 18411
rect 17233 18377 17267 18411
rect 22385 18377 22419 18411
rect 24869 18377 24903 18411
rect 25329 18377 25363 18411
rect 4077 18309 4111 18343
rect 7481 18309 7515 18343
rect 9229 18309 9263 18343
rect 15393 18309 15427 18343
rect 17325 18309 17359 18343
rect 17693 18309 17727 18343
rect 19984 18309 20018 18343
rect 5273 18241 5307 18275
rect 5917 18241 5951 18275
rect 6561 18241 6595 18275
rect 9873 18241 9907 18275
rect 13185 18241 13219 18275
rect 13452 18241 13486 18275
rect 15485 18241 15519 18275
rect 15577 18241 15611 18275
rect 16037 18241 16071 18275
rect 18981 18241 19015 18275
rect 19073 18241 19107 18275
rect 19257 18241 19291 18275
rect 25237 18241 25271 18275
rect 29837 18241 29871 18275
rect 2053 18173 2087 18207
rect 2329 18173 2363 18207
rect 6653 18173 6687 18207
rect 7205 18173 7239 18207
rect 12449 18173 12483 18207
rect 12541 18173 12575 18207
rect 15945 18173 15979 18207
rect 16957 18173 16991 18207
rect 19717 18173 19751 18207
rect 22477 18173 22511 18207
rect 22661 18173 22695 18207
rect 25421 18173 25455 18207
rect 30113 18173 30147 18207
rect 5181 18105 5215 18139
rect 5825 18037 5859 18071
rect 9781 18037 9815 18071
rect 11989 18037 12023 18071
rect 21097 18037 21131 18071
rect 22017 18037 22051 18071
rect 2053 17833 2087 17867
rect 2697 17833 2731 17867
rect 13185 17833 13219 17867
rect 14289 17833 14323 17867
rect 21465 17833 21499 17867
rect 10885 17765 10919 17799
rect 8401 17697 8435 17731
rect 9137 17697 9171 17731
rect 9413 17697 9447 17731
rect 12081 17697 12115 17731
rect 14749 17697 14783 17731
rect 14841 17697 14875 17731
rect 20085 17697 20119 17731
rect 2145 17629 2179 17663
rect 2605 17629 2639 17663
rect 3433 17629 3467 17663
rect 5089 17629 5123 17663
rect 5733 17629 5767 17663
rect 5825 17629 5859 17663
rect 11805 17629 11839 17663
rect 15669 17629 15703 17663
rect 17969 17629 18003 17663
rect 18429 17629 18463 17663
rect 18521 17629 18555 17663
rect 20352 17629 20386 17663
rect 22201 17629 22235 17663
rect 26617 17629 26651 17663
rect 6377 17561 6411 17595
rect 8125 17561 8159 17595
rect 14657 17561 14691 17595
rect 17417 17561 17451 17595
rect 18061 17561 18095 17595
rect 18613 17561 18647 17595
rect 22468 17561 22502 17595
rect 3341 17493 3375 17527
rect 23581 17493 23615 17527
rect 26525 17493 26559 17527
rect 6837 17289 6871 17323
rect 7481 17289 7515 17323
rect 22385 17289 22419 17323
rect 3985 17221 4019 17255
rect 13645 17221 13679 17255
rect 14013 17221 14047 17255
rect 14197 17221 14231 17255
rect 27445 17221 27479 17255
rect 2881 17153 2915 17187
rect 3341 17153 3375 17187
rect 6009 17153 6043 17187
rect 6745 17153 6779 17187
rect 7389 17153 7423 17187
rect 11713 17153 11747 17187
rect 11969 17153 12003 17187
rect 14105 17153 14139 17187
rect 15209 17153 15243 17187
rect 15485 17153 15519 17187
rect 15945 17153 15979 17187
rect 16865 17153 16899 17187
rect 17509 17153 17543 17187
rect 18245 17153 18279 17187
rect 18337 17153 18371 17187
rect 18429 17153 18463 17187
rect 18613 17153 18647 17187
rect 19073 17153 19107 17187
rect 19349 17153 19383 17187
rect 20913 17153 20947 17187
rect 22753 17153 22787 17187
rect 22845 17153 22879 17187
rect 23857 17153 23891 17187
rect 26065 17153 26099 17187
rect 5733 17085 5767 17119
rect 14381 17085 14415 17119
rect 15761 17085 15795 17119
rect 17233 17085 17267 17119
rect 19441 17085 19475 17119
rect 21005 17085 21039 17119
rect 22937 17085 22971 17119
rect 23765 17085 23799 17119
rect 27997 17085 28031 17119
rect 29009 17085 29043 17119
rect 29745 17085 29779 17119
rect 13093 17017 13127 17051
rect 15577 17017 15611 17051
rect 2789 16949 2823 16983
rect 3433 16949 3467 16983
rect 18061 16949 18095 16983
rect 21281 16949 21315 16983
rect 24225 16949 24259 16983
rect 26157 16949 26191 16983
rect 11805 16745 11839 16779
rect 14381 16745 14415 16779
rect 27905 16745 27939 16779
rect 17049 16677 17083 16711
rect 9781 16609 9815 16643
rect 12265 16609 12299 16643
rect 12357 16609 12391 16643
rect 13369 16609 13403 16643
rect 14473 16609 14507 16643
rect 16313 16609 16347 16643
rect 19993 16609 20027 16643
rect 26157 16609 26191 16643
rect 26433 16609 26467 16643
rect 2697 16541 2731 16575
rect 2789 16541 2823 16575
rect 4537 16541 4571 16575
rect 4629 16541 4663 16575
rect 6193 16541 6227 16575
rect 13553 16541 13587 16575
rect 13737 16541 13771 16575
rect 14749 16541 14783 16575
rect 15853 16541 15887 16575
rect 16865 16541 16899 16575
rect 17141 16541 17175 16575
rect 17601 16541 17635 16575
rect 17877 16541 17911 16575
rect 18021 16541 18055 16575
rect 28549 16541 28583 16575
rect 29745 16541 29779 16575
rect 6469 16473 6503 16507
rect 9597 16473 9631 16507
rect 15577 16473 15611 16507
rect 15945 16473 15979 16507
rect 17785 16473 17819 16507
rect 18170 16473 18204 16507
rect 9137 16405 9171 16439
rect 9505 16405 9539 16439
rect 12173 16405 12207 16439
rect 15761 16405 15795 16439
rect 19441 16405 19475 16439
rect 19809 16405 19843 16439
rect 19901 16405 19935 16439
rect 28641 16405 28675 16439
rect 29837 16405 29871 16439
rect 7481 16201 7515 16235
rect 10977 16201 11011 16235
rect 28273 16201 28307 16235
rect 2973 16133 3007 16167
rect 4721 16133 4755 16167
rect 9422 16133 9456 16167
rect 14749 16133 14783 16167
rect 18696 16133 18730 16167
rect 10149 16065 10183 16099
rect 10885 16065 10919 16099
rect 12173 16065 12207 16099
rect 13001 16065 13035 16099
rect 15393 16065 15427 16099
rect 15577 16065 15611 16099
rect 16221 16065 16255 16099
rect 23765 16065 23799 16099
rect 24593 16065 24627 16099
rect 30021 16065 30055 16099
rect 2697 15997 2731 16031
rect 7573 15997 7607 16031
rect 7757 15997 7791 16031
rect 9689 15997 9723 16031
rect 15209 15997 15243 16031
rect 18429 15997 18463 16031
rect 23581 15997 23615 16031
rect 24317 15997 24351 16031
rect 24501 15997 24535 16031
rect 29745 15997 29779 16031
rect 10333 15929 10367 15963
rect 16129 15929 16163 15963
rect 7113 15861 7147 15895
rect 8309 15861 8343 15895
rect 12081 15861 12115 15895
rect 19809 15861 19843 15895
rect 24961 15861 24995 15895
rect 6193 15657 6227 15691
rect 25973 15657 26007 15691
rect 7573 15521 7607 15555
rect 13277 15521 13311 15555
rect 23857 15521 23891 15555
rect 5273 15453 5307 15487
rect 7306 15453 7340 15487
rect 9321 15453 9355 15487
rect 12541 15453 12575 15487
rect 13737 15453 13771 15487
rect 16589 15453 16623 15487
rect 19441 15453 19475 15487
rect 19625 15453 19659 15487
rect 21465 15453 21499 15487
rect 21925 15453 21959 15487
rect 22109 15453 22143 15487
rect 23673 15453 23707 15487
rect 24593 15453 24627 15487
rect 24860 15453 24894 15487
rect 27445 15453 27479 15487
rect 28181 15453 28215 15487
rect 9588 15385 9622 15419
rect 12265 15385 12299 15419
rect 13645 15385 13679 15419
rect 16856 15385 16890 15419
rect 21281 15385 21315 15419
rect 29193 15385 29227 15419
rect 5181 15317 5215 15351
rect 10701 15317 10735 15351
rect 13553 15317 13587 15351
rect 17969 15317 18003 15351
rect 19625 15317 19659 15351
rect 21097 15317 21131 15351
rect 21925 15317 21959 15351
rect 23305 15317 23339 15351
rect 23765 15317 23799 15351
rect 27537 15317 27571 15351
rect 8033 15113 8067 15147
rect 9781 15113 9815 15147
rect 10241 15113 10275 15147
rect 11069 15113 11103 15147
rect 16865 15113 16899 15147
rect 22109 15113 22143 15147
rect 24593 15113 24627 15147
rect 29653 15113 29687 15147
rect 15025 15045 15059 15079
rect 17325 15045 17359 15079
rect 18613 15045 18647 15079
rect 18981 15045 19015 15079
rect 20729 15045 20763 15079
rect 20821 15045 20855 15079
rect 23480 15045 23514 15079
rect 28181 15045 28215 15079
rect 5273 14977 5307 15011
rect 6561 14977 6595 15011
rect 10149 14977 10183 15011
rect 11161 14977 11195 15011
rect 11897 14977 11931 15011
rect 17233 14977 17267 15011
rect 18797 14977 18831 15011
rect 19625 14977 19659 15011
rect 20453 14977 20487 15011
rect 20546 14977 20580 15011
rect 20959 14977 20993 15011
rect 22017 14977 22051 15011
rect 22293 14977 22327 15011
rect 23213 14977 23247 15011
rect 25329 14977 25363 15011
rect 5365 14909 5399 14943
rect 5917 14909 5951 14943
rect 10333 14909 10367 14943
rect 12173 14909 12207 14943
rect 13921 14909 13955 14943
rect 17417 14909 17451 14943
rect 19717 14909 19751 14943
rect 19993 14909 20027 14943
rect 22477 14909 22511 14943
rect 25421 14909 25455 14943
rect 27905 14909 27939 14943
rect 21097 14841 21131 14875
rect 15301 14773 15335 14807
rect 25697 14773 25731 14807
rect 21465 14569 21499 14603
rect 21925 14569 21959 14603
rect 27997 14569 28031 14603
rect 13093 14501 13127 14535
rect 14381 14501 14415 14535
rect 4537 14433 4571 14467
rect 5089 14433 5123 14467
rect 5365 14433 5399 14467
rect 7665 14433 7699 14467
rect 9505 14433 9539 14467
rect 9781 14433 9815 14467
rect 10885 14433 10919 14467
rect 11713 14433 11747 14467
rect 11989 14433 12023 14467
rect 14933 14433 14967 14467
rect 19625 14433 19659 14467
rect 24685 14433 24719 14467
rect 25145 14433 25179 14467
rect 4629 14365 4663 14399
rect 7573 14365 7607 14399
rect 9413 14365 9447 14399
rect 10977 14365 11011 14399
rect 11805 14365 11839 14399
rect 11897 14365 11931 14399
rect 12173 14365 12207 14399
rect 13277 14365 13311 14399
rect 14473 14365 14507 14399
rect 21649 14365 21683 14399
rect 21741 14365 21775 14399
rect 24777 14365 24811 14399
rect 27445 14365 27479 14399
rect 28089 14365 28123 14399
rect 28733 14365 28767 14399
rect 30297 14365 30331 14399
rect 7113 14297 7147 14331
rect 15200 14297 15234 14331
rect 19892 14297 19926 14331
rect 21465 14297 21499 14331
rect 30021 14297 30055 14331
rect 11529 14229 11563 14263
rect 16313 14229 16347 14263
rect 21005 14229 21039 14263
rect 27353 14229 27387 14263
rect 28641 14229 28675 14263
rect 5917 14025 5951 14059
rect 14197 14025 14231 14059
rect 15577 14025 15611 14059
rect 16037 14025 16071 14059
rect 16865 14025 16899 14059
rect 17233 14025 17267 14059
rect 19993 14025 20027 14059
rect 20453 14025 20487 14059
rect 26065 14025 26099 14059
rect 30113 14025 30147 14059
rect 4445 13957 4479 13991
rect 23397 13957 23431 13991
rect 25605 13957 25639 13991
rect 6745 13889 6779 13923
rect 12265 13889 12299 13923
rect 12532 13889 12566 13923
rect 14105 13889 14139 13923
rect 15945 13889 15979 13923
rect 20361 13889 20395 13923
rect 22569 13889 22603 13923
rect 25881 13889 25915 13923
rect 27169 13889 27203 13923
rect 28365 13889 28399 13923
rect 4169 13821 4203 13855
rect 6653 13821 6687 13855
rect 7113 13821 7147 13855
rect 16221 13821 16255 13855
rect 17325 13821 17359 13855
rect 17417 13821 17451 13855
rect 20545 13821 20579 13855
rect 22477 13821 22511 13855
rect 22937 13821 22971 13855
rect 25697 13821 25731 13855
rect 28641 13821 28675 13855
rect 13645 13685 13679 13719
rect 24685 13685 24719 13719
rect 25605 13685 25639 13719
rect 27261 13685 27295 13719
rect 4813 13481 4847 13515
rect 12725 13481 12759 13515
rect 18613 13481 18647 13515
rect 21097 13481 21131 13515
rect 29837 13481 29871 13515
rect 28733 13413 28767 13447
rect 5733 13345 5767 13379
rect 9137 13345 9171 13379
rect 13185 13345 13219 13379
rect 13369 13345 13403 13379
rect 18153 13345 18187 13379
rect 20821 13345 20855 13379
rect 26985 13345 27019 13379
rect 4905 13277 4939 13311
rect 6837 13277 6871 13311
rect 16221 13277 16255 13311
rect 18245 13277 18279 13311
rect 20729 13277 20763 13311
rect 24041 13277 24075 13311
rect 29929 13277 29963 13311
rect 9382 13209 9416 13243
rect 16488 13209 16522 13243
rect 24593 13209 24627 13243
rect 27261 13209 27295 13243
rect 10517 13141 10551 13175
rect 13093 13141 13127 13175
rect 17601 13141 17635 13175
rect 23949 13141 23983 13175
rect 26065 13141 26099 13175
rect 5825 12937 5859 12971
rect 9229 12937 9263 12971
rect 9689 12937 9723 12971
rect 14749 12937 14783 12971
rect 16865 12937 16899 12971
rect 7481 12869 7515 12903
rect 13176 12869 13210 12903
rect 25053 12869 25087 12903
rect 28181 12869 28215 12903
rect 29745 12869 29779 12903
rect 5181 12801 5215 12835
rect 5365 12801 5399 12835
rect 7297 12801 7331 12835
rect 8401 12801 8435 12835
rect 9597 12801 9631 12835
rect 15117 12801 15151 12835
rect 17233 12801 17267 12835
rect 17325 12801 17359 12835
rect 19625 12801 19659 12835
rect 22937 12801 22971 12835
rect 23397 12801 23431 12835
rect 24133 12801 24167 12835
rect 27445 12801 27479 12835
rect 8309 12733 8343 12767
rect 9873 12733 9907 12767
rect 12909 12733 12943 12767
rect 15209 12733 15243 12767
rect 15301 12733 15335 12767
rect 17417 12733 17451 12767
rect 19533 12733 19567 12767
rect 19993 12733 20027 12767
rect 24225 12733 24259 12767
rect 24777 12733 24811 12767
rect 26525 12733 26559 12767
rect 29193 12733 29227 12767
rect 14289 12665 14323 12699
rect 7665 12597 7699 12631
rect 8769 12597 8803 12631
rect 22845 12597 22879 12631
rect 23489 12597 23523 12631
rect 17233 12393 17267 12427
rect 23949 12393 23983 12427
rect 7021 12257 7055 12291
rect 22201 12257 22235 12291
rect 22477 12257 22511 12291
rect 25329 12257 25363 12291
rect 26157 12257 26191 12291
rect 4997 12189 5031 12223
rect 5641 12189 5675 12223
rect 6929 12189 6963 12223
rect 7113 12189 7147 12223
rect 7573 12189 7607 12223
rect 7666 12189 7700 12223
rect 7849 12189 7883 12223
rect 8079 12189 8113 12223
rect 12357 12189 12391 12223
rect 12541 12189 12575 12223
rect 15853 12189 15887 12223
rect 16120 12189 16154 12223
rect 17877 12189 17911 12223
rect 5549 12121 5583 12155
rect 7941 12121 7975 12155
rect 4905 12053 4939 12087
rect 8217 12053 8251 12087
rect 12449 12053 12483 12087
rect 17785 12053 17819 12087
rect 8677 11849 8711 11883
rect 13001 11849 13035 11883
rect 4445 11781 4479 11815
rect 23673 11781 23707 11815
rect 4169 11713 4203 11747
rect 7104 11713 7138 11747
rect 8677 11713 8711 11747
rect 8861 11713 8895 11747
rect 9597 11713 9631 11747
rect 10425 11713 10459 11747
rect 10701 11713 10735 11747
rect 18521 11713 18555 11747
rect 18981 11713 19015 11747
rect 19901 11713 19935 11747
rect 20729 11713 20763 11747
rect 22201 11713 22235 11747
rect 22937 11713 22971 11747
rect 5917 11645 5951 11679
rect 6837 11645 6871 11679
rect 9505 11645 9539 11679
rect 9965 11645 9999 11679
rect 10517 11645 10551 11679
rect 13093 11645 13127 11679
rect 13277 11645 13311 11679
rect 17877 11645 17911 11679
rect 8217 11577 8251 11611
rect 10425 11509 10459 11543
rect 10885 11509 10919 11543
rect 12633 11509 12667 11543
rect 19073 11509 19107 11543
rect 19809 11509 19843 11543
rect 20821 11509 20855 11543
rect 22109 11509 22143 11543
rect 7573 11305 7607 11339
rect 13461 11305 13495 11339
rect 18429 11305 18463 11339
rect 21189 11305 21223 11339
rect 23489 11305 23523 11339
rect 29009 11237 29043 11271
rect 30297 11237 30331 11271
rect 5273 11169 5307 11203
rect 5733 11169 5767 11203
rect 8033 11169 8067 11203
rect 8217 11169 8251 11203
rect 12081 11169 12115 11203
rect 16129 11169 16163 11203
rect 16681 11169 16715 11203
rect 16957 11169 16991 11203
rect 19441 11169 19475 11203
rect 19717 11169 19751 11203
rect 21741 11169 21775 11203
rect 22017 11169 22051 11203
rect 25881 11169 25915 11203
rect 29193 11169 29227 11203
rect 29837 11169 29871 11203
rect 4261 11101 4295 11135
rect 5089 11101 5123 11135
rect 9873 11101 9907 11135
rect 12348 11101 12382 11135
rect 16221 11101 16255 11135
rect 24685 11101 24719 11135
rect 24869 11101 24903 11135
rect 25697 11101 25731 11135
rect 29929 11101 29963 11135
rect 4169 11033 4203 11067
rect 7941 11033 7975 11067
rect 25789 11033 25823 11067
rect 28733 11033 28767 11067
rect 9965 10965 9999 10999
rect 24869 10965 24903 10999
rect 25329 10965 25363 10999
rect 4261 10761 4295 10795
rect 7573 10761 7607 10795
rect 12633 10761 12667 10795
rect 18613 10761 18647 10795
rect 28089 10761 28123 10795
rect 29745 10761 29779 10795
rect 5733 10693 5767 10727
rect 7757 10693 7791 10727
rect 7941 10693 7975 10727
rect 10517 10693 10551 10727
rect 12173 10693 12207 10727
rect 16221 10693 16255 10727
rect 17141 10693 17175 10727
rect 20361 10693 20395 10727
rect 23121 10693 23155 10727
rect 25053 10693 25087 10727
rect 27721 10693 27755 10727
rect 27813 10693 27847 10727
rect 29101 10693 29135 10727
rect 6745 10625 6779 10659
rect 11161 10625 11195 10659
rect 12449 10625 12483 10659
rect 13452 10625 13486 10659
rect 16313 10625 16347 10659
rect 16865 10625 16899 10659
rect 24777 10625 24811 10659
rect 27537 10625 27571 10659
rect 27905 10625 27939 10659
rect 28641 10625 28675 10659
rect 28733 10625 28767 10659
rect 28825 10625 28859 10659
rect 28917 10625 28951 10659
rect 29653 10625 29687 10659
rect 29837 10625 29871 10659
rect 6009 10557 6043 10591
rect 6653 10557 6687 10591
rect 12357 10557 12391 10591
rect 13185 10557 13219 10591
rect 19533 10557 19567 10591
rect 22293 10557 22327 10591
rect 26525 10557 26559 10591
rect 9229 10421 9263 10455
rect 11069 10421 11103 10455
rect 12449 10421 12483 10455
rect 14565 10421 14599 10455
rect 5549 10217 5583 10251
rect 11529 10217 11563 10251
rect 12541 10217 12575 10251
rect 14289 10217 14323 10251
rect 21281 10217 21315 10251
rect 28457 10217 28491 10251
rect 29745 10217 29779 10251
rect 29929 10149 29963 10183
rect 8217 10081 8251 10115
rect 9781 10081 9815 10115
rect 10057 10081 10091 10115
rect 13001 10081 13035 10115
rect 14749 10081 14783 10115
rect 14933 10081 14967 10115
rect 17141 10081 17175 10115
rect 17877 10081 17911 10115
rect 25513 10081 25547 10115
rect 8033 10013 8067 10047
rect 12909 10013 12943 10047
rect 14657 10013 14691 10047
rect 22569 10013 22603 10047
rect 25329 10013 25363 10047
rect 28089 10013 28123 10047
rect 28181 10013 28215 10047
rect 28917 10013 28951 10047
rect 7021 9945 7055 9979
rect 27905 9945 27939 9979
rect 28273 9945 28307 9979
rect 30205 9945 30239 9979
rect 7665 9877 7699 9911
rect 8125 9877 8159 9911
rect 24961 9877 24995 9911
rect 25421 9877 25455 9911
rect 29009 9877 29043 9911
rect 8401 9673 8435 9707
rect 26065 9673 26099 9707
rect 27997 9673 28031 9707
rect 4813 9605 4847 9639
rect 7288 9605 7322 9639
rect 10977 9605 11011 9639
rect 15209 9605 15243 9639
rect 24593 9605 24627 9639
rect 29110 9605 29144 9639
rect 30113 9605 30147 9639
rect 5641 9537 5675 9571
rect 7021 9537 7055 9571
rect 9965 9537 9999 9571
rect 10149 9537 10183 9571
rect 12081 9537 12115 9571
rect 16957 9537 16991 9571
rect 22017 9537 22051 9571
rect 22284 9537 22318 9571
rect 24317 9537 24351 9571
rect 29837 9537 29871 9571
rect 5549 9469 5583 9503
rect 11989 9469 12023 9503
rect 12449 9469 12483 9503
rect 15301 9469 15335 9503
rect 15393 9469 15427 9503
rect 17877 9469 17911 9503
rect 29377 9469 29411 9503
rect 14841 9333 14875 9367
rect 23397 9333 23431 9367
rect 9689 9129 9723 9163
rect 14473 9129 14507 9163
rect 22845 9129 22879 9163
rect 24685 9129 24719 9163
rect 29837 9129 29871 9163
rect 9229 8993 9263 9027
rect 30021 8993 30055 9027
rect 7941 8925 7975 8959
rect 8217 8925 8251 8959
rect 9321 8925 9355 8959
rect 13185 8925 13219 8959
rect 15586 8925 15620 8959
rect 15853 8925 15887 8959
rect 19901 8925 19935 8959
rect 20085 8925 20119 8959
rect 22937 8925 22971 8959
rect 24593 8925 24627 8959
rect 24777 8925 24811 8959
rect 28089 8925 28123 8959
rect 28273 8925 28307 8959
rect 28917 8925 28951 8959
rect 29101 8925 29135 8959
rect 30113 8925 30147 8959
rect 13001 8857 13035 8891
rect 27721 8857 27755 8891
rect 28733 8857 28767 8891
rect 8585 8789 8619 8823
rect 13369 8789 13403 8823
rect 19993 8789 20027 8823
rect 27905 8789 27939 8823
rect 27997 8789 28031 8823
rect 8309 8585 8343 8619
rect 12909 8585 12943 8619
rect 18613 8585 18647 8619
rect 25237 8585 25271 8619
rect 28641 8585 28675 8619
rect 9597 8517 9631 8551
rect 12357 8517 12391 8551
rect 13185 8517 13219 8551
rect 13277 8517 13311 8551
rect 14013 8517 14047 8551
rect 27813 8517 27847 8551
rect 5825 8449 5859 8483
rect 6561 8449 6595 8483
rect 11161 8449 11195 8483
rect 12265 8449 12299 8483
rect 12449 8449 12483 8483
rect 13093 8449 13127 8483
rect 13461 8449 13495 8483
rect 13921 8449 13955 8483
rect 14105 8449 14139 8483
rect 19073 8449 19107 8483
rect 19441 8449 19475 8483
rect 22017 8449 22051 8483
rect 22201 8449 22235 8483
rect 23857 8449 23891 8483
rect 24113 8449 24147 8483
rect 27629 8449 27663 8483
rect 27905 8449 27939 8483
rect 28033 8449 28067 8483
rect 28549 8449 28583 8483
rect 16865 8381 16899 8415
rect 17141 8381 17175 8415
rect 27813 8381 27847 8415
rect 6653 8313 6687 8347
rect 5733 8245 5767 8279
rect 11069 8245 11103 8279
rect 20867 8245 20901 8279
rect 22109 8245 22143 8279
rect 12541 8041 12575 8075
rect 13093 8041 13127 8075
rect 16221 8041 16255 8075
rect 16819 8041 16853 8075
rect 19533 8041 19567 8075
rect 25973 8041 26007 8075
rect 5365 7905 5399 7939
rect 11069 7905 11103 7939
rect 18613 7905 18647 7939
rect 20821 7905 20855 7939
rect 7665 7837 7699 7871
rect 9321 7837 9355 7871
rect 10793 7837 10827 7871
rect 13461 7837 13495 7871
rect 15945 7837 15979 7871
rect 18245 7837 18279 7871
rect 19441 7837 19475 7871
rect 19625 7837 19659 7871
rect 20545 7837 20579 7871
rect 24593 7837 24627 7871
rect 28549 7837 28583 7871
rect 5641 7769 5675 7803
rect 13277 7769 13311 7803
rect 24838 7769 24872 7803
rect 7113 7701 7147 7735
rect 7757 7701 7791 7735
rect 9229 7701 9263 7735
rect 22293 7701 22327 7735
rect 28457 7701 28491 7735
rect 6009 7497 6043 7531
rect 6653 7497 6687 7531
rect 10793 7497 10827 7531
rect 11713 7497 11747 7531
rect 18613 7497 18647 7531
rect 29469 7497 29503 7531
rect 8033 7429 8067 7463
rect 16221 7429 16255 7463
rect 28356 7429 28390 7463
rect 5365 7361 5399 7395
rect 5457 7361 5491 7395
rect 6745 7361 6779 7395
rect 7757 7361 7791 7395
rect 10701 7361 10735 7395
rect 12541 7361 12575 7395
rect 16129 7361 16163 7395
rect 16313 7361 16347 7395
rect 16865 7361 16899 7395
rect 21281 7361 21315 7395
rect 21465 7361 21499 7395
rect 22017 7361 22051 7395
rect 22201 7361 22235 7395
rect 22661 7361 22695 7395
rect 22845 7361 22879 7395
rect 25421 7361 25455 7395
rect 27629 7361 27663 7395
rect 9505 7293 9539 7327
rect 12449 7293 12483 7327
rect 17141 7293 17175 7327
rect 27537 7293 27571 7327
rect 28089 7293 28123 7327
rect 21373 7157 21407 7191
rect 22109 7157 22143 7191
rect 22753 7157 22787 7191
rect 25329 7157 25363 7191
rect 6941 6953 6975 6987
rect 25973 6953 26007 6987
rect 5457 6817 5491 6851
rect 8493 6817 8527 6851
rect 9137 6817 9171 6851
rect 16083 6817 16117 6851
rect 17601 6817 17635 6851
rect 20453 6817 20487 6851
rect 20821 6817 20855 6851
rect 26893 6817 26927 6851
rect 29101 6817 29135 6851
rect 7205 6749 7239 6783
rect 8585 6749 8619 6783
rect 14289 6749 14323 6783
rect 14657 6749 14691 6783
rect 16589 6749 16623 6783
rect 16865 6749 16899 6783
rect 17509 6749 17543 6783
rect 17693 6749 17727 6783
rect 24593 6749 24627 6783
rect 24860 6749 24894 6783
rect 27169 6749 27203 6783
rect 27445 6749 27479 6783
rect 28825 6749 28859 6783
rect 28917 6749 28951 6783
rect 9413 6681 9447 6715
rect 27077 6681 27111 6715
rect 10885 6613 10919 6647
rect 22247 6613 22281 6647
rect 27261 6613 27295 6647
rect 28457 6613 28491 6647
rect 6009 6409 6043 6443
rect 6653 6409 6687 6443
rect 8401 6409 8435 6443
rect 10057 6409 10091 6443
rect 28549 6409 28583 6443
rect 5273 6273 5307 6307
rect 5457 6273 5491 6307
rect 6745 6273 6779 6307
rect 8309 6273 8343 6307
rect 9413 6273 9447 6307
rect 9505 6273 9539 6307
rect 10977 6273 11011 6307
rect 13553 6273 13587 6307
rect 22385 6273 22419 6307
rect 24317 6273 24351 6307
rect 24573 6273 24607 6307
rect 26433 6273 26467 6307
rect 27436 6273 27470 6307
rect 29285 6273 29319 6307
rect 30113 6273 30147 6307
rect 30297 6273 30331 6307
rect 11069 6205 11103 6239
rect 13277 6205 13311 6239
rect 22017 6205 22051 6239
rect 26525 6205 26559 6239
rect 27169 6205 27203 6239
rect 29377 6205 29411 6239
rect 30205 6205 30239 6239
rect 11805 6137 11839 6171
rect 23811 6069 23845 6103
rect 25697 6069 25731 6103
rect 29561 6069 29595 6103
rect 14289 5865 14323 5899
rect 28549 5865 28583 5899
rect 29101 5865 29135 5899
rect 12081 5729 12115 5763
rect 15669 5729 15703 5763
rect 19717 5729 19751 5763
rect 19993 5729 20027 5763
rect 21465 5729 21499 5763
rect 21741 5729 21775 5763
rect 24593 5729 24627 5763
rect 27537 5729 27571 5763
rect 30113 5729 30147 5763
rect 11345 5661 11379 5695
rect 11805 5661 11839 5695
rect 19625 5661 19659 5695
rect 26709 5661 26743 5695
rect 27077 5661 27111 5695
rect 27261 5661 27295 5695
rect 27445 5661 27479 5695
rect 27997 5661 28031 5695
rect 28273 5661 28307 5695
rect 28365 5661 28399 5695
rect 29009 5661 29043 5695
rect 29837 5661 29871 5695
rect 15424 5593 15458 5627
rect 24838 5593 24872 5627
rect 28181 5593 28215 5627
rect 23213 5525 23247 5559
rect 25973 5525 26007 5559
rect 18337 5321 18371 5355
rect 20177 5321 20211 5355
rect 27629 5321 27663 5355
rect 19042 5253 19076 5287
rect 27537 5253 27571 5287
rect 14125 5185 14159 5219
rect 16957 5185 16991 5219
rect 17224 5185 17258 5219
rect 18797 5185 18831 5219
rect 27445 5185 27479 5219
rect 27813 5185 27847 5219
rect 28733 5185 28767 5219
rect 28917 5185 28951 5219
rect 14381 5117 14415 5151
rect 27721 5049 27755 5083
rect 13001 4981 13035 5015
rect 28733 4981 28767 5015
rect 17233 4777 17267 4811
rect 19441 4777 19475 4811
rect 16773 4709 16807 4743
rect 14657 4641 14691 4675
rect 14933 4641 14967 4675
rect 17509 4641 17543 4675
rect 20821 4641 20855 4675
rect 14565 4573 14599 4607
rect 15393 4573 15427 4607
rect 15649 4573 15683 4607
rect 17601 4573 17635 4607
rect 20554 4573 20588 4607
rect 15117 4233 15151 4267
rect 13737 4097 13771 4131
rect 14004 4097 14038 4131
rect 29837 2397 29871 2431
rect 30113 2329 30147 2363
<< metal1 >>
rect 1104 29402 30976 29424
rect 1104 29350 8378 29402
rect 8430 29350 8442 29402
rect 8494 29350 8506 29402
rect 8558 29350 8570 29402
rect 8622 29350 8634 29402
rect 8686 29350 15806 29402
rect 15858 29350 15870 29402
rect 15922 29350 15934 29402
rect 15986 29350 15998 29402
rect 16050 29350 16062 29402
rect 16114 29350 23234 29402
rect 23286 29350 23298 29402
rect 23350 29350 23362 29402
rect 23414 29350 23426 29402
rect 23478 29350 23490 29402
rect 23542 29350 30662 29402
rect 30714 29350 30726 29402
rect 30778 29350 30790 29402
rect 30842 29350 30854 29402
rect 30906 29350 30918 29402
rect 30970 29350 30976 29402
rect 1104 29328 30976 29350
rect 6086 29180 6092 29232
rect 6144 29220 6150 29232
rect 6641 29223 6699 29229
rect 6641 29220 6653 29223
rect 6144 29192 6653 29220
rect 6144 29180 6150 29192
rect 6641 29189 6653 29192
rect 6687 29189 6699 29223
rect 6641 29183 6699 29189
rect 10781 29223 10839 29229
rect 10781 29189 10793 29223
rect 10827 29220 10839 29223
rect 15378 29220 15384 29232
rect 10827 29192 15384 29220
rect 10827 29189 10839 29192
rect 10781 29183 10839 29189
rect 15378 29180 15384 29192
rect 15436 29180 15442 29232
rect 18138 29180 18144 29232
rect 18196 29180 18202 29232
rect 30101 29223 30159 29229
rect 30101 29189 30113 29223
rect 30147 29220 30159 29223
rect 31018 29220 31024 29232
rect 30147 29192 31024 29220
rect 30147 29189 30159 29192
rect 30101 29183 30159 29189
rect 31018 29180 31024 29192
rect 31076 29180 31082 29232
rect 3145 29155 3203 29161
rect 3145 29121 3157 29155
rect 3191 29152 3203 29155
rect 3234 29152 3240 29164
rect 3191 29124 3240 29152
rect 3191 29121 3203 29124
rect 3145 29115 3203 29121
rect 3234 29112 3240 29124
rect 3292 29112 3298 29164
rect 3329 29155 3387 29161
rect 3329 29121 3341 29155
rect 3375 29121 3387 29155
rect 3329 29115 3387 29121
rect 3050 29044 3056 29096
rect 3108 29084 3114 29096
rect 3344 29084 3372 29115
rect 10226 29112 10232 29164
rect 10284 29112 10290 29164
rect 13998 29112 14004 29164
rect 14056 29152 14062 29164
rect 14369 29155 14427 29161
rect 14369 29152 14381 29155
rect 14056 29124 14381 29152
rect 14056 29112 14062 29124
rect 14369 29121 14381 29124
rect 14415 29121 14427 29155
rect 14369 29115 14427 29121
rect 22002 29112 22008 29164
rect 22060 29112 22066 29164
rect 25958 29112 25964 29164
rect 26016 29112 26022 29164
rect 29089 29155 29147 29161
rect 29089 29121 29101 29155
rect 29135 29152 29147 29155
rect 29730 29152 29736 29164
rect 29135 29124 29736 29152
rect 29135 29121 29147 29124
rect 29089 29115 29147 29121
rect 29730 29112 29736 29124
rect 29788 29112 29794 29164
rect 29825 29155 29883 29161
rect 29825 29121 29837 29155
rect 29871 29121 29883 29155
rect 29825 29115 29883 29121
rect 3108 29056 3372 29084
rect 3108 29044 3114 29056
rect 14458 29044 14464 29096
rect 14516 29084 14522 29096
rect 14645 29087 14703 29093
rect 14645 29084 14657 29087
rect 14516 29056 14657 29084
rect 14516 29044 14522 29056
rect 14645 29053 14657 29056
rect 14691 29053 14703 29087
rect 14645 29047 14703 29053
rect 28534 29044 28540 29096
rect 28592 29044 28598 29096
rect 28994 29044 29000 29096
rect 29052 29084 29058 29096
rect 29840 29084 29868 29115
rect 29052 29056 29868 29084
rect 29052 29044 29058 29056
rect 3329 29019 3387 29025
rect 3329 28985 3341 29019
rect 3375 29016 3387 29019
rect 4522 29016 4528 29028
rect 3375 28988 4528 29016
rect 3375 28985 3387 28988
rect 3329 28979 3387 28985
rect 4522 28976 4528 28988
rect 4580 28976 4586 29028
rect 6917 29019 6975 29025
rect 6917 28985 6929 29019
rect 6963 29016 6975 29019
rect 7190 29016 7196 29028
rect 6963 28988 7196 29016
rect 6963 28985 6975 28988
rect 6917 28979 6975 28985
rect 7190 28976 7196 28988
rect 7248 28976 7254 29028
rect 22186 28976 22192 29028
rect 22244 28976 22250 29028
rect 25682 28976 25688 29028
rect 25740 29016 25746 29028
rect 26145 29019 26203 29025
rect 26145 29016 26157 29019
rect 25740 28988 26157 29016
rect 25740 28976 25746 28988
rect 26145 28985 26157 28988
rect 26191 28985 26203 29019
rect 26145 28979 26203 28985
rect 18138 28908 18144 28960
rect 18196 28948 18202 28960
rect 18233 28951 18291 28957
rect 18233 28948 18245 28951
rect 18196 28920 18245 28948
rect 18196 28908 18202 28920
rect 18233 28917 18245 28920
rect 18279 28917 18291 28951
rect 18233 28911 18291 28917
rect 1104 28858 30820 28880
rect 1104 28806 4664 28858
rect 4716 28806 4728 28858
rect 4780 28806 4792 28858
rect 4844 28806 4856 28858
rect 4908 28806 4920 28858
rect 4972 28806 12092 28858
rect 12144 28806 12156 28858
rect 12208 28806 12220 28858
rect 12272 28806 12284 28858
rect 12336 28806 12348 28858
rect 12400 28806 19520 28858
rect 19572 28806 19584 28858
rect 19636 28806 19648 28858
rect 19700 28806 19712 28858
rect 19764 28806 19776 28858
rect 19828 28806 26948 28858
rect 27000 28806 27012 28858
rect 27064 28806 27076 28858
rect 27128 28806 27140 28858
rect 27192 28806 27204 28858
rect 27256 28806 30820 28858
rect 1104 28784 30820 28806
rect 2130 28704 2136 28756
rect 2188 28744 2194 28756
rect 3510 28744 3516 28756
rect 2188 28716 3516 28744
rect 2188 28704 2194 28716
rect 3510 28704 3516 28716
rect 3568 28704 3574 28756
rect 3142 28636 3148 28688
rect 3200 28636 3206 28688
rect 11704 28552 11756 28558
rect 3234 28500 3240 28552
rect 3292 28540 3298 28552
rect 3329 28543 3387 28549
rect 3329 28540 3341 28543
rect 3292 28512 3341 28540
rect 3292 28500 3298 28512
rect 3329 28509 3341 28512
rect 3375 28509 3387 28543
rect 3329 28503 3387 28509
rect 3421 28543 3479 28549
rect 3421 28509 3433 28543
rect 3467 28540 3479 28543
rect 3878 28540 3884 28552
rect 3467 28512 3884 28540
rect 3467 28509 3479 28512
rect 3421 28503 3479 28509
rect 3878 28500 3884 28512
rect 3936 28500 3942 28552
rect 4985 28543 5043 28549
rect 4985 28509 4997 28543
rect 5031 28540 5043 28543
rect 7190 28540 7196 28552
rect 5031 28512 7196 28540
rect 5031 28509 5043 28512
rect 4985 28503 5043 28509
rect 7190 28500 7196 28512
rect 7248 28500 7254 28552
rect 7745 28543 7803 28549
rect 7745 28509 7757 28543
rect 7791 28540 7803 28543
rect 8205 28543 8263 28549
rect 8205 28540 8217 28543
rect 7791 28512 8217 28540
rect 7791 28509 7803 28512
rect 7745 28503 7803 28509
rect 8205 28509 8217 28512
rect 8251 28540 8263 28543
rect 8754 28540 8760 28552
rect 8251 28512 8760 28540
rect 8251 28509 8263 28512
rect 8205 28503 8263 28509
rect 8754 28500 8760 28512
rect 8812 28500 8818 28552
rect 9585 28543 9643 28549
rect 9585 28509 9597 28543
rect 9631 28540 9643 28543
rect 10318 28540 10324 28552
rect 9631 28512 10324 28540
rect 9631 28509 9643 28512
rect 9585 28503 9643 28509
rect 10318 28500 10324 28512
rect 10376 28500 10382 28552
rect 11054 28500 11060 28552
rect 11112 28500 11118 28552
rect 12529 28543 12587 28549
rect 12529 28509 12541 28543
rect 12575 28540 12587 28543
rect 12710 28540 12716 28552
rect 12575 28512 12716 28540
rect 12575 28509 12587 28512
rect 12529 28503 12587 28509
rect 12710 28500 12716 28512
rect 12768 28500 12774 28552
rect 13722 28500 13728 28552
rect 13780 28540 13786 28552
rect 14645 28543 14703 28549
rect 14645 28540 14657 28543
rect 13780 28512 14657 28540
rect 13780 28500 13786 28512
rect 14645 28509 14657 28512
rect 14691 28509 14703 28543
rect 14645 28503 14703 28509
rect 14918 28500 14924 28552
rect 14976 28540 14982 28552
rect 15289 28543 15347 28549
rect 15289 28540 15301 28543
rect 14976 28512 15301 28540
rect 14976 28500 14982 28512
rect 15289 28509 15301 28512
rect 15335 28509 15347 28543
rect 15289 28503 15347 28509
rect 18138 28500 18144 28552
rect 18196 28540 18202 28552
rect 18325 28543 18383 28549
rect 18325 28540 18337 28543
rect 18196 28512 18337 28540
rect 18196 28500 18202 28512
rect 18325 28509 18337 28512
rect 18371 28509 18383 28543
rect 18325 28503 18383 28509
rect 20714 28500 20720 28552
rect 20772 28540 20778 28552
rect 20809 28543 20867 28549
rect 20809 28540 20821 28543
rect 20772 28512 20821 28540
rect 20772 28500 20778 28512
rect 20809 28509 20821 28512
rect 20855 28509 20867 28543
rect 20809 28503 20867 28509
rect 21729 28543 21787 28549
rect 21729 28509 21741 28543
rect 21775 28509 21787 28543
rect 21729 28503 21787 28509
rect 11704 28494 11756 28500
rect 3050 28432 3056 28484
rect 3108 28472 3114 28484
rect 3145 28475 3203 28481
rect 3145 28472 3157 28475
rect 3108 28444 3157 28472
rect 3108 28432 3114 28444
rect 3145 28441 3157 28444
rect 3191 28472 3203 28475
rect 4157 28475 4215 28481
rect 4157 28472 4169 28475
rect 3191 28444 4169 28472
rect 3191 28441 3203 28444
rect 3145 28435 3203 28441
rect 4157 28441 4169 28444
rect 4203 28441 4215 28475
rect 4157 28435 4215 28441
rect 11790 28432 11796 28484
rect 11848 28432 11854 28484
rect 21744 28472 21772 28503
rect 21818 28500 21824 28552
rect 21876 28540 21882 28552
rect 22741 28543 22799 28549
rect 22741 28540 22753 28543
rect 21876 28512 22753 28540
rect 21876 28500 21882 28512
rect 22741 28509 22753 28512
rect 22787 28509 22799 28543
rect 22741 28503 22799 28509
rect 22830 28500 22836 28552
rect 22888 28540 22894 28552
rect 22925 28543 22983 28549
rect 22925 28540 22937 28543
rect 22888 28512 22937 28540
rect 22888 28500 22894 28512
rect 22925 28509 22937 28512
rect 22971 28509 22983 28543
rect 22925 28503 22983 28509
rect 26418 28500 26424 28552
rect 26476 28540 26482 28552
rect 27065 28543 27123 28549
rect 27065 28540 27077 28543
rect 26476 28512 27077 28540
rect 26476 28500 26482 28512
rect 27065 28509 27077 28512
rect 27111 28509 27123 28543
rect 27065 28503 27123 28509
rect 27890 28500 27896 28552
rect 27948 28540 27954 28552
rect 28169 28543 28227 28549
rect 28169 28540 28181 28543
rect 27948 28512 28181 28540
rect 27948 28500 27954 28512
rect 28169 28509 28181 28512
rect 28215 28509 28227 28543
rect 28169 28503 28227 28509
rect 28353 28543 28411 28549
rect 28353 28509 28365 28543
rect 28399 28509 28411 28543
rect 28353 28503 28411 28509
rect 23566 28472 23572 28484
rect 21744 28444 23572 28472
rect 23566 28432 23572 28444
rect 23624 28432 23630 28484
rect 27614 28432 27620 28484
rect 27672 28472 27678 28484
rect 28368 28472 28396 28503
rect 27672 28444 28396 28472
rect 27672 28432 27678 28444
rect 7006 28364 7012 28416
rect 7064 28404 7070 28416
rect 7653 28407 7711 28413
rect 7653 28404 7665 28407
rect 7064 28376 7665 28404
rect 7064 28364 7070 28376
rect 7653 28373 7665 28376
rect 7699 28373 7711 28407
rect 7653 28367 7711 28373
rect 8294 28364 8300 28416
rect 8352 28364 8358 28416
rect 8846 28364 8852 28416
rect 8904 28404 8910 28416
rect 9493 28407 9551 28413
rect 9493 28404 9505 28407
rect 8904 28376 9505 28404
rect 8904 28364 8910 28376
rect 9493 28373 9505 28376
rect 9539 28373 9551 28407
rect 9493 28367 9551 28373
rect 10413 28407 10471 28413
rect 10413 28373 10425 28407
rect 10459 28404 10471 28407
rect 10870 28404 10876 28416
rect 10459 28376 10876 28404
rect 10459 28373 10471 28376
rect 10413 28367 10471 28373
rect 10870 28364 10876 28376
rect 10928 28364 10934 28416
rect 12066 28364 12072 28416
rect 12124 28404 12130 28416
rect 12621 28407 12679 28413
rect 12621 28404 12633 28407
rect 12124 28376 12633 28404
rect 12124 28364 12130 28376
rect 12621 28373 12633 28376
rect 12667 28373 12679 28407
rect 12621 28367 12679 28373
rect 14737 28407 14795 28413
rect 14737 28373 14749 28407
rect 14783 28404 14795 28407
rect 15286 28404 15292 28416
rect 14783 28376 15292 28404
rect 14783 28373 14795 28376
rect 14737 28367 14795 28373
rect 15286 28364 15292 28376
rect 15344 28364 15350 28416
rect 15381 28407 15439 28413
rect 15381 28373 15393 28407
rect 15427 28404 15439 28407
rect 16206 28404 16212 28416
rect 15427 28376 16212 28404
rect 15427 28373 15439 28376
rect 15381 28367 15439 28373
rect 16206 28364 16212 28376
rect 16264 28364 16270 28416
rect 18509 28407 18567 28413
rect 18509 28373 18521 28407
rect 18555 28404 18567 28407
rect 18598 28404 18604 28416
rect 18555 28376 18604 28404
rect 18555 28373 18567 28376
rect 18509 28367 18567 28373
rect 18598 28364 18604 28376
rect 18656 28364 18662 28416
rect 20898 28364 20904 28416
rect 20956 28364 20962 28416
rect 21637 28407 21695 28413
rect 21637 28373 21649 28407
rect 21683 28404 21695 28407
rect 22370 28404 22376 28416
rect 21683 28376 22376 28404
rect 21683 28373 21695 28376
rect 21637 28367 21695 28373
rect 22370 28364 22376 28376
rect 22428 28364 22434 28416
rect 23750 28364 23756 28416
rect 23808 28364 23814 28416
rect 27157 28407 27215 28413
rect 27157 28373 27169 28407
rect 27203 28404 27215 28407
rect 27430 28404 27436 28416
rect 27203 28376 27436 28404
rect 27203 28373 27215 28376
rect 27157 28367 27215 28373
rect 27430 28364 27436 28376
rect 27488 28364 27494 28416
rect 29178 28364 29184 28416
rect 29236 28364 29242 28416
rect 1104 28314 30976 28336
rect 1104 28262 8378 28314
rect 8430 28262 8442 28314
rect 8494 28262 8506 28314
rect 8558 28262 8570 28314
rect 8622 28262 8634 28314
rect 8686 28262 15806 28314
rect 15858 28262 15870 28314
rect 15922 28262 15934 28314
rect 15986 28262 15998 28314
rect 16050 28262 16062 28314
rect 16114 28262 23234 28314
rect 23286 28262 23298 28314
rect 23350 28262 23362 28314
rect 23414 28262 23426 28314
rect 23478 28262 23490 28314
rect 23542 28262 30662 28314
rect 30714 28262 30726 28314
rect 30778 28262 30790 28314
rect 30842 28262 30854 28314
rect 30906 28262 30918 28314
rect 30970 28262 30976 28314
rect 1104 28240 30976 28262
rect 12710 28160 12716 28212
rect 12768 28160 12774 28212
rect 13814 28160 13820 28212
rect 13872 28200 13878 28212
rect 14918 28200 14924 28212
rect 13872 28172 14924 28200
rect 13872 28160 13878 28172
rect 14918 28160 14924 28172
rect 14976 28160 14982 28212
rect 15286 28160 15292 28212
rect 15344 28200 15350 28212
rect 18141 28203 18199 28209
rect 18141 28200 18153 28203
rect 15344 28172 15976 28200
rect 15344 28160 15350 28172
rect 2866 28132 2872 28144
rect 2700 28104 2872 28132
rect 2700 28005 2728 28104
rect 2866 28092 2872 28104
rect 2924 28132 2930 28144
rect 2924 28104 4016 28132
rect 2924 28092 2930 28104
rect 2958 28073 2964 28076
rect 2952 28027 2964 28073
rect 2958 28024 2964 28027
rect 3016 28024 3022 28076
rect 3988 28008 4016 28104
rect 4522 28092 4528 28144
rect 4580 28132 4586 28144
rect 4770 28135 4828 28141
rect 4770 28132 4782 28135
rect 4580 28104 4782 28132
rect 4580 28092 4586 28104
rect 4770 28101 4782 28104
rect 4816 28101 4828 28135
rect 4770 28095 4828 28101
rect 8573 28135 8631 28141
rect 8573 28101 8585 28135
rect 8619 28132 8631 28135
rect 8846 28132 8852 28144
rect 8619 28104 8852 28132
rect 8619 28101 8631 28104
rect 8573 28095 8631 28101
rect 8846 28092 8852 28104
rect 8904 28092 8910 28144
rect 12728 28132 12756 28160
rect 11164 28104 12756 28132
rect 6920 28076 6972 28082
rect 8294 28024 8300 28076
rect 8352 28024 8358 28076
rect 9674 28024 9680 28076
rect 9732 28024 9738 28076
rect 11164 28073 11192 28104
rect 13354 28092 13360 28144
rect 13412 28092 13418 28144
rect 15470 28092 15476 28144
rect 15528 28092 15534 28144
rect 15948 28141 15976 28172
rect 17604 28172 18153 28200
rect 15933 28135 15991 28141
rect 15933 28101 15945 28135
rect 15979 28101 15991 28135
rect 15933 28095 15991 28101
rect 11149 28067 11207 28073
rect 11149 28033 11161 28067
rect 11195 28033 11207 28067
rect 11149 28027 11207 28033
rect 12066 28024 12072 28076
rect 12124 28024 12130 28076
rect 16206 28024 16212 28076
rect 16264 28024 16270 28076
rect 17604 28073 17632 28172
rect 18141 28169 18153 28172
rect 18187 28200 18199 28203
rect 18782 28200 18788 28212
rect 18187 28172 18788 28200
rect 18187 28169 18199 28172
rect 18141 28163 18199 28169
rect 18782 28160 18788 28172
rect 18840 28160 18846 28212
rect 23566 28160 23572 28212
rect 23624 28200 23630 28212
rect 24213 28203 24271 28209
rect 24213 28200 24225 28203
rect 23624 28172 24225 28200
rect 23624 28160 23630 28172
rect 24213 28169 24225 28172
rect 24259 28169 24271 28203
rect 24213 28163 24271 28169
rect 18874 28092 18880 28144
rect 18932 28092 18938 28144
rect 23750 28092 23756 28144
rect 23808 28092 23814 28144
rect 27430 28092 27436 28144
rect 27488 28092 27494 28144
rect 28166 28092 28172 28144
rect 28224 28092 28230 28144
rect 17589 28067 17647 28073
rect 17589 28033 17601 28067
rect 17635 28033 17647 28067
rect 17589 28027 17647 28033
rect 20806 28024 20812 28076
rect 20864 28024 20870 28076
rect 21082 28024 21088 28076
rect 21140 28064 21146 28076
rect 21818 28064 21824 28076
rect 21140 28036 21824 28064
rect 21140 28024 21146 28036
rect 21818 28024 21824 28036
rect 21876 28024 21882 28076
rect 29454 28024 29460 28076
rect 29512 28024 29518 28076
rect 6920 28018 6972 28024
rect 2685 27999 2743 28005
rect 2685 27965 2697 27999
rect 2731 27965 2743 27999
rect 2685 27959 2743 27965
rect 3970 27956 3976 28008
rect 4028 27996 4034 28008
rect 4525 27999 4583 28005
rect 4525 27996 4537 27999
rect 4028 27968 4537 27996
rect 4028 27956 4034 27968
rect 4525 27965 4537 27968
rect 4571 27965 4583 27999
rect 4525 27959 4583 27965
rect 7009 27999 7067 28005
rect 7009 27965 7021 27999
rect 7055 27996 7067 27999
rect 7374 27996 7380 28008
rect 7055 27968 7380 27996
rect 7055 27965 7067 27968
rect 7009 27959 7067 27965
rect 7374 27956 7380 27968
rect 7432 27956 7438 28008
rect 7650 27956 7656 28008
rect 7708 27996 7714 28008
rect 7745 27999 7803 28005
rect 7745 27996 7757 27999
rect 7708 27968 7757 27996
rect 7708 27956 7714 27968
rect 7745 27965 7757 27968
rect 7791 27965 7803 27999
rect 7745 27959 7803 27965
rect 12345 27999 12403 28005
rect 12345 27965 12357 27999
rect 12391 27996 12403 27999
rect 13630 27996 13636 28008
rect 12391 27968 13636 27996
rect 12391 27965 12403 27968
rect 12345 27959 12403 27965
rect 13630 27956 13636 27968
rect 13688 27956 13694 28008
rect 17497 27999 17555 28005
rect 17497 27965 17509 27999
rect 17543 27996 17555 27999
rect 19613 27999 19671 28005
rect 19613 27996 19625 27999
rect 17543 27968 19625 27996
rect 17543 27965 17555 27968
rect 17497 27959 17555 27965
rect 19613 27965 19625 27968
rect 19659 27965 19671 27999
rect 19613 27959 19671 27965
rect 19886 27956 19892 28008
rect 19944 27956 19950 28008
rect 21358 27956 21364 28008
rect 21416 27956 21422 28008
rect 22465 27999 22523 28005
rect 22465 27965 22477 27999
rect 22511 27965 22523 27999
rect 22465 27959 22523 27965
rect 10045 27931 10103 27937
rect 10045 27897 10057 27931
rect 10091 27928 10103 27931
rect 10318 27928 10324 27940
rect 10091 27900 10324 27928
rect 10091 27897 10103 27900
rect 10045 27891 10103 27897
rect 10318 27888 10324 27900
rect 10376 27928 10382 27940
rect 11882 27928 11888 27940
rect 10376 27900 11888 27928
rect 10376 27888 10382 27900
rect 11882 27888 11888 27900
rect 11940 27888 11946 27940
rect 13722 27888 13728 27940
rect 13780 27928 13786 27940
rect 14461 27931 14519 27937
rect 14461 27928 14473 27931
rect 13780 27900 14473 27928
rect 13780 27888 13786 27900
rect 14461 27897 14473 27900
rect 14507 27897 14519 27931
rect 14461 27891 14519 27897
rect 3878 27820 3884 27872
rect 3936 27860 3942 27872
rect 4065 27863 4123 27869
rect 4065 27860 4077 27863
rect 3936 27832 4077 27860
rect 3936 27820 3942 27832
rect 4065 27829 4077 27832
rect 4111 27829 4123 27863
rect 4065 27823 4123 27829
rect 5902 27820 5908 27872
rect 5960 27820 5966 27872
rect 11057 27863 11115 27869
rect 11057 27829 11069 27863
rect 11103 27860 11115 27863
rect 11146 27860 11152 27872
rect 11103 27832 11152 27860
rect 11103 27829 11115 27832
rect 11057 27823 11115 27829
rect 11146 27820 11152 27832
rect 11204 27820 11210 27872
rect 22480 27860 22508 27959
rect 22738 27956 22744 28008
rect 22796 27956 22802 28008
rect 26602 27956 26608 28008
rect 26660 27996 26666 28008
rect 27157 27999 27215 28005
rect 27157 27996 27169 27999
rect 26660 27968 27169 27996
rect 26660 27956 26666 27968
rect 27157 27965 27169 27968
rect 27203 27965 27215 27999
rect 27157 27959 27215 27965
rect 23474 27860 23480 27872
rect 22480 27832 23480 27860
rect 23474 27820 23480 27832
rect 23532 27820 23538 27872
rect 28902 27820 28908 27872
rect 28960 27820 28966 27872
rect 29549 27863 29607 27869
rect 29549 27829 29561 27863
rect 29595 27860 29607 27863
rect 29914 27860 29920 27872
rect 29595 27832 29920 27860
rect 29595 27829 29607 27832
rect 29549 27823 29607 27829
rect 29914 27820 29920 27832
rect 29972 27820 29978 27872
rect 1104 27770 30820 27792
rect 1104 27718 4664 27770
rect 4716 27718 4728 27770
rect 4780 27718 4792 27770
rect 4844 27718 4856 27770
rect 4908 27718 4920 27770
rect 4972 27718 12092 27770
rect 12144 27718 12156 27770
rect 12208 27718 12220 27770
rect 12272 27718 12284 27770
rect 12336 27718 12348 27770
rect 12400 27718 19520 27770
rect 19572 27718 19584 27770
rect 19636 27718 19648 27770
rect 19700 27718 19712 27770
rect 19764 27718 19776 27770
rect 19828 27718 26948 27770
rect 27000 27718 27012 27770
rect 27064 27718 27076 27770
rect 27128 27718 27140 27770
rect 27192 27718 27204 27770
rect 27256 27718 30820 27770
rect 1104 27696 30820 27718
rect 2317 27659 2375 27665
rect 2317 27625 2329 27659
rect 2363 27656 2375 27659
rect 2363 27628 2774 27656
rect 2363 27625 2375 27628
rect 2317 27619 2375 27625
rect 2746 27588 2774 27628
rect 2958 27616 2964 27668
rect 3016 27616 3022 27668
rect 3329 27659 3387 27665
rect 3329 27625 3341 27659
rect 3375 27656 3387 27659
rect 3878 27656 3884 27668
rect 3375 27628 3884 27656
rect 3375 27625 3387 27628
rect 3329 27619 3387 27625
rect 3344 27588 3372 27619
rect 3878 27616 3884 27628
rect 3936 27656 3942 27668
rect 6904 27659 6962 27665
rect 3936 27628 4936 27656
rect 3936 27616 3942 27628
rect 2746 27560 3372 27588
rect 4908 27588 4936 27628
rect 6904 27625 6916 27659
rect 6950 27656 6962 27659
rect 7006 27656 7012 27668
rect 6950 27628 7012 27656
rect 6950 27625 6962 27628
rect 6904 27619 6962 27625
rect 7006 27616 7012 27628
rect 7064 27616 7070 27668
rect 10962 27616 10968 27668
rect 11020 27616 11026 27668
rect 11146 27665 11152 27668
rect 11136 27659 11152 27665
rect 11136 27625 11148 27659
rect 11136 27619 11152 27625
rect 11146 27616 11152 27619
rect 11204 27616 11210 27668
rect 19521 27659 19579 27665
rect 19521 27625 19533 27659
rect 19567 27656 19579 27659
rect 19886 27656 19892 27668
rect 19567 27628 19892 27656
rect 19567 27625 19579 27628
rect 19521 27619 19579 27625
rect 19886 27616 19892 27628
rect 19944 27616 19950 27668
rect 20898 27616 20904 27668
rect 20956 27656 20962 27668
rect 22109 27659 22167 27665
rect 22109 27656 22121 27659
rect 20956 27628 22121 27656
rect 20956 27616 20962 27628
rect 22109 27625 22121 27628
rect 22155 27625 22167 27659
rect 22109 27619 22167 27625
rect 22738 27616 22744 27668
rect 22796 27656 22802 27668
rect 22925 27659 22983 27665
rect 22925 27656 22937 27659
rect 22796 27628 22937 27656
rect 22796 27616 22802 27628
rect 22925 27625 22937 27628
rect 22971 27625 22983 27659
rect 22925 27619 22983 27625
rect 26602 27616 26608 27668
rect 26660 27616 26666 27668
rect 4908 27560 5028 27588
rect 3234 27520 3240 27532
rect 2746 27492 3240 27520
rect 2746 27452 2774 27492
rect 3234 27480 3240 27492
rect 3292 27520 3298 27532
rect 3421 27523 3479 27529
rect 3421 27520 3433 27523
rect 3292 27492 3433 27520
rect 3292 27480 3298 27492
rect 3421 27489 3433 27492
rect 3467 27520 3479 27523
rect 3878 27520 3884 27532
rect 3467 27492 3884 27520
rect 3467 27489 3479 27492
rect 3421 27483 3479 27489
rect 3878 27480 3884 27492
rect 3936 27480 3942 27532
rect 3970 27480 3976 27532
rect 4028 27480 4034 27532
rect 5000 27520 5028 27560
rect 5810 27548 5816 27600
rect 5868 27548 5874 27600
rect 9674 27588 9680 27600
rect 9232 27560 9680 27588
rect 5000 27492 6132 27520
rect 2148 27424 2774 27452
rect 2148 27393 2176 27424
rect 3142 27412 3148 27464
rect 3200 27412 3206 27464
rect 3896 27452 3924 27480
rect 5902 27452 5908 27464
rect 3896 27424 5908 27452
rect 5902 27412 5908 27424
rect 5960 27452 5966 27464
rect 6104 27461 6132 27492
rect 7374 27480 7380 27532
rect 7432 27520 7438 27532
rect 9232 27529 9260 27560
rect 9674 27548 9680 27560
rect 9732 27548 9738 27600
rect 10980 27588 11008 27616
rect 9968 27560 11008 27588
rect 9968 27529 9996 27560
rect 13630 27548 13636 27600
rect 13688 27548 13694 27600
rect 20806 27588 20812 27600
rect 18432 27560 20812 27588
rect 9217 27523 9275 27529
rect 7432 27492 8892 27520
rect 7432 27480 7438 27492
rect 5997 27455 6055 27461
rect 5997 27452 6009 27455
rect 5960 27424 6009 27452
rect 5960 27412 5966 27424
rect 5997 27421 6009 27424
rect 6043 27421 6055 27455
rect 5997 27415 6055 27421
rect 6089 27455 6147 27461
rect 6089 27421 6101 27455
rect 6135 27421 6147 27455
rect 6089 27415 6147 27421
rect 6638 27412 6644 27464
rect 6696 27412 6702 27464
rect 8864 27452 8892 27492
rect 9217 27489 9229 27523
rect 9263 27489 9275 27523
rect 9953 27523 10011 27529
rect 9953 27520 9965 27523
rect 9217 27483 9275 27489
rect 9324 27492 9965 27520
rect 9324 27452 9352 27492
rect 9953 27489 9965 27492
rect 9999 27489 10011 27523
rect 11698 27520 11704 27532
rect 9953 27483 10011 27489
rect 10060 27492 11704 27520
rect 8864 27424 9352 27452
rect 10060 27438 10088 27492
rect 11698 27480 11704 27492
rect 11756 27480 11762 27532
rect 15470 27480 15476 27532
rect 15528 27480 15534 27532
rect 14648 27464 14700 27470
rect 10870 27412 10876 27464
rect 10928 27412 10934 27464
rect 13725 27455 13783 27461
rect 13725 27421 13737 27455
rect 13771 27452 13783 27455
rect 13814 27452 13820 27464
rect 13771 27424 13820 27452
rect 13771 27421 13783 27424
rect 13725 27415 13783 27421
rect 13814 27412 13820 27424
rect 13872 27412 13878 27464
rect 14090 27412 14096 27464
rect 14148 27452 14154 27464
rect 14553 27455 14611 27461
rect 14553 27452 14565 27455
rect 14148 27424 14565 27452
rect 14148 27412 14154 27424
rect 14553 27421 14565 27424
rect 14599 27421 14611 27455
rect 14553 27415 14611 27421
rect 18233 27455 18291 27461
rect 18233 27421 18245 27455
rect 18279 27452 18291 27455
rect 18432 27452 18460 27560
rect 20806 27548 20812 27560
rect 20864 27548 20870 27600
rect 23474 27548 23480 27600
rect 23532 27588 23538 27600
rect 23569 27591 23627 27597
rect 23569 27588 23581 27591
rect 23532 27560 23581 27588
rect 23532 27548 23538 27560
rect 23569 27557 23581 27560
rect 23615 27557 23627 27591
rect 23569 27551 23627 27557
rect 23658 27548 23664 27600
rect 23716 27588 23722 27600
rect 28994 27588 29000 27600
rect 23716 27560 29000 27588
rect 23716 27548 23722 27560
rect 28994 27548 29000 27560
rect 29052 27548 29058 27600
rect 18874 27480 18880 27532
rect 18932 27480 18938 27532
rect 21082 27520 21088 27532
rect 19168 27492 21088 27520
rect 18279 27424 18460 27452
rect 18509 27455 18567 27461
rect 18279 27421 18291 27424
rect 18233 27415 18291 27421
rect 18509 27421 18521 27455
rect 18555 27452 18567 27455
rect 19168 27452 19196 27492
rect 21082 27480 21088 27492
rect 21140 27480 21146 27532
rect 22370 27480 22376 27532
rect 22428 27480 22434 27532
rect 25777 27523 25835 27529
rect 25777 27489 25789 27523
rect 25823 27520 25835 27523
rect 25866 27520 25872 27532
rect 25823 27492 25872 27520
rect 25823 27489 25835 27492
rect 25777 27483 25835 27489
rect 25866 27480 25872 27492
rect 25924 27480 25930 27532
rect 26050 27480 26056 27532
rect 26108 27480 26114 27532
rect 28166 27480 28172 27532
rect 28224 27480 28230 27532
rect 18555 27424 19196 27452
rect 19613 27455 19671 27461
rect 18555 27421 18567 27424
rect 18509 27415 18567 27421
rect 19613 27421 19625 27455
rect 19659 27452 19671 27455
rect 23017 27455 23075 27461
rect 19659 27424 20668 27452
rect 19659 27421 19671 27424
rect 19613 27415 19671 27421
rect 2133 27387 2191 27393
rect 2133 27353 2145 27387
rect 2179 27353 2191 27387
rect 2133 27347 2191 27353
rect 2424 27356 3556 27384
rect 2314 27276 2320 27328
rect 2372 27325 2378 27328
rect 2372 27319 2391 27325
rect 2379 27316 2391 27319
rect 2424 27316 2452 27356
rect 2379 27288 2452 27316
rect 2501 27319 2559 27325
rect 2379 27285 2391 27288
rect 2372 27279 2391 27285
rect 2501 27285 2513 27319
rect 2547 27316 2559 27319
rect 3418 27316 3424 27328
rect 2547 27288 3424 27316
rect 2547 27285 2559 27288
rect 2501 27279 2559 27285
rect 2372 27276 2378 27279
rect 3418 27276 3424 27288
rect 3476 27276 3482 27328
rect 3528 27316 3556 27356
rect 3602 27344 3608 27396
rect 3660 27384 3666 27396
rect 4218 27387 4276 27393
rect 4218 27384 4230 27387
rect 3660 27356 4230 27384
rect 3660 27344 3666 27356
rect 4218 27353 4230 27356
rect 4264 27353 4276 27387
rect 4218 27347 4276 27353
rect 5813 27387 5871 27393
rect 5813 27353 5825 27387
rect 5859 27353 5871 27387
rect 5813 27347 5871 27353
rect 5353 27319 5411 27325
rect 5353 27316 5365 27319
rect 3528 27288 5365 27316
rect 5353 27285 5365 27288
rect 5399 27316 5411 27319
rect 5828 27316 5856 27347
rect 7650 27344 7656 27396
rect 7708 27344 7714 27396
rect 11790 27344 11796 27396
rect 11848 27344 11854 27396
rect 14108 27384 14136 27412
rect 14648 27406 14700 27412
rect 12452 27356 14136 27384
rect 5399 27288 5856 27316
rect 8389 27319 8447 27325
rect 5399 27285 5411 27288
rect 5353 27279 5411 27285
rect 8389 27285 8401 27319
rect 8435 27316 8447 27319
rect 8754 27316 8760 27328
rect 8435 27288 8760 27316
rect 8435 27285 8447 27288
rect 8389 27279 8447 27285
rect 8754 27276 8760 27288
rect 8812 27316 8818 27328
rect 9306 27316 9312 27328
rect 8812 27288 9312 27316
rect 8812 27276 8818 27288
rect 9306 27276 9312 27288
rect 9364 27276 9370 27328
rect 11054 27276 11060 27328
rect 11112 27316 11118 27328
rect 12452 27316 12480 27356
rect 11112 27288 12480 27316
rect 12621 27319 12679 27325
rect 11112 27276 11118 27288
rect 12621 27285 12633 27319
rect 12667 27316 12679 27319
rect 12710 27316 12716 27328
rect 12667 27288 12716 27316
rect 12667 27285 12679 27288
rect 12621 27279 12679 27285
rect 12710 27276 12716 27288
rect 12768 27276 12774 27328
rect 20640 27325 20668 27424
rect 23017 27421 23029 27455
rect 23063 27452 23075 27455
rect 23566 27452 23572 27464
rect 23063 27424 23572 27452
rect 23063 27421 23075 27424
rect 23017 27415 23075 27421
rect 23566 27412 23572 27424
rect 23624 27412 23630 27464
rect 23661 27455 23719 27461
rect 23661 27421 23673 27455
rect 23707 27421 23719 27455
rect 23661 27415 23719 27421
rect 25685 27455 25743 27461
rect 25685 27421 25697 27455
rect 25731 27452 25743 27455
rect 26418 27452 26424 27464
rect 25731 27424 26424 27452
rect 25731 27421 25743 27424
rect 25685 27415 25743 27421
rect 21358 27344 21364 27396
rect 21416 27344 21422 27396
rect 22922 27344 22928 27396
rect 22980 27384 22986 27396
rect 23676 27384 23704 27415
rect 26418 27412 26424 27424
rect 26476 27412 26482 27464
rect 26513 27455 26571 27461
rect 26513 27421 26525 27455
rect 26559 27452 26571 27455
rect 26602 27452 26608 27464
rect 26559 27424 26608 27452
rect 26559 27421 26571 27424
rect 26513 27415 26571 27421
rect 26602 27412 26608 27424
rect 26660 27412 26666 27464
rect 27614 27412 27620 27464
rect 27672 27412 27678 27464
rect 27890 27412 27896 27464
rect 27948 27412 27954 27464
rect 28721 27455 28779 27461
rect 28721 27421 28733 27455
rect 28767 27452 28779 27455
rect 28902 27452 28908 27464
rect 28767 27424 28908 27452
rect 28767 27421 28779 27424
rect 28721 27415 28779 27421
rect 26142 27384 26148 27396
rect 22980 27356 26148 27384
rect 22980 27344 22986 27356
rect 26142 27344 26148 27356
rect 26200 27344 26206 27396
rect 26436 27384 26464 27412
rect 28736 27384 28764 27415
rect 28902 27412 28908 27424
rect 28960 27412 28966 27464
rect 26436 27356 28764 27384
rect 20625 27319 20683 27325
rect 20625 27285 20637 27319
rect 20671 27316 20683 27319
rect 20714 27316 20720 27328
rect 20671 27288 20720 27316
rect 20671 27285 20683 27288
rect 20625 27279 20683 27285
rect 20714 27276 20720 27288
rect 20772 27276 20778 27328
rect 20806 27276 20812 27328
rect 20864 27316 20870 27328
rect 27614 27316 27620 27328
rect 20864 27288 27620 27316
rect 20864 27276 20870 27288
rect 27614 27276 27620 27288
rect 27672 27276 27678 27328
rect 28813 27319 28871 27325
rect 28813 27285 28825 27319
rect 28859 27316 28871 27319
rect 30190 27316 30196 27328
rect 28859 27288 30196 27316
rect 28859 27285 28871 27288
rect 28813 27279 28871 27285
rect 30190 27276 30196 27288
rect 30248 27276 30254 27328
rect 1104 27226 30976 27248
rect 1104 27174 8378 27226
rect 8430 27174 8442 27226
rect 8494 27174 8506 27226
rect 8558 27174 8570 27226
rect 8622 27174 8634 27226
rect 8686 27174 15806 27226
rect 15858 27174 15870 27226
rect 15922 27174 15934 27226
rect 15986 27174 15998 27226
rect 16050 27174 16062 27226
rect 16114 27174 23234 27226
rect 23286 27174 23298 27226
rect 23350 27174 23362 27226
rect 23414 27174 23426 27226
rect 23478 27174 23490 27226
rect 23542 27174 30662 27226
rect 30714 27174 30726 27226
rect 30778 27174 30790 27226
rect 30842 27174 30854 27226
rect 30906 27174 30918 27226
rect 30970 27174 30976 27226
rect 1104 27152 30976 27174
rect 3326 27072 3332 27124
rect 3384 27112 3390 27124
rect 5810 27112 5816 27124
rect 3384 27084 5816 27112
rect 3384 27072 3390 27084
rect 5810 27072 5816 27084
rect 5868 27072 5874 27124
rect 6638 27072 6644 27124
rect 6696 27112 6702 27124
rect 7377 27115 7435 27121
rect 7377 27112 7389 27115
rect 6696 27084 7389 27112
rect 6696 27072 6702 27084
rect 7377 27081 7389 27084
rect 7423 27081 7435 27115
rect 7377 27075 7435 27081
rect 19429 27115 19487 27121
rect 19429 27081 19441 27115
rect 19475 27112 19487 27115
rect 23658 27112 23664 27124
rect 19475 27084 23664 27112
rect 19475 27081 19487 27084
rect 19429 27075 19487 27081
rect 23658 27072 23664 27084
rect 23716 27072 23722 27124
rect 3136 27047 3194 27053
rect 3136 27013 3148 27047
rect 3182 27044 3194 27047
rect 5169 27047 5227 27053
rect 5169 27044 5181 27047
rect 3182 27016 5181 27044
rect 3182 27013 3194 27016
rect 3136 27007 3194 27013
rect 5169 27013 5181 27016
rect 5215 27013 5227 27047
rect 5169 27007 5227 27013
rect 11698 27004 11704 27056
rect 11756 27044 11762 27056
rect 11756 27016 12848 27044
rect 11756 27004 11762 27016
rect 2866 26936 2872 26988
rect 2924 26936 2930 26988
rect 3418 26936 3424 26988
rect 3476 26976 3482 26988
rect 4801 26979 4859 26985
rect 4801 26976 4813 26979
rect 3476 26948 4813 26976
rect 3476 26936 3482 26948
rect 4801 26945 4813 26948
rect 4847 26945 4859 26979
rect 4801 26939 4859 26945
rect 4982 26936 4988 26988
rect 5040 26936 5046 26988
rect 6825 26979 6883 26985
rect 6825 26945 6837 26979
rect 6871 26976 6883 26979
rect 7469 26979 7527 26985
rect 7469 26976 7481 26979
rect 6871 26948 7481 26976
rect 6871 26945 6883 26948
rect 6825 26939 6883 26945
rect 7469 26945 7481 26948
rect 7515 26976 7527 26979
rect 8294 26976 8300 26988
rect 7515 26948 8300 26976
rect 7515 26945 7527 26948
rect 7469 26939 7527 26945
rect 8294 26936 8300 26948
rect 8352 26936 8358 26988
rect 11882 26936 11888 26988
rect 11940 26936 11946 26988
rect 12820 26976 12848 27016
rect 13354 27004 13360 27056
rect 13412 27004 13418 27056
rect 14642 27044 14648 27056
rect 13464 27016 14648 27044
rect 13464 26976 13492 27016
rect 14642 27004 14648 27016
rect 14700 27004 14706 27056
rect 23566 27004 23572 27056
rect 23624 27044 23630 27056
rect 23624 27016 23704 27044
rect 23624 27004 23630 27016
rect 12820 26962 13492 26976
rect 12820 26948 13478 26962
rect 14090 26936 14096 26988
rect 14148 26936 14154 26988
rect 16045 26979 16103 26985
rect 16045 26945 16057 26979
rect 16091 26976 16103 26979
rect 16206 26976 16212 26988
rect 16091 26948 16212 26976
rect 16091 26945 16103 26948
rect 16045 26939 16103 26945
rect 16206 26936 16212 26948
rect 16264 26936 16270 26988
rect 18316 26979 18374 26985
rect 18316 26945 18328 26979
rect 18362 26976 18374 26979
rect 18598 26976 18604 26988
rect 18362 26948 18604 26976
rect 18362 26945 18374 26948
rect 18316 26939 18374 26945
rect 18598 26936 18604 26948
rect 18656 26976 18662 26988
rect 20070 26976 20076 26988
rect 18656 26948 20076 26976
rect 18656 26936 18662 26948
rect 20070 26936 20076 26948
rect 20128 26936 20134 26988
rect 23676 26985 23704 27016
rect 29178 27004 29184 27056
rect 29236 27004 29242 27056
rect 29914 27004 29920 27056
rect 29972 27004 29978 27056
rect 24946 26985 24952 26988
rect 23661 26979 23719 26985
rect 23661 26945 23673 26979
rect 23707 26945 23719 26979
rect 23661 26939 23719 26945
rect 24940 26939 24952 26985
rect 24946 26936 24952 26939
rect 25004 26936 25010 26988
rect 30190 26936 30196 26988
rect 30248 26936 30254 26988
rect 4709 26911 4767 26917
rect 4709 26908 4721 26911
rect 4264 26880 4721 26908
rect 4264 26852 4292 26880
rect 4709 26877 4721 26880
rect 4755 26877 4767 26911
rect 4709 26871 4767 26877
rect 11790 26868 11796 26920
rect 11848 26868 11854 26920
rect 16301 26911 16359 26917
rect 16301 26877 16313 26911
rect 16347 26908 16359 26911
rect 16574 26908 16580 26920
rect 16347 26880 16580 26908
rect 16347 26877 16359 26880
rect 16301 26871 16359 26877
rect 16574 26868 16580 26880
rect 16632 26868 16638 26920
rect 18046 26868 18052 26920
rect 18104 26868 18110 26920
rect 23106 26868 23112 26920
rect 23164 26908 23170 26920
rect 23569 26911 23627 26917
rect 23569 26908 23581 26911
rect 23164 26880 23581 26908
rect 23164 26868 23170 26880
rect 23569 26877 23581 26880
rect 23615 26877 23627 26911
rect 23569 26871 23627 26877
rect 24578 26868 24584 26920
rect 24636 26908 24642 26920
rect 24673 26911 24731 26917
rect 24673 26908 24685 26911
rect 24636 26880 24685 26908
rect 24636 26868 24642 26880
rect 24673 26877 24685 26880
rect 24719 26877 24731 26911
rect 24673 26871 24731 26877
rect 4246 26800 4252 26852
rect 4304 26800 4310 26852
rect 25866 26800 25872 26852
rect 25924 26840 25930 26852
rect 26053 26843 26111 26849
rect 26053 26840 26065 26843
rect 25924 26812 26065 26840
rect 25924 26800 25930 26812
rect 26053 26809 26065 26812
rect 26099 26809 26111 26843
rect 26053 26803 26111 26809
rect 6730 26732 6736 26784
rect 6788 26732 6794 26784
rect 12253 26775 12311 26781
rect 12253 26741 12265 26775
rect 12299 26772 12311 26775
rect 12894 26772 12900 26784
rect 12299 26744 12900 26772
rect 12299 26741 12311 26744
rect 12253 26735 12311 26741
rect 12894 26732 12900 26744
rect 12952 26732 12958 26784
rect 14921 26775 14979 26781
rect 14921 26741 14933 26775
rect 14967 26772 14979 26775
rect 15010 26772 15016 26784
rect 14967 26744 15016 26772
rect 14967 26741 14979 26744
rect 14921 26735 14979 26741
rect 15010 26732 15016 26744
rect 15068 26732 15074 26784
rect 24029 26775 24087 26781
rect 24029 26741 24041 26775
rect 24075 26772 24087 26775
rect 25958 26772 25964 26784
rect 24075 26744 25964 26772
rect 24075 26741 24087 26744
rect 24029 26735 24087 26741
rect 25958 26732 25964 26744
rect 26016 26732 26022 26784
rect 26142 26732 26148 26784
rect 26200 26772 26206 26784
rect 28445 26775 28503 26781
rect 28445 26772 28457 26775
rect 26200 26744 28457 26772
rect 26200 26732 26206 26744
rect 28445 26741 28457 26744
rect 28491 26772 28503 26775
rect 29454 26772 29460 26784
rect 28491 26744 29460 26772
rect 28491 26741 28503 26744
rect 28445 26735 28503 26741
rect 29454 26732 29460 26744
rect 29512 26732 29518 26784
rect 1104 26682 30820 26704
rect 1104 26630 4664 26682
rect 4716 26630 4728 26682
rect 4780 26630 4792 26682
rect 4844 26630 4856 26682
rect 4908 26630 4920 26682
rect 4972 26630 12092 26682
rect 12144 26630 12156 26682
rect 12208 26630 12220 26682
rect 12272 26630 12284 26682
rect 12336 26630 12348 26682
rect 12400 26630 19520 26682
rect 19572 26630 19584 26682
rect 19636 26630 19648 26682
rect 19700 26630 19712 26682
rect 19764 26630 19776 26682
rect 19828 26630 26948 26682
rect 27000 26630 27012 26682
rect 27064 26630 27076 26682
rect 27128 26630 27140 26682
rect 27192 26630 27204 26682
rect 27256 26630 30820 26682
rect 1104 26608 30820 26630
rect 3421 26571 3479 26577
rect 3421 26537 3433 26571
rect 3467 26568 3479 26571
rect 3602 26568 3608 26580
rect 3467 26540 3608 26568
rect 3467 26537 3479 26540
rect 3421 26531 3479 26537
rect 3602 26528 3608 26540
rect 3660 26528 3666 26580
rect 3878 26528 3884 26580
rect 3936 26568 3942 26580
rect 3936 26540 4568 26568
rect 3936 26528 3942 26540
rect 3326 26460 3332 26512
rect 3384 26460 3390 26512
rect 2314 26392 2320 26444
rect 2372 26432 2378 26444
rect 4540 26432 4568 26540
rect 11790 26528 11796 26580
rect 11848 26568 11854 26580
rect 12158 26568 12164 26580
rect 11848 26540 12164 26568
rect 11848 26528 11854 26540
rect 12158 26528 12164 26540
rect 12216 26568 12222 26580
rect 12529 26571 12587 26577
rect 12529 26568 12541 26571
rect 12216 26540 12541 26568
rect 12216 26528 12222 26540
rect 12529 26537 12541 26540
rect 12575 26537 12587 26571
rect 12529 26531 12587 26537
rect 16206 26528 16212 26580
rect 16264 26568 16270 26580
rect 16301 26571 16359 26577
rect 16301 26568 16313 26571
rect 16264 26540 16313 26568
rect 16264 26528 16270 26540
rect 16301 26537 16313 26540
rect 16347 26537 16359 26571
rect 16301 26531 16359 26537
rect 24857 26571 24915 26577
rect 24857 26537 24869 26571
rect 24903 26568 24915 26571
rect 24946 26568 24952 26580
rect 24903 26540 24952 26568
rect 24903 26537 24915 26540
rect 24857 26531 24915 26537
rect 24946 26528 24952 26540
rect 25004 26528 25010 26580
rect 26050 26528 26056 26580
rect 26108 26528 26114 26580
rect 26142 26528 26148 26580
rect 26200 26568 26206 26580
rect 26513 26571 26571 26577
rect 26513 26568 26525 26571
rect 26200 26540 26525 26568
rect 26200 26528 26206 26540
rect 26513 26537 26525 26540
rect 26559 26537 26571 26571
rect 26513 26531 26571 26537
rect 7374 26500 7380 26512
rect 6472 26472 7380 26500
rect 6472 26441 6500 26472
rect 7374 26460 7380 26472
rect 7432 26460 7438 26512
rect 8297 26503 8355 26509
rect 8297 26469 8309 26503
rect 8343 26500 8355 26503
rect 8343 26472 11192 26500
rect 8343 26469 8355 26472
rect 8297 26463 8355 26469
rect 4617 26435 4675 26441
rect 4617 26432 4629 26435
rect 2372 26404 4384 26432
rect 4540 26404 4629 26432
rect 2372 26392 2378 26404
rect 3418 26324 3424 26376
rect 3476 26324 3482 26376
rect 3786 26324 3792 26376
rect 3844 26364 3850 26376
rect 3844 26336 4200 26364
rect 3844 26324 3850 26336
rect 3050 26256 3056 26308
rect 3108 26296 3114 26308
rect 3145 26299 3203 26305
rect 3145 26296 3157 26299
rect 3108 26268 3157 26296
rect 3108 26256 3114 26268
rect 3145 26265 3157 26268
rect 3191 26296 3203 26299
rect 3970 26296 3976 26308
rect 3191 26268 3976 26296
rect 3191 26265 3203 26268
rect 3145 26259 3203 26265
rect 3970 26256 3976 26268
rect 4028 26256 4034 26308
rect 4065 26299 4123 26305
rect 4065 26265 4077 26299
rect 4111 26265 4123 26299
rect 4172 26296 4200 26336
rect 4246 26324 4252 26376
rect 4304 26324 4310 26376
rect 4356 26373 4384 26404
rect 4617 26401 4629 26404
rect 4663 26401 4675 26435
rect 4617 26395 4675 26401
rect 6457 26435 6515 26441
rect 6457 26401 6469 26435
rect 6503 26401 6515 26435
rect 6457 26395 6515 26401
rect 8018 26392 8024 26444
rect 8076 26392 8082 26444
rect 9401 26435 9459 26441
rect 9401 26401 9413 26435
rect 9447 26401 9459 26435
rect 9401 26395 9459 26401
rect 6920 26376 6972 26382
rect 4341 26367 4399 26373
rect 4341 26333 4353 26367
rect 4387 26333 4399 26367
rect 4341 26327 4399 26333
rect 7929 26367 7987 26373
rect 7929 26333 7941 26367
rect 7975 26364 7987 26367
rect 8294 26364 8300 26376
rect 7975 26336 8300 26364
rect 7975 26333 7987 26336
rect 7929 26327 7987 26333
rect 8294 26324 8300 26336
rect 8352 26324 8358 26376
rect 9306 26324 9312 26376
rect 9364 26324 9370 26376
rect 9416 26364 9444 26395
rect 9674 26392 9680 26444
rect 9732 26392 9738 26444
rect 11164 26432 11192 26472
rect 15028 26472 15884 26500
rect 15028 26444 15056 26472
rect 11164 26404 11284 26432
rect 10226 26364 10232 26376
rect 9416 26336 10232 26364
rect 10226 26324 10232 26336
rect 10284 26324 10290 26376
rect 11146 26324 11152 26376
rect 11204 26324 11210 26376
rect 11256 26364 11284 26404
rect 14550 26392 14556 26444
rect 14608 26392 14614 26444
rect 15010 26392 15016 26444
rect 15068 26392 15074 26444
rect 15194 26392 15200 26444
rect 15252 26432 15258 26444
rect 15856 26441 15884 26472
rect 23106 26460 23112 26512
rect 23164 26500 23170 26512
rect 23201 26503 23259 26509
rect 23201 26500 23213 26503
rect 23164 26472 23213 26500
rect 23164 26460 23170 26472
rect 23201 26469 23213 26472
rect 23247 26469 23259 26503
rect 25866 26500 25872 26512
rect 23201 26463 23259 26469
rect 25332 26472 25872 26500
rect 15657 26435 15715 26441
rect 15657 26432 15669 26435
rect 15252 26404 15669 26432
rect 15252 26392 15258 26404
rect 15657 26401 15669 26404
rect 15703 26401 15715 26435
rect 15657 26395 15715 26401
rect 15841 26435 15899 26441
rect 15841 26401 15853 26435
rect 15887 26401 15899 26435
rect 20806 26432 20812 26444
rect 15841 26395 15899 26401
rect 20272 26404 20812 26432
rect 12986 26364 12992 26376
rect 11256 26336 12992 26364
rect 12986 26324 12992 26336
rect 13044 26324 13050 26376
rect 14918 26324 14924 26376
rect 14976 26324 14982 26376
rect 15672 26336 15976 26364
rect 6920 26318 6972 26324
rect 15672 26308 15700 26336
rect 4433 26299 4491 26305
rect 4433 26296 4445 26299
rect 4172 26268 4445 26296
rect 4065 26259 4123 26265
rect 4433 26265 4445 26268
rect 4479 26265 4491 26299
rect 4433 26259 4491 26265
rect 4080 26228 4108 26259
rect 7282 26256 7288 26308
rect 7340 26256 7346 26308
rect 11416 26299 11474 26305
rect 11416 26265 11428 26299
rect 11462 26296 11474 26299
rect 11698 26296 11704 26308
rect 11462 26268 11704 26296
rect 11462 26265 11474 26268
rect 11416 26259 11474 26265
rect 11698 26256 11704 26268
rect 11756 26256 11762 26308
rect 15654 26256 15660 26308
rect 15712 26256 15718 26308
rect 15948 26305 15976 26336
rect 18782 26324 18788 26376
rect 18840 26324 18846 26376
rect 20272 26373 20300 26404
rect 20806 26392 20812 26404
rect 20864 26392 20870 26444
rect 25332 26441 25360 26472
rect 25866 26460 25872 26472
rect 25924 26460 25930 26512
rect 25317 26435 25375 26441
rect 25317 26401 25329 26435
rect 25363 26401 25375 26435
rect 25317 26395 25375 26401
rect 25406 26392 25412 26444
rect 25464 26392 25470 26444
rect 25958 26392 25964 26444
rect 26016 26432 26022 26444
rect 26145 26435 26203 26441
rect 26145 26432 26157 26435
rect 26016 26404 26157 26432
rect 26016 26392 26022 26404
rect 26145 26401 26157 26404
rect 26191 26401 26203 26435
rect 26145 26395 26203 26401
rect 27614 26392 27620 26444
rect 27672 26432 27678 26444
rect 27672 26404 28396 26432
rect 27672 26392 27678 26404
rect 20257 26367 20315 26373
rect 20257 26333 20269 26367
rect 20303 26333 20315 26367
rect 20257 26327 20315 26333
rect 20441 26367 20499 26373
rect 20441 26333 20453 26367
rect 20487 26364 20499 26367
rect 21082 26364 21088 26376
rect 20487 26336 21088 26364
rect 20487 26333 20499 26336
rect 20441 26327 20499 26333
rect 21082 26324 21088 26336
rect 21140 26324 21146 26376
rect 21818 26324 21824 26376
rect 21876 26324 21882 26376
rect 26326 26324 26332 26376
rect 26384 26324 26390 26376
rect 27890 26324 27896 26376
rect 27948 26364 27954 26376
rect 28368 26373 28396 26404
rect 28169 26367 28227 26373
rect 28169 26364 28181 26367
rect 27948 26336 28181 26364
rect 27948 26324 27954 26336
rect 28169 26333 28181 26336
rect 28215 26333 28227 26367
rect 28169 26327 28227 26333
rect 28353 26367 28411 26373
rect 28353 26333 28365 26367
rect 28399 26333 28411 26367
rect 28353 26327 28411 26333
rect 29914 26324 29920 26376
rect 29972 26324 29978 26376
rect 15933 26299 15991 26305
rect 15933 26265 15945 26299
rect 15979 26296 15991 26299
rect 22088 26299 22146 26305
rect 15979 26268 16033 26296
rect 18340 26268 18828 26296
rect 15979 26265 15991 26268
rect 15933 26259 15991 26265
rect 4154 26228 4160 26240
rect 4080 26200 4160 26228
rect 4154 26188 4160 26200
rect 4212 26188 4218 26240
rect 15948 26228 15976 26259
rect 18340 26228 18368 26268
rect 15948 26200 18368 26228
rect 18414 26188 18420 26240
rect 18472 26228 18478 26240
rect 18693 26231 18751 26237
rect 18693 26228 18705 26231
rect 18472 26200 18705 26228
rect 18472 26188 18478 26200
rect 18693 26197 18705 26200
rect 18739 26197 18751 26231
rect 18800 26228 18828 26268
rect 19352 26268 19564 26296
rect 19352 26228 19380 26268
rect 18800 26200 19380 26228
rect 18693 26191 18751 26197
rect 19426 26188 19432 26240
rect 19484 26188 19490 26240
rect 19536 26228 19564 26268
rect 22088 26265 22100 26299
rect 22134 26296 22146 26299
rect 22278 26296 22284 26308
rect 22134 26268 22284 26296
rect 22134 26265 22146 26268
rect 22088 26259 22146 26265
rect 22278 26256 22284 26268
rect 22336 26256 22342 26308
rect 25225 26299 25283 26305
rect 25225 26296 25237 26299
rect 22388 26268 25237 26296
rect 22002 26228 22008 26240
rect 19536 26200 22008 26228
rect 22002 26188 22008 26200
rect 22060 26188 22066 26240
rect 22186 26188 22192 26240
rect 22244 26228 22250 26240
rect 22388 26228 22416 26268
rect 25225 26265 25237 26268
rect 25271 26296 25283 26299
rect 25498 26296 25504 26308
rect 25271 26268 25504 26296
rect 25271 26265 25283 26268
rect 25225 26259 25283 26265
rect 25498 26256 25504 26268
rect 25556 26256 25562 26308
rect 26050 26256 26056 26308
rect 26108 26256 26114 26308
rect 26602 26256 26608 26308
rect 26660 26296 26666 26308
rect 29932 26296 29960 26324
rect 26660 26268 29960 26296
rect 26660 26256 26666 26268
rect 22244 26200 22416 26228
rect 22244 26188 22250 26200
rect 29178 26188 29184 26240
rect 29236 26188 29242 26240
rect 29822 26188 29828 26240
rect 29880 26188 29886 26240
rect 1104 26138 30976 26160
rect 1104 26086 8378 26138
rect 8430 26086 8442 26138
rect 8494 26086 8506 26138
rect 8558 26086 8570 26138
rect 8622 26086 8634 26138
rect 8686 26086 15806 26138
rect 15858 26086 15870 26138
rect 15922 26086 15934 26138
rect 15986 26086 15998 26138
rect 16050 26086 16062 26138
rect 16114 26086 23234 26138
rect 23286 26086 23298 26138
rect 23350 26086 23362 26138
rect 23414 26086 23426 26138
rect 23478 26086 23490 26138
rect 23542 26086 30662 26138
rect 30714 26086 30726 26138
rect 30778 26086 30790 26138
rect 30842 26086 30854 26138
rect 30906 26086 30918 26138
rect 30970 26086 30976 26138
rect 1104 26064 30976 26086
rect 2866 25984 2872 26036
rect 2924 25984 2930 26036
rect 8294 25984 8300 26036
rect 8352 25984 8358 26036
rect 10226 25984 10232 26036
rect 10284 25984 10290 26036
rect 11698 25984 11704 26036
rect 11756 25984 11762 26036
rect 12158 25984 12164 26036
rect 12216 25984 12222 26036
rect 20993 26027 21051 26033
rect 20993 26024 21005 26027
rect 18708 25996 21005 26024
rect 6730 25916 6736 25968
rect 6788 25956 6794 25968
rect 6825 25959 6883 25965
rect 6825 25956 6837 25959
rect 6788 25928 6837 25956
rect 6788 25916 6794 25928
rect 6825 25925 6837 25928
rect 6871 25925 6883 25959
rect 6825 25919 6883 25925
rect 7282 25916 7288 25968
rect 7340 25916 7346 25968
rect 12894 25916 12900 25968
rect 12952 25916 12958 25968
rect 18708 25965 18736 25996
rect 20993 25993 21005 25996
rect 21039 25993 21051 26027
rect 20993 25987 21051 25993
rect 22278 25984 22284 26036
rect 22336 25984 22342 26036
rect 22741 26027 22799 26033
rect 22741 25993 22753 26027
rect 22787 26024 22799 26027
rect 23106 26024 23112 26036
rect 22787 25996 23112 26024
rect 22787 25993 22799 25996
rect 22741 25987 22799 25993
rect 23106 25984 23112 25996
rect 23164 25984 23170 26036
rect 29914 25984 29920 26036
rect 29972 25984 29978 26036
rect 18693 25959 18751 25965
rect 18693 25925 18705 25959
rect 18739 25925 18751 25959
rect 18693 25919 18751 25925
rect 19426 25916 19432 25968
rect 19484 25916 19490 25968
rect 29178 25916 29184 25968
rect 29236 25916 29242 25968
rect 4338 25848 4344 25900
rect 4396 25848 4402 25900
rect 9116 25891 9174 25897
rect 9116 25857 9128 25891
rect 9162 25888 9174 25891
rect 9490 25888 9496 25900
rect 9162 25860 9496 25888
rect 9162 25857 9174 25860
rect 9116 25851 9174 25857
rect 9490 25848 9496 25860
rect 9548 25848 9554 25900
rect 11698 25848 11704 25900
rect 11756 25888 11762 25900
rect 12069 25891 12127 25897
rect 12069 25888 12081 25891
rect 11756 25860 12081 25888
rect 11756 25848 11762 25860
rect 12069 25857 12081 25860
rect 12115 25857 12127 25891
rect 12069 25851 12127 25857
rect 13173 25891 13231 25897
rect 13173 25857 13185 25891
rect 13219 25888 13231 25891
rect 14550 25888 14556 25900
rect 13219 25860 14556 25888
rect 13219 25857 13231 25860
rect 13173 25851 13231 25857
rect 14550 25848 14556 25860
rect 14608 25848 14614 25900
rect 18414 25848 18420 25900
rect 18472 25848 18478 25900
rect 20901 25891 20959 25897
rect 20901 25888 20913 25891
rect 20456 25860 20913 25888
rect 20456 25832 20484 25860
rect 20901 25857 20913 25860
rect 20947 25857 20959 25891
rect 20901 25851 20959 25857
rect 22002 25848 22008 25900
rect 22060 25888 22066 25900
rect 22649 25891 22707 25897
rect 22649 25888 22661 25891
rect 22060 25860 22661 25888
rect 22060 25848 22066 25860
rect 22649 25857 22661 25860
rect 22695 25888 22707 25891
rect 24670 25888 24676 25900
rect 22695 25860 24676 25888
rect 22695 25857 22707 25860
rect 22649 25851 22707 25857
rect 24670 25848 24676 25860
rect 24728 25848 24734 25900
rect 24854 25897 24860 25900
rect 24848 25851 24860 25897
rect 24854 25848 24860 25851
rect 24912 25848 24918 25900
rect 6546 25780 6552 25832
rect 6604 25780 6610 25832
rect 8849 25823 8907 25829
rect 8849 25789 8861 25823
rect 8895 25789 8907 25823
rect 8849 25783 8907 25789
rect 8864 25684 8892 25783
rect 11974 25780 11980 25832
rect 12032 25820 12038 25832
rect 12253 25823 12311 25829
rect 12253 25820 12265 25823
rect 12032 25792 12265 25820
rect 12032 25780 12038 25792
rect 12253 25789 12265 25792
rect 12299 25789 12311 25823
rect 12253 25783 12311 25789
rect 12986 25780 12992 25832
rect 13044 25780 13050 25832
rect 20438 25780 20444 25832
rect 20496 25780 20502 25832
rect 22833 25823 22891 25829
rect 22833 25789 22845 25823
rect 22879 25789 22891 25823
rect 22833 25783 22891 25789
rect 15102 25752 15108 25764
rect 13096 25724 15108 25752
rect 9122 25684 9128 25696
rect 8864 25656 9128 25684
rect 9122 25644 9128 25656
rect 9180 25644 9186 25696
rect 13096 25693 13124 25724
rect 15102 25712 15108 25724
rect 15160 25712 15166 25764
rect 22646 25712 22652 25764
rect 22704 25752 22710 25764
rect 22848 25752 22876 25783
rect 24578 25780 24584 25832
rect 24636 25780 24642 25832
rect 27982 25780 27988 25832
rect 28040 25820 28046 25832
rect 28169 25823 28227 25829
rect 28169 25820 28181 25823
rect 28040 25792 28181 25820
rect 28040 25780 28046 25792
rect 28169 25789 28181 25792
rect 28215 25789 28227 25823
rect 28169 25783 28227 25789
rect 28445 25823 28503 25829
rect 28445 25789 28457 25823
rect 28491 25820 28503 25823
rect 29822 25820 29828 25832
rect 28491 25792 29828 25820
rect 28491 25789 28503 25792
rect 28445 25783 28503 25789
rect 29822 25780 29828 25792
rect 29880 25780 29886 25832
rect 22704 25724 22876 25752
rect 22704 25712 22710 25724
rect 13081 25687 13139 25693
rect 13081 25653 13093 25687
rect 13127 25653 13139 25687
rect 13081 25647 13139 25653
rect 13170 25644 13176 25696
rect 13228 25684 13234 25696
rect 13357 25687 13415 25693
rect 13357 25684 13369 25687
rect 13228 25656 13369 25684
rect 13228 25644 13234 25656
rect 13357 25653 13369 25656
rect 13403 25653 13415 25687
rect 13357 25647 13415 25653
rect 25958 25644 25964 25696
rect 26016 25644 26022 25696
rect 1104 25594 30820 25616
rect 1104 25542 4664 25594
rect 4716 25542 4728 25594
rect 4780 25542 4792 25594
rect 4844 25542 4856 25594
rect 4908 25542 4920 25594
rect 4972 25542 12092 25594
rect 12144 25542 12156 25594
rect 12208 25542 12220 25594
rect 12272 25542 12284 25594
rect 12336 25542 12348 25594
rect 12400 25542 19520 25594
rect 19572 25542 19584 25594
rect 19636 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 26948 25594
rect 27000 25542 27012 25594
rect 27064 25542 27076 25594
rect 27128 25542 27140 25594
rect 27192 25542 27204 25594
rect 27256 25542 30820 25594
rect 1104 25520 30820 25542
rect 4157 25483 4215 25489
rect 4157 25449 4169 25483
rect 4203 25480 4215 25483
rect 4982 25480 4988 25492
rect 4203 25452 4988 25480
rect 4203 25449 4215 25452
rect 4157 25443 4215 25449
rect 4982 25440 4988 25452
rect 5040 25440 5046 25492
rect 8018 25440 8024 25492
rect 8076 25480 8082 25492
rect 8113 25483 8171 25489
rect 8113 25480 8125 25483
rect 8076 25452 8125 25480
rect 8076 25440 8082 25452
rect 8113 25449 8125 25452
rect 8159 25449 8171 25483
rect 8113 25443 8171 25449
rect 9490 25440 9496 25492
rect 9548 25440 9554 25492
rect 24765 25483 24823 25489
rect 24765 25449 24777 25483
rect 24811 25480 24823 25483
rect 24854 25480 24860 25492
rect 24811 25452 24860 25480
rect 24811 25449 24823 25452
rect 24765 25443 24823 25449
rect 24854 25440 24860 25452
rect 24912 25440 24918 25492
rect 27982 25440 27988 25492
rect 28040 25440 28046 25492
rect 11146 25412 11152 25424
rect 7760 25384 11152 25412
rect 2961 25279 3019 25285
rect 2961 25245 2973 25279
rect 3007 25245 3019 25279
rect 2961 25239 3019 25245
rect 2976 25208 3004 25239
rect 3142 25236 3148 25288
rect 3200 25236 3206 25288
rect 3234 25236 3240 25288
rect 3292 25236 3298 25288
rect 3973 25279 4031 25285
rect 3973 25245 3985 25279
rect 4019 25276 4031 25279
rect 4062 25276 4068 25288
rect 4019 25248 4068 25276
rect 4019 25245 4031 25248
rect 3973 25239 4031 25245
rect 4062 25236 4068 25248
rect 4120 25236 4126 25288
rect 4154 25236 4160 25288
rect 4212 25236 4218 25288
rect 6733 25279 6791 25285
rect 6733 25245 6745 25279
rect 6779 25276 6791 25279
rect 6822 25276 6828 25288
rect 6779 25248 6828 25276
rect 6779 25245 6791 25248
rect 6733 25239 6791 25245
rect 6822 25236 6828 25248
rect 6880 25276 6886 25288
rect 7760 25276 7788 25384
rect 11146 25372 11152 25384
rect 11204 25372 11210 25424
rect 19981 25415 20039 25421
rect 19981 25381 19993 25415
rect 20027 25412 20039 25415
rect 26326 25412 26332 25424
rect 20027 25384 26332 25412
rect 20027 25381 20039 25384
rect 19981 25375 20039 25381
rect 26326 25372 26332 25384
rect 26384 25372 26390 25424
rect 10137 25347 10195 25353
rect 10137 25313 10149 25347
rect 10183 25344 10195 25347
rect 11790 25344 11796 25356
rect 10183 25316 11796 25344
rect 10183 25313 10195 25316
rect 10137 25307 10195 25313
rect 11790 25304 11796 25316
rect 11848 25344 11854 25356
rect 11974 25344 11980 25356
rect 11848 25316 11980 25344
rect 11848 25304 11854 25316
rect 11974 25304 11980 25316
rect 12032 25304 12038 25356
rect 19518 25304 19524 25356
rect 19576 25304 19582 25356
rect 22646 25304 22652 25356
rect 22704 25344 22710 25356
rect 25317 25347 25375 25353
rect 25317 25344 25329 25347
rect 22704 25316 25329 25344
rect 22704 25304 22710 25316
rect 25317 25313 25329 25316
rect 25363 25344 25375 25347
rect 25406 25344 25412 25356
rect 25363 25316 25412 25344
rect 25363 25313 25375 25316
rect 25317 25307 25375 25313
rect 25406 25304 25412 25316
rect 25464 25304 25470 25356
rect 25958 25304 25964 25356
rect 26016 25344 26022 25356
rect 26053 25347 26111 25353
rect 26053 25344 26065 25347
rect 26016 25316 26065 25344
rect 26016 25304 26022 25316
rect 26053 25313 26065 25316
rect 26099 25313 26111 25347
rect 26053 25307 26111 25313
rect 26418 25304 26424 25356
rect 26476 25344 26482 25356
rect 26513 25347 26571 25353
rect 26513 25344 26525 25347
rect 26476 25316 26525 25344
rect 26476 25304 26482 25316
rect 26513 25313 26525 25316
rect 26559 25313 26571 25347
rect 26513 25307 26571 25313
rect 30101 25347 30159 25353
rect 30101 25313 30113 25347
rect 30147 25344 30159 25347
rect 31018 25344 31024 25356
rect 30147 25316 31024 25344
rect 30147 25313 30159 25316
rect 30101 25307 30159 25313
rect 31018 25304 31024 25316
rect 31076 25304 31082 25356
rect 6880 25248 7788 25276
rect 9953 25279 10011 25285
rect 6880 25236 6886 25248
rect 9953 25245 9965 25279
rect 9999 25276 10011 25279
rect 10226 25276 10232 25288
rect 9999 25248 10232 25276
rect 9999 25245 10011 25248
rect 9953 25239 10011 25245
rect 10226 25236 10232 25248
rect 10284 25236 10290 25288
rect 18782 25236 18788 25288
rect 18840 25276 18846 25288
rect 19613 25279 19671 25285
rect 19613 25276 19625 25279
rect 18840 25248 19625 25276
rect 18840 25236 18846 25248
rect 19613 25245 19625 25248
rect 19659 25245 19671 25279
rect 19613 25239 19671 25245
rect 22738 25236 22744 25288
rect 22796 25236 22802 25288
rect 22922 25236 22928 25288
rect 22980 25236 22986 25288
rect 25225 25279 25283 25285
rect 25225 25245 25237 25279
rect 25271 25276 25283 25279
rect 25976 25276 26004 25304
rect 25271 25248 26004 25276
rect 26145 25279 26203 25285
rect 25271 25245 25283 25248
rect 25225 25239 25283 25245
rect 26145 25245 26157 25279
rect 26191 25276 26203 25279
rect 26602 25276 26608 25288
rect 26191 25248 26608 25276
rect 26191 25245 26203 25248
rect 26145 25239 26203 25245
rect 26602 25236 26608 25248
rect 26660 25236 26666 25288
rect 27798 25236 27804 25288
rect 27856 25276 27862 25288
rect 27893 25279 27951 25285
rect 27893 25276 27905 25279
rect 27856 25248 27905 25276
rect 27856 25236 27862 25248
rect 27893 25245 27905 25248
rect 27939 25276 27951 25279
rect 28721 25279 28779 25285
rect 28721 25276 28733 25279
rect 27939 25248 28733 25276
rect 27939 25245 27951 25248
rect 27893 25239 27951 25245
rect 28721 25245 28733 25248
rect 28767 25276 28779 25279
rect 28902 25276 28908 25288
rect 28767 25248 28908 25276
rect 28767 25245 28779 25248
rect 28721 25239 28779 25245
rect 28902 25236 28908 25248
rect 28960 25236 28966 25288
rect 29822 25236 29828 25288
rect 29880 25236 29886 25288
rect 5258 25208 5264 25220
rect 2976 25180 5264 25208
rect 5258 25168 5264 25180
rect 5316 25168 5322 25220
rect 7006 25217 7012 25220
rect 7000 25171 7012 25217
rect 7006 25168 7012 25171
rect 7064 25168 7070 25220
rect 10778 25168 10784 25220
rect 10836 25168 10842 25220
rect 12529 25211 12587 25217
rect 12529 25177 12541 25211
rect 12575 25208 12587 25211
rect 14550 25208 14556 25220
rect 12575 25180 14556 25208
rect 12575 25177 12587 25180
rect 12529 25171 12587 25177
rect 14550 25168 14556 25180
rect 14608 25168 14614 25220
rect 2777 25143 2835 25149
rect 2777 25109 2789 25143
rect 2823 25140 2835 25143
rect 2866 25140 2872 25152
rect 2823 25112 2872 25140
rect 2823 25109 2835 25112
rect 2777 25103 2835 25109
rect 2866 25100 2872 25112
rect 2924 25100 2930 25152
rect 9858 25100 9864 25152
rect 9916 25100 9922 25152
rect 22925 25143 22983 25149
rect 22925 25109 22937 25143
rect 22971 25140 22983 25143
rect 23658 25140 23664 25152
rect 22971 25112 23664 25140
rect 22971 25109 22983 25112
rect 22925 25103 22983 25109
rect 23658 25100 23664 25112
rect 23716 25100 23722 25152
rect 25038 25100 25044 25152
rect 25096 25140 25102 25152
rect 25133 25143 25191 25149
rect 25133 25140 25145 25143
rect 25096 25112 25145 25140
rect 25096 25100 25102 25112
rect 25133 25109 25145 25112
rect 25179 25109 25191 25143
rect 25133 25103 25191 25109
rect 28442 25100 28448 25152
rect 28500 25140 28506 25152
rect 28629 25143 28687 25149
rect 28629 25140 28641 25143
rect 28500 25112 28641 25140
rect 28500 25100 28506 25112
rect 28629 25109 28641 25112
rect 28675 25109 28687 25143
rect 28629 25103 28687 25109
rect 1104 25050 30976 25072
rect 1104 24998 8378 25050
rect 8430 24998 8442 25050
rect 8494 24998 8506 25050
rect 8558 24998 8570 25050
rect 8622 24998 8634 25050
rect 8686 24998 15806 25050
rect 15858 24998 15870 25050
rect 15922 24998 15934 25050
rect 15986 24998 15998 25050
rect 16050 24998 16062 25050
rect 16114 24998 23234 25050
rect 23286 24998 23298 25050
rect 23350 24998 23362 25050
rect 23414 24998 23426 25050
rect 23478 24998 23490 25050
rect 23542 24998 30662 25050
rect 30714 24998 30726 25050
rect 30778 24998 30790 25050
rect 30842 24998 30854 25050
rect 30906 24998 30918 25050
rect 30970 24998 30976 25050
rect 1104 24976 30976 24998
rect 5905 24939 5963 24945
rect 5905 24905 5917 24939
rect 5951 24936 5963 24939
rect 6546 24936 6552 24948
rect 5951 24908 6552 24936
rect 5951 24905 5963 24908
rect 5905 24899 5963 24905
rect 6546 24896 6552 24908
rect 6604 24896 6610 24948
rect 6917 24939 6975 24945
rect 6917 24905 6929 24939
rect 6963 24936 6975 24939
rect 7006 24936 7012 24948
rect 6963 24908 7012 24936
rect 6963 24905 6975 24908
rect 6917 24899 6975 24905
rect 7006 24896 7012 24908
rect 7064 24896 7070 24948
rect 7377 24939 7435 24945
rect 7377 24905 7389 24939
rect 7423 24936 7435 24939
rect 8018 24936 8024 24948
rect 7423 24908 8024 24936
rect 7423 24905 7435 24908
rect 7377 24899 7435 24905
rect 8018 24896 8024 24908
rect 8076 24896 8082 24948
rect 8481 24939 8539 24945
rect 8481 24905 8493 24939
rect 8527 24936 8539 24939
rect 11146 24936 11152 24948
rect 8527 24908 11152 24936
rect 8527 24905 8539 24908
rect 8481 24899 8539 24905
rect 11146 24896 11152 24908
rect 11204 24896 11210 24948
rect 11698 24896 11704 24948
rect 11756 24936 11762 24948
rect 18230 24936 18236 24948
rect 11756 24908 18236 24936
rect 11756 24896 11762 24908
rect 18230 24896 18236 24908
rect 18288 24936 18294 24948
rect 22186 24936 22192 24948
rect 18288 24908 22192 24936
rect 18288 24896 18294 24908
rect 22186 24896 22192 24908
rect 22244 24896 22250 24948
rect 7285 24871 7343 24877
rect 7285 24837 7297 24871
rect 7331 24868 7343 24871
rect 15654 24868 15660 24880
rect 7331 24840 15660 24868
rect 7331 24837 7343 24840
rect 7285 24831 7343 24837
rect 15654 24828 15660 24840
rect 15712 24828 15718 24880
rect 28442 24828 28448 24880
rect 28500 24828 28506 24880
rect 2797 24803 2855 24809
rect 2797 24769 2809 24803
rect 2843 24800 2855 24803
rect 2958 24800 2964 24812
rect 2843 24772 2964 24800
rect 2843 24769 2855 24772
rect 2797 24763 2855 24769
rect 2958 24760 2964 24772
rect 3016 24760 3022 24812
rect 3050 24760 3056 24812
rect 3108 24760 3114 24812
rect 3510 24760 3516 24812
rect 3568 24760 3574 24812
rect 5997 24803 6055 24809
rect 5997 24769 6009 24803
rect 6043 24800 6055 24803
rect 6730 24800 6736 24812
rect 6043 24772 6736 24800
rect 6043 24769 6055 24772
rect 5997 24763 6055 24769
rect 6730 24760 6736 24772
rect 6788 24760 6794 24812
rect 8573 24803 8631 24809
rect 8573 24769 8585 24803
rect 8619 24800 8631 24803
rect 8754 24800 8760 24812
rect 8619 24772 8760 24800
rect 8619 24769 8631 24772
rect 8573 24763 8631 24769
rect 8754 24760 8760 24772
rect 8812 24760 8818 24812
rect 11977 24803 12035 24809
rect 11977 24769 11989 24803
rect 12023 24800 12035 24803
rect 12621 24803 12679 24809
rect 12023 24772 12434 24800
rect 12023 24769 12035 24772
rect 11977 24763 12035 24769
rect 7561 24735 7619 24741
rect 7561 24701 7573 24735
rect 7607 24732 7619 24735
rect 8665 24735 8723 24741
rect 8665 24732 8677 24735
rect 7607 24704 8677 24732
rect 7607 24701 7619 24704
rect 7561 24695 7619 24701
rect 8665 24701 8677 24704
rect 8711 24732 8723 24735
rect 9950 24732 9956 24744
rect 8711 24704 9956 24732
rect 8711 24701 8723 24704
rect 8665 24695 8723 24701
rect 9950 24692 9956 24704
rect 10008 24692 10014 24744
rect 12406 24732 12434 24772
rect 12621 24769 12633 24803
rect 12667 24800 12679 24803
rect 13998 24800 14004 24812
rect 12667 24772 14004 24800
rect 12667 24769 12679 24772
rect 12621 24763 12679 24769
rect 13998 24760 14004 24772
rect 14056 24760 14062 24812
rect 14090 24760 14096 24812
rect 14148 24760 14154 24812
rect 14642 24760 14648 24812
rect 14700 24760 14706 24812
rect 15930 24800 15936 24812
rect 14844 24772 15936 24800
rect 13354 24732 13360 24744
rect 12406 24704 13360 24732
rect 13354 24692 13360 24704
rect 13412 24692 13418 24744
rect 14016 24732 14044 24760
rect 14844 24732 14872 24772
rect 15930 24760 15936 24772
rect 15988 24760 15994 24812
rect 17580 24803 17638 24809
rect 17580 24769 17592 24803
rect 17626 24800 17638 24803
rect 17862 24800 17868 24812
rect 17626 24772 17868 24800
rect 17626 24769 17638 24772
rect 17580 24763 17638 24769
rect 17862 24760 17868 24772
rect 17920 24760 17926 24812
rect 19981 24803 20039 24809
rect 19981 24769 19993 24803
rect 20027 24800 20039 24803
rect 20438 24800 20444 24812
rect 20027 24772 20444 24800
rect 20027 24769 20039 24772
rect 19981 24763 20039 24769
rect 20438 24760 20444 24772
rect 20496 24760 20502 24812
rect 22097 24803 22155 24809
rect 22097 24800 22109 24803
rect 20548 24772 22109 24800
rect 14016 24704 14872 24732
rect 15010 24692 15016 24744
rect 15068 24692 15074 24744
rect 15102 24692 15108 24744
rect 15160 24732 15166 24744
rect 15565 24735 15623 24741
rect 15565 24732 15577 24735
rect 15160 24704 15577 24732
rect 15160 24692 15166 24704
rect 15565 24701 15577 24704
rect 15611 24701 15623 24735
rect 15565 24695 15623 24701
rect 16025 24735 16083 24741
rect 16025 24701 16037 24735
rect 16071 24732 16083 24735
rect 16298 24732 16304 24744
rect 16071 24704 16304 24732
rect 16071 24701 16083 24704
rect 16025 24695 16083 24701
rect 16298 24692 16304 24704
rect 16356 24692 16362 24744
rect 16574 24692 16580 24744
rect 16632 24732 16638 24744
rect 17313 24735 17371 24741
rect 17313 24732 17325 24735
rect 16632 24704 17325 24732
rect 16632 24692 16638 24704
rect 17313 24701 17325 24704
rect 17359 24701 17371 24735
rect 17313 24695 17371 24701
rect 11330 24624 11336 24676
rect 11388 24664 11394 24676
rect 12529 24667 12587 24673
rect 12529 24664 12541 24667
rect 11388 24636 12541 24664
rect 11388 24624 11394 24636
rect 12529 24633 12541 24636
rect 12575 24633 12587 24667
rect 12529 24627 12587 24633
rect 1673 24599 1731 24605
rect 1673 24565 1685 24599
rect 1719 24596 1731 24599
rect 3418 24596 3424 24608
rect 1719 24568 3424 24596
rect 1719 24565 1731 24568
rect 1673 24559 1731 24565
rect 3418 24556 3424 24568
rect 3476 24556 3482 24608
rect 4338 24556 4344 24608
rect 4396 24596 4402 24608
rect 4801 24599 4859 24605
rect 4801 24596 4813 24599
rect 4396 24568 4813 24596
rect 4396 24556 4402 24568
rect 4801 24565 4813 24568
rect 4847 24565 4859 24599
rect 4801 24559 4859 24565
rect 8110 24556 8116 24608
rect 8168 24556 8174 24608
rect 11606 24556 11612 24608
rect 11664 24596 11670 24608
rect 11885 24599 11943 24605
rect 11885 24596 11897 24599
rect 11664 24568 11897 24596
rect 11664 24556 11670 24568
rect 11885 24565 11897 24568
rect 11931 24565 11943 24599
rect 17328 24596 17356 24695
rect 19886 24692 19892 24744
rect 19944 24692 19950 24744
rect 18693 24667 18751 24673
rect 18693 24633 18705 24667
rect 18739 24664 18751 24667
rect 19334 24664 19340 24676
rect 18739 24636 19340 24664
rect 18739 24633 18751 24636
rect 18693 24627 18751 24633
rect 19334 24624 19340 24636
rect 19392 24664 19398 24676
rect 19518 24664 19524 24676
rect 19392 24636 19524 24664
rect 19392 24624 19398 24636
rect 19518 24624 19524 24636
rect 19576 24624 19582 24676
rect 20548 24664 20576 24772
rect 22097 24769 22109 24772
rect 22143 24769 22155 24803
rect 22097 24763 22155 24769
rect 22186 24760 22192 24812
rect 22244 24800 22250 24812
rect 23293 24803 23351 24809
rect 23293 24800 23305 24803
rect 22244 24772 23305 24800
rect 22244 24760 22250 24772
rect 23293 24769 23305 24772
rect 23339 24769 23351 24803
rect 23293 24763 23351 24769
rect 25685 24803 25743 24809
rect 25685 24769 25697 24803
rect 25731 24800 25743 24803
rect 27798 24800 27804 24812
rect 25731 24772 27804 24800
rect 25731 24769 25743 24772
rect 25685 24763 25743 24769
rect 27798 24760 27804 24772
rect 27856 24760 27862 24812
rect 29546 24760 29552 24812
rect 29604 24760 29610 24812
rect 21358 24692 21364 24744
rect 21416 24732 21422 24744
rect 21818 24732 21824 24744
rect 21416 24704 21824 24732
rect 21416 24692 21422 24704
rect 21818 24692 21824 24704
rect 21876 24732 21882 24744
rect 22281 24735 22339 24741
rect 22281 24732 22293 24735
rect 21876 24704 22293 24732
rect 21876 24692 21882 24704
rect 22281 24701 22293 24704
rect 22327 24732 22339 24735
rect 24578 24732 24584 24744
rect 22327 24704 24584 24732
rect 22327 24701 22339 24704
rect 22281 24695 22339 24701
rect 24578 24692 24584 24704
rect 24636 24692 24642 24744
rect 25774 24692 25780 24744
rect 25832 24692 25838 24744
rect 26050 24692 26056 24744
rect 26108 24692 26114 24744
rect 28169 24735 28227 24741
rect 28169 24701 28181 24735
rect 28215 24701 28227 24735
rect 28169 24695 28227 24701
rect 19628 24636 20576 24664
rect 18506 24596 18512 24608
rect 17328 24568 18512 24596
rect 11885 24559 11943 24565
rect 18506 24556 18512 24568
rect 18564 24596 18570 24608
rect 19628 24596 19656 24636
rect 18564 24568 19656 24596
rect 18564 24556 18570 24568
rect 20346 24556 20352 24608
rect 20404 24556 20410 24608
rect 23106 24556 23112 24608
rect 23164 24596 23170 24608
rect 24581 24599 24639 24605
rect 24581 24596 24593 24599
rect 23164 24568 24593 24596
rect 23164 24556 23170 24568
rect 24581 24565 24593 24568
rect 24627 24565 24639 24599
rect 28184 24596 28212 24695
rect 28902 24692 28908 24744
rect 28960 24732 28966 24744
rect 29917 24735 29975 24741
rect 29917 24732 29929 24735
rect 28960 24704 29929 24732
rect 28960 24692 28966 24704
rect 29917 24701 29929 24704
rect 29963 24701 29975 24735
rect 29917 24695 29975 24701
rect 28258 24596 28264 24608
rect 28184 24568 28264 24596
rect 24581 24559 24639 24565
rect 28258 24556 28264 24568
rect 28316 24556 28322 24608
rect 1104 24506 30820 24528
rect 1104 24454 4664 24506
rect 4716 24454 4728 24506
rect 4780 24454 4792 24506
rect 4844 24454 4856 24506
rect 4908 24454 4920 24506
rect 4972 24454 12092 24506
rect 12144 24454 12156 24506
rect 12208 24454 12220 24506
rect 12272 24454 12284 24506
rect 12336 24454 12348 24506
rect 12400 24454 19520 24506
rect 19572 24454 19584 24506
rect 19636 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 26948 24506
rect 27000 24454 27012 24506
rect 27064 24454 27076 24506
rect 27128 24454 27140 24506
rect 27192 24454 27204 24506
rect 27256 24454 30820 24506
rect 1104 24432 30820 24454
rect 2958 24352 2964 24404
rect 3016 24352 3022 24404
rect 3234 24352 3240 24404
rect 3292 24392 3298 24404
rect 3970 24392 3976 24404
rect 3292 24364 3976 24392
rect 3292 24352 3298 24364
rect 3970 24352 3976 24364
rect 4028 24392 4034 24404
rect 4157 24395 4215 24401
rect 4157 24392 4169 24395
rect 4028 24364 4169 24392
rect 4028 24352 4034 24364
rect 4157 24361 4169 24364
rect 4203 24361 4215 24395
rect 4157 24355 4215 24361
rect 15930 24352 15936 24404
rect 15988 24392 15994 24404
rect 16025 24395 16083 24401
rect 16025 24392 16037 24395
rect 15988 24364 16037 24392
rect 15988 24352 15994 24364
rect 16025 24361 16037 24364
rect 16071 24361 16083 24395
rect 16025 24355 16083 24361
rect 17862 24352 17868 24404
rect 17920 24352 17926 24404
rect 22738 24352 22744 24404
rect 22796 24352 22802 24404
rect 3142 24284 3148 24336
rect 3200 24324 3206 24336
rect 4341 24327 4399 24333
rect 3200 24296 3648 24324
rect 3200 24284 3206 24296
rect 2409 24259 2467 24265
rect 2409 24225 2421 24259
rect 2455 24256 2467 24259
rect 2455 24228 2774 24256
rect 2455 24225 2467 24228
rect 2409 24219 2467 24225
rect 2314 24148 2320 24200
rect 2372 24148 2378 24200
rect 2501 24191 2559 24197
rect 2501 24157 2513 24191
rect 2547 24157 2559 24191
rect 2746 24188 2774 24228
rect 3145 24191 3203 24197
rect 3145 24188 3157 24191
rect 2746 24160 3157 24188
rect 2501 24151 2559 24157
rect 3145 24157 3157 24160
rect 3191 24157 3203 24191
rect 3145 24151 3203 24157
rect 2516 24120 2544 24151
rect 3252 24120 3280 24296
rect 3418 24216 3424 24268
rect 3476 24216 3482 24268
rect 3620 24256 3648 24296
rect 4341 24293 4353 24327
rect 4387 24324 4399 24327
rect 5166 24324 5172 24336
rect 4387 24296 5172 24324
rect 4387 24293 4399 24296
rect 4341 24287 4399 24293
rect 5166 24284 5172 24296
rect 5224 24284 5230 24336
rect 4801 24259 4859 24265
rect 4801 24256 4813 24259
rect 3620 24228 4813 24256
rect 4801 24225 4813 24228
rect 4847 24225 4859 24259
rect 4801 24219 4859 24225
rect 7374 24216 7380 24268
rect 7432 24216 7438 24268
rect 11330 24216 11336 24268
rect 11388 24216 11394 24268
rect 11606 24216 11612 24268
rect 11664 24216 11670 24268
rect 13354 24216 13360 24268
rect 13412 24216 13418 24268
rect 18414 24216 18420 24268
rect 18472 24216 18478 24268
rect 19886 24216 19892 24268
rect 19944 24216 19950 24268
rect 19978 24216 19984 24268
rect 20036 24216 20042 24268
rect 21358 24216 21364 24268
rect 21416 24216 21422 24268
rect 25130 24216 25136 24268
rect 25188 24216 25194 24268
rect 25961 24259 26019 24265
rect 25961 24225 25973 24259
rect 26007 24256 26019 24259
rect 26142 24256 26148 24268
rect 26007 24228 26148 24256
rect 26007 24225 26019 24228
rect 25961 24219 26019 24225
rect 26142 24216 26148 24228
rect 26200 24216 26206 24268
rect 27614 24216 27620 24268
rect 27672 24256 27678 24268
rect 29181 24259 29239 24265
rect 27672 24228 28396 24256
rect 27672 24216 27678 24228
rect 3329 24191 3387 24197
rect 3329 24157 3341 24191
rect 3375 24157 3387 24191
rect 3329 24151 3387 24157
rect 2516 24092 3280 24120
rect 3344 24052 3372 24151
rect 3436 24120 3464 24216
rect 6920 24200 6972 24206
rect 4154 24148 4160 24200
rect 4212 24188 4218 24200
rect 4985 24191 5043 24197
rect 4985 24188 4997 24191
rect 4212 24160 4997 24188
rect 4212 24148 4218 24160
rect 4985 24157 4997 24160
rect 5031 24157 5043 24191
rect 4985 24151 5043 24157
rect 5077 24191 5135 24197
rect 5077 24157 5089 24191
rect 5123 24157 5135 24191
rect 5077 24151 5135 24157
rect 3973 24123 4031 24129
rect 3973 24120 3985 24123
rect 3436 24092 3985 24120
rect 3973 24089 3985 24092
rect 4019 24120 4031 24123
rect 5092 24120 5120 24151
rect 13446 24148 13452 24200
rect 13504 24188 13510 24200
rect 14277 24191 14335 24197
rect 14277 24188 14289 24191
rect 13504 24160 14289 24188
rect 13504 24148 13510 24160
rect 14277 24157 14289 24160
rect 14323 24157 14335 24191
rect 14277 24151 14335 24157
rect 18230 24148 18236 24200
rect 18288 24148 18294 24200
rect 18325 24191 18383 24197
rect 18325 24157 18337 24191
rect 18371 24188 18383 24191
rect 19334 24188 19340 24200
rect 18371 24160 19340 24188
rect 18371 24157 18383 24160
rect 18325 24151 18383 24157
rect 19334 24148 19340 24160
rect 19392 24148 19398 24200
rect 22922 24148 22928 24200
rect 22980 24188 22986 24200
rect 23385 24191 23443 24197
rect 23385 24188 23397 24191
rect 22980 24160 23397 24188
rect 22980 24148 22986 24160
rect 23385 24157 23397 24160
rect 23431 24157 23443 24191
rect 23385 24151 23443 24157
rect 24946 24148 24952 24200
rect 25004 24188 25010 24200
rect 26053 24191 26111 24197
rect 26053 24188 26065 24191
rect 25004 24160 26065 24188
rect 25004 24148 25010 24160
rect 26053 24157 26065 24160
rect 26099 24157 26111 24191
rect 26053 24151 26111 24157
rect 26326 24148 26332 24200
rect 26384 24148 26390 24200
rect 27890 24148 27896 24200
rect 27948 24188 27954 24200
rect 28166 24188 28172 24200
rect 27948 24160 28172 24188
rect 27948 24148 27954 24160
rect 28166 24148 28172 24160
rect 28224 24148 28230 24200
rect 28368 24197 28396 24228
rect 29181 24225 29193 24259
rect 29227 24256 29239 24259
rect 29546 24256 29552 24268
rect 29227 24228 29552 24256
rect 29227 24225 29239 24228
rect 29181 24219 29239 24225
rect 29546 24216 29552 24228
rect 29604 24216 29610 24268
rect 28353 24191 28411 24197
rect 28353 24157 28365 24191
rect 28399 24188 28411 24191
rect 28442 24188 28448 24200
rect 28399 24160 28448 24188
rect 28399 24157 28411 24160
rect 28353 24151 28411 24157
rect 28442 24148 28448 24160
rect 28500 24148 28506 24200
rect 6920 24142 6972 24148
rect 4019 24092 5120 24120
rect 6825 24123 6883 24129
rect 4019 24089 4031 24092
rect 3973 24083 4031 24089
rect 6825 24089 6837 24123
rect 6871 24089 6883 24123
rect 6825 24083 6883 24089
rect 4154 24052 4160 24064
rect 4212 24061 4218 24064
rect 4212 24055 4231 24061
rect 3344 24024 4160 24052
rect 4154 24012 4160 24024
rect 4219 24021 4231 24055
rect 6840 24052 6868 24083
rect 12618 24080 12624 24132
rect 12676 24080 12682 24132
rect 14090 24080 14096 24132
rect 14148 24120 14154 24132
rect 14553 24123 14611 24129
rect 14553 24120 14565 24123
rect 14148 24092 14565 24120
rect 14148 24080 14154 24092
rect 14553 24089 14565 24092
rect 14599 24089 14611 24123
rect 14553 24083 14611 24089
rect 15010 24080 15016 24132
rect 15068 24080 15074 24132
rect 21628 24123 21686 24129
rect 21628 24089 21640 24123
rect 21674 24120 21686 24123
rect 22002 24120 22008 24132
rect 21674 24092 22008 24120
rect 21674 24089 21686 24092
rect 21628 24083 21686 24089
rect 22002 24080 22008 24092
rect 22060 24080 22066 24132
rect 22738 24080 22744 24132
rect 22796 24120 22802 24132
rect 23201 24123 23259 24129
rect 23201 24120 23213 24123
rect 22796 24092 23213 24120
rect 22796 24080 22802 24092
rect 23201 24089 23213 24092
rect 23247 24089 23259 24123
rect 23201 24083 23259 24089
rect 24670 24080 24676 24132
rect 24728 24120 24734 24132
rect 28534 24120 28540 24132
rect 24728 24092 28540 24120
rect 24728 24080 24734 24092
rect 7098 24052 7104 24064
rect 6840 24024 7104 24052
rect 4212 24015 4231 24021
rect 4212 24012 4218 24015
rect 7098 24012 7104 24024
rect 7156 24012 7162 24064
rect 19426 24012 19432 24064
rect 19484 24012 19490 24064
rect 19797 24055 19855 24061
rect 19797 24021 19809 24055
rect 19843 24052 19855 24055
rect 20162 24052 20168 24064
rect 19843 24024 20168 24052
rect 19843 24021 19855 24024
rect 19797 24015 19855 24021
rect 20162 24012 20168 24024
rect 20220 24052 20226 24064
rect 22370 24052 22376 24064
rect 20220 24024 22376 24052
rect 20220 24012 20226 24024
rect 22370 24012 22376 24024
rect 22428 24012 22434 24064
rect 23566 24012 23572 24064
rect 23624 24012 23630 24064
rect 24581 24055 24639 24061
rect 24581 24021 24593 24055
rect 24627 24052 24639 24055
rect 24854 24052 24860 24064
rect 24627 24024 24860 24052
rect 24627 24021 24639 24024
rect 24581 24015 24639 24021
rect 24854 24012 24860 24024
rect 24912 24012 24918 24064
rect 24964 24061 24992 24092
rect 28534 24080 28540 24092
rect 28592 24080 28598 24132
rect 24949 24055 25007 24061
rect 24949 24021 24961 24055
rect 24995 24021 25007 24055
rect 24949 24015 25007 24021
rect 25041 24055 25099 24061
rect 25041 24021 25053 24055
rect 25087 24052 25099 24055
rect 25774 24052 25780 24064
rect 25087 24024 25780 24052
rect 25087 24021 25099 24024
rect 25041 24015 25099 24021
rect 25774 24012 25780 24024
rect 25832 24012 25838 24064
rect 26142 24012 26148 24064
rect 26200 24012 26206 24064
rect 1104 23962 30976 23984
rect 1104 23910 8378 23962
rect 8430 23910 8442 23962
rect 8494 23910 8506 23962
rect 8558 23910 8570 23962
rect 8622 23910 8634 23962
rect 8686 23910 15806 23962
rect 15858 23910 15870 23962
rect 15922 23910 15934 23962
rect 15986 23910 15998 23962
rect 16050 23910 16062 23962
rect 16114 23910 23234 23962
rect 23286 23910 23298 23962
rect 23350 23910 23362 23962
rect 23414 23910 23426 23962
rect 23478 23910 23490 23962
rect 23542 23910 30662 23962
rect 30714 23910 30726 23962
rect 30778 23910 30790 23962
rect 30842 23910 30854 23962
rect 30906 23910 30918 23962
rect 30970 23910 30976 23962
rect 1104 23888 30976 23910
rect 2746 23820 3004 23848
rect 2314 23740 2320 23792
rect 2372 23780 2378 23792
rect 2746 23780 2774 23820
rect 2866 23789 2872 23792
rect 2860 23780 2872 23789
rect 2372 23752 2774 23780
rect 2827 23752 2872 23780
rect 2372 23740 2378 23752
rect 2860 23743 2872 23752
rect 2866 23740 2872 23743
rect 2924 23740 2930 23792
rect 2976 23780 3004 23820
rect 3970 23808 3976 23860
rect 4028 23808 4034 23860
rect 5258 23808 5264 23860
rect 5316 23808 5322 23860
rect 13446 23808 13452 23860
rect 13504 23808 13510 23860
rect 14090 23808 14096 23860
rect 14148 23808 14154 23860
rect 16298 23808 16304 23860
rect 16356 23808 16362 23860
rect 19886 23808 19892 23860
rect 19944 23808 19950 23860
rect 22002 23808 22008 23860
rect 22060 23808 22066 23860
rect 22465 23851 22523 23857
rect 22465 23817 22477 23851
rect 22511 23848 22523 23851
rect 22738 23848 22744 23860
rect 22511 23820 22744 23848
rect 22511 23817 22523 23820
rect 22465 23811 22523 23817
rect 22738 23808 22744 23820
rect 22796 23808 22802 23860
rect 26053 23851 26111 23857
rect 26053 23817 26065 23851
rect 26099 23848 26111 23851
rect 26326 23848 26332 23860
rect 26099 23820 26332 23848
rect 26099 23817 26111 23820
rect 26053 23811 26111 23817
rect 26326 23808 26332 23820
rect 26384 23808 26390 23860
rect 28258 23808 28264 23860
rect 28316 23848 28322 23860
rect 28353 23851 28411 23857
rect 28353 23848 28365 23851
rect 28316 23820 28365 23848
rect 28316 23808 28322 23820
rect 28353 23817 28365 23820
rect 28399 23817 28411 23851
rect 28353 23811 28411 23817
rect 4062 23780 4068 23792
rect 2976 23752 4068 23780
rect 4062 23740 4068 23752
rect 4120 23780 4126 23792
rect 4120 23752 5120 23780
rect 4120 23740 4126 23752
rect 2593 23715 2651 23721
rect 2593 23681 2605 23715
rect 2639 23712 2651 23715
rect 2682 23712 2688 23724
rect 2639 23684 2688 23712
rect 2639 23681 2651 23684
rect 2593 23675 2651 23681
rect 2682 23672 2688 23684
rect 2740 23672 2746 23724
rect 4709 23715 4767 23721
rect 4709 23681 4721 23715
rect 4755 23712 4767 23715
rect 4982 23712 4988 23724
rect 4755 23684 4988 23712
rect 4755 23681 4767 23684
rect 4709 23675 4767 23681
rect 4982 23672 4988 23684
rect 5040 23672 5046 23724
rect 5092 23656 5120 23752
rect 6914 23740 6920 23792
rect 6972 23780 6978 23792
rect 7837 23783 7895 23789
rect 7837 23780 7849 23783
rect 6972 23752 7849 23780
rect 6972 23740 6978 23752
rect 7837 23749 7849 23752
rect 7883 23749 7895 23783
rect 7837 23743 7895 23749
rect 9585 23783 9643 23789
rect 9585 23749 9597 23783
rect 9631 23780 9643 23783
rect 10778 23780 10784 23792
rect 9631 23752 10784 23780
rect 9631 23749 9643 23752
rect 9585 23743 9643 23749
rect 10778 23740 10784 23752
rect 10836 23740 10842 23792
rect 11974 23740 11980 23792
rect 12032 23780 12038 23792
rect 12529 23783 12587 23789
rect 12032 23752 12480 23780
rect 12032 23740 12038 23752
rect 5166 23672 5172 23724
rect 5224 23672 5230 23724
rect 5353 23715 5411 23721
rect 5353 23681 5365 23715
rect 5399 23681 5411 23715
rect 5353 23675 5411 23681
rect 10137 23715 10195 23721
rect 10137 23681 10149 23715
rect 10183 23712 10195 23715
rect 10183 23684 10364 23712
rect 10183 23681 10195 23684
rect 10137 23675 10195 23681
rect 5074 23604 5080 23656
rect 5132 23644 5138 23656
rect 5368 23644 5396 23675
rect 5132 23616 5396 23644
rect 5132 23604 5138 23616
rect 9674 23604 9680 23656
rect 9732 23644 9738 23656
rect 10229 23647 10287 23653
rect 10229 23644 10241 23647
rect 9732 23616 10241 23644
rect 9732 23604 9738 23616
rect 10229 23613 10241 23616
rect 10275 23613 10287 23647
rect 10336 23644 10364 23684
rect 10410 23672 10416 23724
rect 10468 23672 10474 23724
rect 11054 23672 11060 23724
rect 11112 23712 11118 23724
rect 11793 23715 11851 23721
rect 11793 23712 11805 23715
rect 11112 23684 11805 23712
rect 11112 23672 11118 23684
rect 11793 23681 11805 23684
rect 11839 23681 11851 23715
rect 12452 23712 12480 23752
rect 12529 23749 12541 23783
rect 12575 23780 12587 23783
rect 12618 23780 12624 23792
rect 12575 23752 12624 23780
rect 12575 23749 12587 23752
rect 12529 23743 12587 23749
rect 12618 23740 12624 23752
rect 12676 23740 12682 23792
rect 14642 23780 14648 23792
rect 13096 23752 14648 23780
rect 13096 23712 13124 23752
rect 14642 23740 14648 23752
rect 14700 23740 14706 23792
rect 18776 23783 18834 23789
rect 18776 23749 18788 23783
rect 18822 23780 18834 23783
rect 19426 23780 19432 23792
rect 18822 23752 19432 23780
rect 18822 23749 18834 23752
rect 18776 23743 18834 23749
rect 19426 23740 19432 23752
rect 19484 23740 19490 23792
rect 23106 23740 23112 23792
rect 23164 23780 23170 23792
rect 23385 23783 23443 23789
rect 23385 23780 23397 23783
rect 23164 23752 23397 23780
rect 23164 23740 23170 23752
rect 23385 23749 23397 23752
rect 23431 23749 23443 23783
rect 23385 23743 23443 23749
rect 25133 23783 25191 23789
rect 25133 23749 25145 23783
rect 25179 23780 25191 23783
rect 28166 23780 28172 23792
rect 25179 23752 28172 23780
rect 25179 23749 25191 23752
rect 25133 23743 25191 23749
rect 28166 23740 28172 23752
rect 28224 23740 28230 23792
rect 12452 23698 13124 23712
rect 12466 23684 13124 23698
rect 13357 23715 13415 23721
rect 11793 23675 11851 23681
rect 13357 23681 13369 23715
rect 13403 23712 13415 23715
rect 13722 23712 13728 23724
rect 13403 23684 13728 23712
rect 13403 23681 13415 23684
rect 13357 23675 13415 23681
rect 11238 23644 11244 23656
rect 10336 23616 11244 23644
rect 10229 23607 10287 23613
rect 11238 23604 11244 23616
rect 11296 23604 11302 23656
rect 12986 23604 12992 23656
rect 13044 23644 13050 23656
rect 13372 23644 13400 23675
rect 13722 23672 13728 23684
rect 13780 23672 13786 23724
rect 13998 23672 14004 23724
rect 14056 23672 14062 23724
rect 15188 23715 15246 23721
rect 15188 23681 15200 23715
rect 15234 23712 15246 23715
rect 15470 23712 15476 23724
rect 15234 23684 15476 23712
rect 15234 23681 15246 23684
rect 15188 23675 15246 23681
rect 15470 23672 15476 23684
rect 15528 23672 15534 23724
rect 18506 23672 18512 23724
rect 18564 23672 18570 23724
rect 20714 23672 20720 23724
rect 20772 23712 20778 23724
rect 20993 23715 21051 23721
rect 20993 23712 21005 23715
rect 20772 23684 21005 23712
rect 20772 23672 20778 23684
rect 20993 23681 21005 23684
rect 21039 23681 21051 23715
rect 20993 23675 21051 23681
rect 22370 23672 22376 23724
rect 22428 23712 22434 23724
rect 25682 23712 25688 23724
rect 22428 23684 25688 23712
rect 22428 23672 22434 23684
rect 25682 23672 25688 23684
rect 25740 23672 25746 23724
rect 25958 23672 25964 23724
rect 26016 23712 26022 23724
rect 26237 23715 26295 23721
rect 26237 23712 26249 23715
rect 26016 23684 26249 23712
rect 26016 23672 26022 23684
rect 26237 23681 26249 23684
rect 26283 23681 26295 23715
rect 26237 23675 26295 23681
rect 26510 23672 26516 23724
rect 26568 23672 26574 23724
rect 28445 23715 28503 23721
rect 28445 23681 28457 23715
rect 28491 23712 28503 23715
rect 28902 23712 28908 23724
rect 28491 23684 28908 23712
rect 28491 23681 28503 23684
rect 28445 23675 28503 23681
rect 28902 23672 28908 23684
rect 28960 23672 28966 23724
rect 13044 23616 13400 23644
rect 13044 23604 13050 23616
rect 14918 23604 14924 23656
rect 14976 23604 14982 23656
rect 20898 23604 20904 23656
rect 20956 23604 20962 23656
rect 22646 23604 22652 23656
rect 22704 23604 22710 23656
rect 26418 23604 26424 23656
rect 26476 23604 26482 23656
rect 20346 23536 20352 23588
rect 20404 23576 20410 23588
rect 20404 23548 26280 23576
rect 20404 23536 20410 23548
rect 4522 23468 4528 23520
rect 4580 23468 4586 23520
rect 10134 23468 10140 23520
rect 10192 23468 10198 23520
rect 10597 23511 10655 23517
rect 10597 23477 10609 23511
rect 10643 23508 10655 23511
rect 11514 23508 11520 23520
rect 10643 23480 11520 23508
rect 10643 23477 10655 23480
rect 10597 23471 10655 23477
rect 11514 23468 11520 23480
rect 11572 23468 11578 23520
rect 18414 23468 18420 23520
rect 18472 23508 18478 23520
rect 19978 23508 19984 23520
rect 18472 23480 19984 23508
rect 18472 23468 18478 23480
rect 19978 23468 19984 23480
rect 20036 23468 20042 23520
rect 21361 23511 21419 23517
rect 21361 23477 21373 23511
rect 21407 23508 21419 23511
rect 23014 23508 23020 23520
rect 21407 23480 23020 23508
rect 21407 23477 21419 23480
rect 21361 23471 21419 23477
rect 23014 23468 23020 23480
rect 23072 23468 23078 23520
rect 26252 23517 26280 23548
rect 26237 23511 26295 23517
rect 26237 23477 26249 23511
rect 26283 23477 26295 23511
rect 26237 23471 26295 23477
rect 1104 23418 30820 23440
rect 1104 23366 4664 23418
rect 4716 23366 4728 23418
rect 4780 23366 4792 23418
rect 4844 23366 4856 23418
rect 4908 23366 4920 23418
rect 4972 23366 12092 23418
rect 12144 23366 12156 23418
rect 12208 23366 12220 23418
rect 12272 23366 12284 23418
rect 12336 23366 12348 23418
rect 12400 23366 19520 23418
rect 19572 23366 19584 23418
rect 19636 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 26948 23418
rect 27000 23366 27012 23418
rect 27064 23366 27076 23418
rect 27128 23366 27140 23418
rect 27192 23366 27204 23418
rect 27256 23366 30820 23418
rect 1104 23344 30820 23366
rect 4246 23264 4252 23316
rect 4304 23264 4310 23316
rect 4982 23264 4988 23316
rect 5040 23264 5046 23316
rect 6730 23264 6736 23316
rect 6788 23304 6794 23316
rect 7561 23307 7619 23313
rect 7561 23304 7573 23307
rect 6788 23276 7573 23304
rect 6788 23264 6794 23276
rect 7561 23273 7573 23276
rect 7607 23273 7619 23307
rect 7561 23267 7619 23273
rect 9677 23307 9735 23313
rect 9677 23273 9689 23307
rect 9723 23304 9735 23307
rect 10134 23304 10140 23316
rect 9723 23276 10140 23304
rect 9723 23273 9735 23276
rect 9677 23267 9735 23273
rect 3053 23239 3111 23245
rect 3053 23205 3065 23239
rect 3099 23236 3111 23239
rect 5166 23236 5172 23248
rect 3099 23208 5172 23236
rect 3099 23205 3111 23208
rect 3053 23199 3111 23205
rect 5166 23196 5172 23208
rect 5224 23196 5230 23248
rect 2314 23168 2320 23180
rect 1688 23140 2320 23168
rect 1688 23109 1716 23140
rect 2314 23128 2320 23140
rect 2372 23128 2378 23180
rect 1673 23103 1731 23109
rect 1673 23069 1685 23103
rect 1719 23069 1731 23103
rect 1673 23063 1731 23069
rect 1854 23060 1860 23112
rect 1912 23060 1918 23112
rect 2869 23103 2927 23109
rect 2869 23100 2881 23103
rect 2746 23072 2881 23100
rect 1765 23035 1823 23041
rect 1765 23001 1777 23035
rect 1811 23032 1823 23035
rect 2746 23032 2774 23072
rect 2869 23069 2881 23072
rect 2915 23069 2927 23103
rect 2869 23063 2927 23069
rect 3145 23103 3203 23109
rect 3145 23069 3157 23103
rect 3191 23100 3203 23103
rect 3694 23100 3700 23112
rect 3191 23072 3700 23100
rect 3191 23069 3203 23072
rect 3145 23063 3203 23069
rect 3694 23060 3700 23072
rect 3752 23060 3758 23112
rect 4341 23103 4399 23109
rect 4341 23069 4353 23103
rect 4387 23100 4399 23103
rect 4522 23100 4528 23112
rect 4387 23072 4528 23100
rect 4387 23069 4399 23072
rect 4341 23063 4399 23069
rect 4522 23060 4528 23072
rect 4580 23060 4586 23112
rect 5169 23103 5227 23109
rect 5169 23069 5181 23103
rect 5215 23069 5227 23103
rect 5169 23063 5227 23069
rect 1811 23004 2774 23032
rect 1811 23001 1823 23004
rect 1765 22995 1823 23001
rect 2314 22924 2320 22976
rect 2372 22964 2378 22976
rect 2685 22967 2743 22973
rect 2685 22964 2697 22967
rect 2372 22936 2697 22964
rect 2372 22924 2378 22936
rect 2685 22933 2697 22936
rect 2731 22933 2743 22967
rect 2685 22927 2743 22933
rect 4154 22924 4160 22976
rect 4212 22964 4218 22976
rect 5184 22964 5212 23063
rect 5810 23060 5816 23112
rect 5868 23060 5874 23112
rect 7576 23100 7604 23267
rect 10134 23264 10140 23276
rect 10192 23264 10198 23316
rect 11885 23307 11943 23313
rect 11885 23273 11897 23307
rect 11931 23304 11943 23307
rect 11974 23304 11980 23316
rect 11931 23276 11980 23304
rect 11931 23273 11943 23276
rect 11885 23267 11943 23273
rect 11974 23264 11980 23276
rect 12032 23264 12038 23316
rect 15470 23264 15476 23316
rect 15528 23264 15534 23316
rect 21082 23264 21088 23316
rect 21140 23264 21146 23316
rect 23661 23307 23719 23313
rect 23661 23273 23673 23307
rect 23707 23304 23719 23307
rect 24946 23304 24952 23316
rect 23707 23276 24952 23304
rect 23707 23273 23719 23276
rect 23661 23267 23719 23273
rect 24946 23264 24952 23276
rect 25004 23264 25010 23316
rect 25774 23264 25780 23316
rect 25832 23304 25838 23316
rect 25961 23307 26019 23313
rect 25961 23304 25973 23307
rect 25832 23276 25973 23304
rect 25832 23264 25838 23276
rect 25961 23273 25973 23276
rect 26007 23273 26019 23307
rect 25961 23267 26019 23273
rect 26421 23307 26479 23313
rect 26421 23273 26433 23307
rect 26467 23304 26479 23307
rect 26510 23304 26516 23316
rect 26467 23276 26516 23304
rect 26467 23273 26479 23276
rect 26421 23267 26479 23273
rect 26510 23264 26516 23276
rect 26568 23264 26574 23316
rect 11238 23196 11244 23248
rect 11296 23236 11302 23248
rect 12621 23239 12679 23245
rect 12621 23236 12633 23239
rect 11296 23208 12633 23236
rect 11296 23196 11302 23208
rect 12621 23205 12633 23208
rect 12667 23205 12679 23239
rect 12621 23199 12679 23205
rect 23106 23196 23112 23248
rect 23164 23196 23170 23248
rect 23566 23196 23572 23248
rect 23624 23196 23630 23248
rect 8754 23128 8760 23180
rect 8812 23168 8818 23180
rect 9217 23171 9275 23177
rect 9217 23168 9229 23171
rect 8812 23140 9229 23168
rect 8812 23128 8818 23140
rect 9217 23137 9229 23140
rect 9263 23137 9275 23171
rect 9217 23131 9275 23137
rect 13081 23171 13139 23177
rect 13081 23137 13093 23171
rect 13127 23168 13139 23171
rect 15654 23168 15660 23180
rect 13127 23140 15660 23168
rect 13127 23137 13139 23140
rect 13081 23131 13139 23137
rect 15654 23128 15660 23140
rect 15712 23128 15718 23180
rect 16117 23171 16175 23177
rect 16117 23137 16129 23171
rect 16163 23168 16175 23171
rect 16574 23168 16580 23180
rect 16163 23140 16580 23168
rect 16163 23137 16175 23140
rect 16117 23131 16175 23137
rect 16574 23128 16580 23140
rect 16632 23128 16638 23180
rect 19978 23128 19984 23180
rect 20036 23128 20042 23180
rect 23124 23168 23152 23196
rect 23584 23168 23612 23196
rect 22572 23140 23152 23168
rect 23400 23140 23612 23168
rect 9309 23103 9367 23109
rect 9309 23100 9321 23103
rect 7576 23072 9321 23100
rect 9309 23069 9321 23072
rect 9355 23069 9367 23103
rect 9309 23063 9367 23069
rect 10413 23103 10471 23109
rect 10413 23069 10425 23103
rect 10459 23100 10471 23103
rect 10778 23100 10784 23112
rect 10459 23072 10784 23100
rect 10459 23069 10471 23072
rect 10413 23063 10471 23069
rect 10778 23060 10784 23072
rect 10836 23060 10842 23112
rect 12989 23103 13047 23109
rect 12989 23069 13001 23103
rect 13035 23100 13047 23103
rect 13354 23100 13360 23112
rect 13035 23072 13360 23100
rect 13035 23069 13047 23072
rect 12989 23063 13047 23069
rect 13354 23060 13360 23072
rect 13412 23060 13418 23112
rect 15933 23103 15991 23109
rect 15933 23069 15945 23103
rect 15979 23100 15991 23103
rect 16298 23100 16304 23112
rect 15979 23072 16304 23100
rect 15979 23069 15991 23072
rect 15933 23063 15991 23069
rect 16298 23060 16304 23072
rect 16356 23060 16362 23112
rect 19889 23103 19947 23109
rect 19889 23069 19901 23103
rect 19935 23100 19947 23103
rect 20898 23100 20904 23112
rect 19935 23072 20904 23100
rect 19935 23069 19947 23072
rect 19889 23063 19947 23069
rect 20898 23060 20904 23072
rect 20956 23060 20962 23112
rect 22572 23109 22600 23140
rect 22557 23103 22615 23109
rect 22557 23069 22569 23103
rect 22603 23069 22615 23103
rect 22557 23063 22615 23069
rect 23014 23060 23020 23112
rect 23072 23060 23078 23112
rect 23106 23060 23112 23112
rect 23164 23060 23170 23112
rect 23400 23109 23428 23140
rect 24578 23128 24584 23180
rect 24636 23128 24642 23180
rect 25866 23128 25872 23180
rect 25924 23168 25930 23180
rect 26697 23171 26755 23177
rect 26697 23168 26709 23171
rect 25924 23140 26709 23168
rect 25924 23128 25930 23140
rect 26697 23137 26709 23140
rect 26743 23137 26755 23171
rect 26697 23131 26755 23137
rect 23385 23103 23443 23109
rect 23385 23069 23397 23103
rect 23431 23069 23443 23103
rect 23385 23063 23443 23069
rect 23523 23103 23581 23109
rect 23523 23069 23535 23103
rect 23569 23100 23581 23103
rect 23658 23100 23664 23112
rect 23569 23072 23664 23100
rect 23569 23069 23581 23072
rect 23523 23063 23581 23069
rect 23658 23060 23664 23072
rect 23716 23060 23722 23112
rect 24854 23109 24860 23112
rect 24848 23100 24860 23109
rect 24815 23072 24860 23100
rect 24848 23063 24860 23072
rect 24854 23060 24860 23063
rect 24912 23060 24918 23112
rect 26789 23103 26847 23109
rect 26789 23069 26801 23103
rect 26835 23069 26847 23103
rect 26789 23063 26847 23069
rect 6086 22992 6092 23044
rect 6144 22992 6150 23044
rect 7098 22992 7104 23044
rect 7156 22992 7162 23044
rect 21450 22992 21456 23044
rect 21508 23032 21514 23044
rect 23293 23035 23351 23041
rect 23293 23032 23305 23035
rect 21508 23004 23305 23032
rect 21508 22992 21514 23004
rect 23293 23001 23305 23004
rect 23339 23001 23351 23035
rect 26804 23032 26832 23063
rect 28534 23060 28540 23112
rect 28592 23060 28598 23112
rect 28902 23060 28908 23112
rect 28960 23100 28966 23112
rect 29181 23103 29239 23109
rect 29181 23100 29193 23103
rect 28960 23072 29193 23100
rect 28960 23060 28966 23072
rect 29181 23069 29193 23072
rect 29227 23069 29239 23103
rect 29181 23063 29239 23069
rect 28920 23032 28948 23060
rect 26804 23004 28948 23032
rect 23293 22995 23351 23001
rect 14734 22964 14740 22976
rect 4212 22936 14740 22964
rect 4212 22924 4218 22936
rect 14734 22924 14740 22936
rect 14792 22924 14798 22976
rect 15470 22924 15476 22976
rect 15528 22964 15534 22976
rect 15841 22967 15899 22973
rect 15841 22964 15853 22967
rect 15528 22936 15853 22964
rect 15528 22924 15534 22936
rect 15841 22933 15853 22936
rect 15887 22933 15899 22967
rect 15841 22927 15899 22933
rect 19426 22924 19432 22976
rect 19484 22924 19490 22976
rect 19797 22967 19855 22973
rect 19797 22933 19809 22967
rect 19843 22964 19855 22967
rect 20070 22964 20076 22976
rect 19843 22936 20076 22964
rect 19843 22933 19855 22936
rect 19797 22927 19855 22933
rect 20070 22924 20076 22936
rect 20128 22964 20134 22976
rect 21266 22964 21272 22976
rect 20128 22936 21272 22964
rect 20128 22924 20134 22936
rect 21266 22924 21272 22936
rect 21324 22964 21330 22976
rect 22370 22964 22376 22976
rect 21324 22936 22376 22964
rect 21324 22924 21330 22936
rect 22370 22924 22376 22936
rect 22428 22964 22434 22976
rect 25038 22964 25044 22976
rect 22428 22936 25044 22964
rect 22428 22924 22434 22936
rect 25038 22924 25044 22936
rect 25096 22924 25102 22976
rect 28350 22924 28356 22976
rect 28408 22964 28414 22976
rect 28445 22967 28503 22973
rect 28445 22964 28457 22967
rect 28408 22936 28457 22964
rect 28408 22924 28414 22936
rect 28445 22933 28457 22936
rect 28491 22933 28503 22967
rect 28445 22927 28503 22933
rect 28626 22924 28632 22976
rect 28684 22964 28690 22976
rect 29089 22967 29147 22973
rect 29089 22964 29101 22967
rect 28684 22936 29101 22964
rect 28684 22924 28690 22936
rect 29089 22933 29101 22936
rect 29135 22933 29147 22967
rect 29089 22927 29147 22933
rect 1104 22874 30976 22896
rect 1104 22822 8378 22874
rect 8430 22822 8442 22874
rect 8494 22822 8506 22874
rect 8558 22822 8570 22874
rect 8622 22822 8634 22874
rect 8686 22822 15806 22874
rect 15858 22822 15870 22874
rect 15922 22822 15934 22874
rect 15986 22822 15998 22874
rect 16050 22822 16062 22874
rect 16114 22822 23234 22874
rect 23286 22822 23298 22874
rect 23350 22822 23362 22874
rect 23414 22822 23426 22874
rect 23478 22822 23490 22874
rect 23542 22822 30662 22874
rect 30714 22822 30726 22874
rect 30778 22822 30790 22874
rect 30842 22822 30854 22874
rect 30906 22822 30918 22874
rect 30970 22822 30976 22874
rect 1104 22800 30976 22822
rect 2041 22763 2099 22769
rect 2041 22729 2053 22763
rect 2087 22760 2099 22763
rect 4062 22760 4068 22772
rect 2087 22732 4068 22760
rect 2087 22729 2099 22732
rect 2041 22723 2099 22729
rect 4062 22720 4068 22732
rect 4120 22720 4126 22772
rect 6086 22720 6092 22772
rect 6144 22760 6150 22772
rect 6641 22763 6699 22769
rect 6641 22760 6653 22763
rect 6144 22732 6653 22760
rect 6144 22720 6150 22732
rect 6641 22729 6653 22732
rect 6687 22729 6699 22763
rect 6641 22723 6699 22729
rect 8754 22720 8760 22772
rect 8812 22720 8818 22772
rect 15654 22720 15660 22772
rect 15712 22760 15718 22772
rect 15841 22763 15899 22769
rect 15841 22760 15853 22763
rect 15712 22732 15853 22760
rect 15712 22720 15718 22732
rect 15841 22729 15853 22732
rect 15887 22729 15899 22763
rect 20162 22760 20168 22772
rect 15841 22723 15899 22729
rect 17788 22732 20168 22760
rect 1854 22652 1860 22704
rect 1912 22692 1918 22704
rect 3326 22692 3332 22704
rect 1912 22664 3332 22692
rect 1912 22652 1918 22664
rect 1964 22633 1992 22664
rect 3326 22652 3332 22664
rect 3384 22692 3390 22704
rect 5445 22695 5503 22701
rect 5445 22692 5457 22695
rect 3384 22664 5457 22692
rect 3384 22652 3390 22664
rect 5445 22661 5457 22664
rect 5491 22661 5503 22695
rect 5445 22655 5503 22661
rect 7644 22695 7702 22701
rect 7644 22661 7656 22695
rect 7690 22692 7702 22695
rect 8110 22692 8116 22704
rect 7690 22664 8116 22692
rect 7690 22661 7702 22664
rect 7644 22655 7702 22661
rect 8110 22652 8116 22664
rect 8168 22652 8174 22704
rect 9766 22692 9772 22704
rect 8680 22664 9772 22692
rect 1949 22627 2007 22633
rect 1949 22593 1961 22627
rect 1995 22593 2007 22627
rect 1949 22587 2007 22593
rect 2222 22584 2228 22636
rect 2280 22584 2286 22636
rect 2958 22633 2964 22636
rect 2952 22587 2964 22633
rect 2958 22584 2964 22587
rect 3016 22584 3022 22636
rect 4246 22584 4252 22636
rect 4304 22624 4310 22636
rect 4525 22627 4583 22633
rect 4525 22624 4537 22627
rect 4304 22596 4537 22624
rect 4304 22584 4310 22596
rect 4525 22593 4537 22596
rect 4571 22624 4583 22627
rect 4571 22596 5120 22624
rect 4571 22593 4583 22596
rect 4525 22587 4583 22593
rect 2682 22516 2688 22568
rect 2740 22516 2746 22568
rect 4801 22559 4859 22565
rect 4801 22525 4813 22559
rect 4847 22556 4859 22559
rect 4982 22556 4988 22568
rect 4847 22528 4988 22556
rect 4847 22525 4859 22528
rect 4801 22519 4859 22525
rect 4982 22516 4988 22528
rect 5040 22516 5046 22568
rect 5092 22556 5120 22596
rect 5166 22584 5172 22636
rect 5224 22624 5230 22636
rect 5629 22627 5687 22633
rect 5629 22624 5641 22627
rect 5224 22596 5641 22624
rect 5224 22584 5230 22596
rect 5629 22593 5641 22596
rect 5675 22593 5687 22627
rect 5629 22587 5687 22593
rect 6730 22584 6736 22636
rect 6788 22584 6794 22636
rect 6822 22584 6828 22636
rect 6880 22624 6886 22636
rect 7377 22627 7435 22633
rect 7377 22624 7389 22627
rect 6880 22596 7389 22624
rect 6880 22584 6886 22596
rect 7377 22593 7389 22596
rect 7423 22624 7435 22627
rect 8680 22624 8708 22664
rect 9766 22652 9772 22664
rect 9824 22652 9830 22704
rect 11514 22652 11520 22704
rect 11572 22692 11578 22704
rect 12897 22695 12955 22701
rect 12897 22692 12909 22695
rect 11572 22664 12909 22692
rect 11572 22652 11578 22664
rect 12897 22661 12909 22664
rect 12943 22661 12955 22695
rect 12897 22655 12955 22661
rect 14734 22652 14740 22704
rect 14792 22652 14798 22704
rect 17788 22701 17816 22732
rect 20162 22720 20168 22732
rect 20220 22720 20226 22772
rect 20257 22763 20315 22769
rect 20257 22729 20269 22763
rect 20303 22760 20315 22763
rect 20898 22760 20904 22772
rect 20303 22732 20904 22760
rect 20303 22729 20315 22732
rect 20257 22723 20315 22729
rect 20898 22720 20904 22732
rect 20956 22720 20962 22772
rect 21450 22720 21456 22772
rect 21508 22720 21514 22772
rect 22370 22720 22376 22772
rect 22428 22720 22434 22772
rect 23106 22720 23112 22772
rect 23164 22760 23170 22772
rect 23201 22763 23259 22769
rect 23201 22760 23213 22763
rect 23164 22732 23213 22760
rect 23164 22720 23170 22732
rect 23201 22729 23213 22732
rect 23247 22729 23259 22763
rect 23201 22723 23259 22729
rect 25866 22720 25872 22772
rect 25924 22720 25930 22772
rect 28902 22720 28908 22772
rect 28960 22760 28966 22772
rect 30101 22763 30159 22769
rect 30101 22760 30113 22763
rect 28960 22732 30113 22760
rect 28960 22720 28966 22732
rect 30101 22729 30113 22732
rect 30147 22729 30159 22763
rect 30101 22723 30159 22729
rect 17773 22695 17831 22701
rect 17773 22661 17785 22695
rect 17819 22661 17831 22695
rect 17773 22655 17831 22661
rect 19144 22695 19202 22701
rect 19144 22661 19156 22695
rect 19190 22692 19202 22695
rect 19426 22692 19432 22704
rect 19190 22664 19432 22692
rect 19190 22661 19202 22664
rect 19144 22655 19202 22661
rect 19426 22652 19432 22664
rect 19484 22652 19490 22704
rect 22278 22652 22284 22704
rect 22336 22692 22342 22704
rect 23014 22692 23020 22704
rect 22336 22664 23020 22692
rect 22336 22652 22342 22664
rect 23014 22652 23020 22664
rect 23072 22692 23078 22704
rect 23569 22695 23627 22701
rect 23569 22692 23581 22695
rect 23072 22664 23581 22692
rect 23072 22652 23078 22664
rect 23569 22661 23581 22664
rect 23615 22661 23627 22695
rect 23569 22655 23627 22661
rect 28626 22652 28632 22704
rect 28684 22652 28690 22704
rect 29178 22652 29184 22704
rect 29236 22652 29242 22704
rect 7423 22596 8708 22624
rect 7423 22593 7435 22596
rect 7377 22587 7435 22593
rect 8754 22584 8760 22636
rect 8812 22624 8818 22636
rect 9401 22627 9459 22633
rect 9401 22624 9413 22627
rect 8812 22596 9413 22624
rect 8812 22584 8818 22596
rect 9401 22593 9413 22596
rect 9447 22593 9459 22627
rect 9401 22587 9459 22593
rect 11422 22584 11428 22636
rect 11480 22624 11486 22636
rect 12069 22627 12127 22633
rect 12069 22624 12081 22627
rect 11480 22596 12081 22624
rect 11480 22584 11486 22596
rect 12069 22593 12081 22596
rect 12115 22593 12127 22627
rect 12069 22587 12127 22593
rect 12253 22627 12311 22633
rect 12253 22593 12265 22627
rect 12299 22624 12311 22627
rect 12710 22624 12716 22636
rect 12299 22596 12716 22624
rect 12299 22593 12311 22596
rect 12253 22587 12311 22593
rect 12710 22584 12716 22596
rect 12768 22584 12774 22636
rect 13170 22584 13176 22636
rect 13228 22584 13234 22636
rect 15933 22627 15991 22633
rect 15933 22624 15945 22627
rect 13280 22596 15945 22624
rect 5258 22556 5264 22568
rect 5092 22528 5264 22556
rect 5258 22516 5264 22528
rect 5316 22516 5322 22568
rect 5813 22559 5871 22565
rect 5813 22525 5825 22559
rect 5859 22525 5871 22559
rect 5813 22519 5871 22525
rect 9493 22559 9551 22565
rect 9493 22525 9505 22559
rect 9539 22556 9551 22559
rect 9674 22556 9680 22568
rect 9539 22528 9680 22556
rect 9539 22525 9551 22528
rect 9493 22519 9551 22525
rect 3694 22448 3700 22500
rect 3752 22488 3758 22500
rect 5828 22488 5856 22519
rect 9674 22516 9680 22528
rect 9732 22516 9738 22568
rect 9769 22559 9827 22565
rect 9769 22525 9781 22559
rect 9815 22556 9827 22559
rect 10410 22556 10416 22568
rect 9815 22528 10416 22556
rect 9815 22525 9827 22528
rect 9769 22519 9827 22525
rect 10410 22516 10416 22528
rect 10468 22516 10474 22568
rect 11146 22516 11152 22568
rect 11204 22556 11210 22568
rect 13280 22556 13308 22596
rect 15933 22593 15945 22596
rect 15979 22624 15991 22627
rect 16945 22627 17003 22633
rect 16945 22624 16957 22627
rect 15979 22596 16957 22624
rect 15979 22593 15991 22596
rect 15933 22587 15991 22593
rect 16945 22593 16957 22596
rect 16991 22593 17003 22627
rect 16945 22587 17003 22593
rect 18506 22584 18512 22636
rect 18564 22624 18570 22636
rect 18877 22627 18935 22633
rect 18877 22624 18889 22627
rect 18564 22596 18889 22624
rect 18564 22584 18570 22596
rect 18877 22593 18889 22596
rect 18923 22593 18935 22627
rect 18877 22587 18935 22593
rect 21269 22627 21327 22633
rect 21269 22593 21281 22627
rect 21315 22593 21327 22627
rect 21269 22587 21327 22593
rect 21453 22627 21511 22633
rect 21453 22593 21465 22627
rect 21499 22624 21511 22627
rect 23106 22624 23112 22636
rect 21499 22596 23112 22624
rect 21499 22593 21511 22596
rect 21453 22587 21511 22593
rect 11204 22528 13308 22556
rect 15749 22559 15807 22565
rect 11204 22516 11210 22528
rect 15749 22525 15761 22559
rect 15795 22525 15807 22559
rect 21284 22556 21312 22587
rect 23106 22584 23112 22596
rect 23164 22624 23170 22636
rect 23385 22627 23443 22633
rect 23385 22624 23397 22627
rect 23164 22596 23397 22624
rect 23164 22584 23170 22596
rect 23385 22593 23397 22596
rect 23431 22593 23443 22627
rect 23385 22587 23443 22593
rect 24489 22627 24547 22633
rect 24489 22593 24501 22627
rect 24535 22624 24547 22627
rect 24578 22624 24584 22636
rect 24535 22596 24584 22624
rect 24535 22593 24547 22596
rect 24489 22587 24547 22593
rect 24578 22584 24584 22596
rect 24636 22584 24642 22636
rect 24762 22633 24768 22636
rect 24756 22587 24768 22633
rect 24762 22584 24768 22587
rect 24820 22584 24826 22636
rect 28350 22584 28356 22636
rect 28408 22584 28414 22636
rect 22278 22556 22284 22568
rect 21284 22528 22284 22556
rect 15749 22519 15807 22525
rect 3752 22460 5856 22488
rect 3752 22448 3758 22460
rect 13078 22448 13084 22500
rect 13136 22448 13142 22500
rect 15764 22488 15792 22519
rect 22278 22516 22284 22528
rect 22336 22556 22342 22568
rect 22465 22559 22523 22565
rect 22465 22556 22477 22559
rect 22336 22528 22477 22556
rect 22336 22516 22342 22528
rect 22465 22525 22477 22528
rect 22511 22525 22523 22559
rect 22465 22519 22523 22525
rect 22557 22559 22615 22565
rect 22557 22525 22569 22559
rect 22603 22525 22615 22559
rect 22557 22519 22615 22525
rect 16574 22488 16580 22500
rect 15764 22460 16580 22488
rect 16574 22448 16580 22460
rect 16632 22488 16638 22500
rect 17402 22488 17408 22500
rect 16632 22460 17408 22488
rect 16632 22448 16638 22460
rect 17402 22448 17408 22460
rect 17460 22448 17466 22500
rect 20346 22448 20352 22500
rect 20404 22488 20410 22500
rect 20404 22460 22232 22488
rect 20404 22448 20410 22460
rect 2225 22423 2283 22429
rect 2225 22389 2237 22423
rect 2271 22420 2283 22423
rect 3050 22420 3056 22432
rect 2271 22392 3056 22420
rect 2271 22389 2283 22392
rect 2225 22383 2283 22389
rect 3050 22380 3056 22392
rect 3108 22380 3114 22432
rect 4065 22423 4123 22429
rect 4065 22389 4077 22423
rect 4111 22420 4123 22423
rect 4154 22420 4160 22432
rect 4111 22392 4160 22420
rect 4111 22389 4123 22392
rect 4065 22383 4123 22389
rect 4154 22380 4160 22392
rect 4212 22380 4218 22432
rect 4982 22380 4988 22432
rect 5040 22420 5046 22432
rect 6822 22420 6828 22432
rect 5040 22392 6828 22420
rect 5040 22380 5046 22392
rect 6822 22380 6828 22392
rect 6880 22380 6886 22432
rect 12437 22423 12495 22429
rect 12437 22389 12449 22423
rect 12483 22420 12495 22423
rect 12526 22420 12532 22432
rect 12483 22392 12532 22420
rect 12483 22389 12495 22392
rect 12437 22383 12495 22389
rect 12526 22380 12532 22392
rect 12584 22380 12590 22432
rect 13173 22423 13231 22429
rect 13173 22389 13185 22423
rect 13219 22420 13231 22423
rect 14734 22420 14740 22432
rect 13219 22392 14740 22420
rect 13219 22389 13231 22392
rect 13173 22383 13231 22389
rect 14734 22380 14740 22392
rect 14792 22380 14798 22432
rect 15010 22380 15016 22432
rect 15068 22380 15074 22432
rect 16301 22423 16359 22429
rect 16301 22389 16313 22423
rect 16347 22420 16359 22423
rect 16666 22420 16672 22432
rect 16347 22392 16672 22420
rect 16347 22389 16359 22392
rect 16301 22383 16359 22389
rect 16666 22380 16672 22392
rect 16724 22380 16730 22432
rect 22005 22423 22063 22429
rect 22005 22389 22017 22423
rect 22051 22420 22063 22423
rect 22094 22420 22100 22432
rect 22051 22392 22100 22420
rect 22051 22389 22063 22392
rect 22005 22383 22063 22389
rect 22094 22380 22100 22392
rect 22152 22380 22158 22432
rect 22204 22420 22232 22460
rect 22572 22420 22600 22519
rect 25130 22420 25136 22432
rect 22204 22392 25136 22420
rect 25130 22380 25136 22392
rect 25188 22380 25194 22432
rect 1104 22330 30820 22352
rect 1104 22278 4664 22330
rect 4716 22278 4728 22330
rect 4780 22278 4792 22330
rect 4844 22278 4856 22330
rect 4908 22278 4920 22330
rect 4972 22278 12092 22330
rect 12144 22278 12156 22330
rect 12208 22278 12220 22330
rect 12272 22278 12284 22330
rect 12336 22278 12348 22330
rect 12400 22278 19520 22330
rect 19572 22278 19584 22330
rect 19636 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 26948 22330
rect 27000 22278 27012 22330
rect 27064 22278 27076 22330
rect 27128 22278 27140 22330
rect 27192 22278 27204 22330
rect 27256 22278 30820 22330
rect 1104 22256 30820 22278
rect 3421 22219 3479 22225
rect 3421 22185 3433 22219
rect 3467 22216 3479 22219
rect 3694 22216 3700 22228
rect 3467 22188 3700 22216
rect 3467 22185 3479 22188
rect 3421 22179 3479 22185
rect 3694 22176 3700 22188
rect 3752 22176 3758 22228
rect 5629 22219 5687 22225
rect 5629 22185 5641 22219
rect 5675 22216 5687 22219
rect 5810 22216 5816 22228
rect 5675 22188 5816 22216
rect 5675 22185 5687 22188
rect 5629 22179 5687 22185
rect 5810 22176 5816 22188
rect 5868 22176 5874 22228
rect 15565 22219 15623 22225
rect 15565 22185 15577 22219
rect 15611 22216 15623 22219
rect 15654 22216 15660 22228
rect 15611 22188 15660 22216
rect 15611 22185 15623 22188
rect 15565 22179 15623 22185
rect 15654 22176 15660 22188
rect 15712 22176 15718 22228
rect 24762 22176 24768 22228
rect 24820 22176 24826 22228
rect 5258 22108 5264 22160
rect 5316 22148 5322 22160
rect 9122 22148 9128 22160
rect 5316 22120 9128 22148
rect 5316 22108 5322 22120
rect 9122 22108 9128 22120
rect 9180 22108 9186 22160
rect 11790 22148 11796 22160
rect 11624 22120 11796 22148
rect 6822 22080 6828 22092
rect 6472 22052 6828 22080
rect 6472 22024 6500 22052
rect 6822 22040 6828 22052
rect 6880 22040 6886 22092
rect 10134 22040 10140 22092
rect 10192 22040 10198 22092
rect 10410 22040 10416 22092
rect 10468 22040 10474 22092
rect 11422 22040 11428 22092
rect 11480 22040 11486 22092
rect 11624 22089 11652 22120
rect 11790 22108 11796 22120
rect 11848 22148 11854 22160
rect 15194 22148 15200 22160
rect 11848 22120 15200 22148
rect 11848 22108 11854 22120
rect 15194 22108 15200 22120
rect 15252 22108 15258 22160
rect 11609 22083 11667 22089
rect 11609 22049 11621 22083
rect 11655 22080 11667 22083
rect 14737 22083 14795 22089
rect 11655 22052 11689 22080
rect 12176 22052 13216 22080
rect 11655 22049 11667 22052
rect 11609 22043 11667 22049
rect 2041 22015 2099 22021
rect 2041 21981 2053 22015
rect 2087 22012 2099 22015
rect 2682 22012 2688 22024
rect 2087 21984 2688 22012
rect 2087 21981 2099 21984
rect 2041 21975 2099 21981
rect 2682 21972 2688 21984
rect 2740 21972 2746 22024
rect 4982 21972 4988 22024
rect 5040 21972 5046 22024
rect 5718 21972 5724 22024
rect 5776 21972 5782 22024
rect 6086 21972 6092 22024
rect 6144 22012 6150 22024
rect 6273 22015 6331 22021
rect 6273 22012 6285 22015
rect 6144 21984 6285 22012
rect 6144 21972 6150 21984
rect 6273 21981 6285 21984
rect 6319 21981 6331 22015
rect 6273 21975 6331 21981
rect 6454 21972 6460 22024
rect 6512 21972 6518 22024
rect 10042 21972 10048 22024
rect 10100 21972 10106 22024
rect 12176 22021 12204 22052
rect 12161 22015 12219 22021
rect 12161 21981 12173 22015
rect 12207 21981 12219 22015
rect 12161 21975 12219 21981
rect 12345 22015 12403 22021
rect 12345 21981 12357 22015
rect 12391 22012 12403 22015
rect 12986 22012 12992 22024
rect 12391 21984 12992 22012
rect 12391 21981 12403 21984
rect 12345 21975 12403 21981
rect 12986 21972 12992 21984
rect 13044 21972 13050 22024
rect 13188 21956 13216 22052
rect 14737 22049 14749 22083
rect 14783 22080 14795 22083
rect 14918 22080 14924 22092
rect 14783 22052 14924 22080
rect 14783 22049 14795 22052
rect 14737 22043 14795 22049
rect 14918 22040 14924 22052
rect 14976 22040 14982 22092
rect 16945 22083 17003 22089
rect 16945 22049 16957 22083
rect 16991 22080 17003 22083
rect 18506 22080 18512 22092
rect 16991 22052 18512 22080
rect 16991 22049 17003 22052
rect 16945 22043 17003 22049
rect 14936 22012 14964 22040
rect 14936 21984 16574 22012
rect 2314 21953 2320 21956
rect 2308 21944 2320 21953
rect 2275 21916 2320 21944
rect 2308 21907 2320 21916
rect 2314 21904 2320 21907
rect 2372 21904 2378 21956
rect 4154 21904 4160 21956
rect 4212 21904 4218 21956
rect 7006 21904 7012 21956
rect 7064 21904 7070 21956
rect 13170 21904 13176 21956
rect 13228 21904 13234 21956
rect 15010 21904 15016 21956
rect 15068 21904 15074 21956
rect 16546 21944 16574 21984
rect 16666 21972 16672 22024
rect 16724 22021 16730 22024
rect 16724 21975 16736 22021
rect 16724 21972 16730 21975
rect 16960 21944 16988 22043
rect 18506 22040 18512 22052
rect 18564 22040 18570 22092
rect 20806 22040 20812 22092
rect 20864 22080 20870 22092
rect 21453 22083 21511 22089
rect 21453 22080 21465 22083
rect 20864 22052 21465 22080
rect 20864 22040 20870 22052
rect 21453 22049 21465 22052
rect 21499 22049 21511 22083
rect 21453 22043 21511 22049
rect 25130 22040 25136 22092
rect 25188 22080 25194 22092
rect 25317 22083 25375 22089
rect 25317 22080 25329 22083
rect 25188 22052 25329 22080
rect 25188 22040 25194 22052
rect 25317 22049 25329 22052
rect 25363 22049 25375 22083
rect 25317 22043 25375 22049
rect 25958 22040 25964 22092
rect 26016 22040 26022 22092
rect 26234 22040 26240 22092
rect 26292 22040 26298 22092
rect 29178 22040 29184 22092
rect 29236 22040 29242 22092
rect 17865 22015 17923 22021
rect 17865 21981 17877 22015
rect 17911 22012 17923 22015
rect 18138 22012 18144 22024
rect 17911 21984 18144 22012
rect 17911 21981 17923 21984
rect 17865 21975 17923 21981
rect 18138 21972 18144 21984
rect 18196 21972 18202 22024
rect 21174 21972 21180 22024
rect 21232 22012 21238 22024
rect 22830 22012 22836 22024
rect 21232 21984 22836 22012
rect 21232 21972 21238 21984
rect 22830 21972 22836 21984
rect 22888 21972 22894 22024
rect 25225 22015 25283 22021
rect 25225 21981 25237 22015
rect 25271 22012 25283 22015
rect 25866 22012 25872 22024
rect 25271 21984 25872 22012
rect 25271 21981 25283 21984
rect 25225 21975 25283 21981
rect 25866 21972 25872 21984
rect 25924 21972 25930 22024
rect 26329 22015 26387 22021
rect 26329 21981 26341 22015
rect 26375 22012 26387 22015
rect 27433 22015 27491 22021
rect 27433 22012 27445 22015
rect 26375 21984 27445 22012
rect 26375 21981 26387 21984
rect 26329 21975 26387 21981
rect 27433 21981 27445 21984
rect 27479 22012 27491 22015
rect 27614 22012 27620 22024
rect 27479 21984 27620 22012
rect 27479 21981 27491 21984
rect 27433 21975 27491 21981
rect 27614 21972 27620 21984
rect 27672 21972 27678 22024
rect 28166 21972 28172 22024
rect 28224 21972 28230 22024
rect 28442 21972 28448 22024
rect 28500 21972 28506 22024
rect 29362 21972 29368 22024
rect 29420 22012 29426 22024
rect 29825 22015 29883 22021
rect 29825 22012 29837 22015
rect 29420 21984 29837 22012
rect 29420 21972 29426 21984
rect 29825 21981 29837 21984
rect 29871 21981 29883 22015
rect 29825 21975 29883 21981
rect 16546 21916 16988 21944
rect 17218 21904 17224 21956
rect 17276 21944 17282 21956
rect 17589 21947 17647 21953
rect 17589 21944 17601 21947
rect 17276 21916 17601 21944
rect 17276 21904 17282 21916
rect 17589 21913 17601 21916
rect 17635 21913 17647 21947
rect 17589 21907 17647 21913
rect 22925 21947 22983 21953
rect 22925 21913 22937 21947
rect 22971 21913 22983 21947
rect 22925 21907 22983 21913
rect 23293 21947 23351 21953
rect 23293 21913 23305 21947
rect 23339 21944 23351 21947
rect 23566 21944 23572 21956
rect 23339 21916 23572 21944
rect 23339 21913 23351 21916
rect 23293 21907 23351 21913
rect 10870 21836 10876 21888
rect 10928 21876 10934 21888
rect 10965 21879 11023 21885
rect 10965 21876 10977 21879
rect 10928 21848 10977 21876
rect 10928 21836 10934 21848
rect 10965 21845 10977 21848
rect 11011 21845 11023 21879
rect 10965 21839 11023 21845
rect 11146 21836 11152 21888
rect 11204 21876 11210 21888
rect 11333 21879 11391 21885
rect 11333 21876 11345 21879
rect 11204 21848 11345 21876
rect 11204 21836 11210 21848
rect 11333 21845 11345 21848
rect 11379 21845 11391 21879
rect 11333 21839 11391 21845
rect 12250 21836 12256 21888
rect 12308 21836 12314 21888
rect 12434 21836 12440 21888
rect 12492 21876 12498 21888
rect 12805 21879 12863 21885
rect 12805 21876 12817 21879
rect 12492 21848 12817 21876
rect 12492 21836 12498 21848
rect 12805 21845 12817 21848
rect 12851 21845 12863 21879
rect 15028 21876 15056 21904
rect 22940 21876 22968 21907
rect 23566 21904 23572 21916
rect 23624 21904 23630 21956
rect 25133 21947 25191 21953
rect 25133 21913 25145 21947
rect 25179 21944 25191 21947
rect 25682 21944 25688 21956
rect 25179 21916 25688 21944
rect 25179 21913 25191 21916
rect 25133 21907 25191 21913
rect 25682 21904 25688 21916
rect 25740 21904 25746 21956
rect 30101 21947 30159 21953
rect 30101 21913 30113 21947
rect 30147 21944 30159 21947
rect 31018 21944 31024 21956
rect 30147 21916 31024 21944
rect 30147 21913 30159 21916
rect 30101 21907 30159 21913
rect 31018 21904 31024 21916
rect 31076 21904 31082 21956
rect 15028 21848 22968 21876
rect 27525 21879 27583 21885
rect 12805 21839 12863 21845
rect 27525 21845 27537 21879
rect 27571 21876 27583 21879
rect 27890 21876 27896 21888
rect 27571 21848 27896 21876
rect 27571 21845 27583 21848
rect 27525 21839 27583 21845
rect 27890 21836 27896 21848
rect 27948 21836 27954 21888
rect 1104 21786 30976 21808
rect 1104 21734 8378 21786
rect 8430 21734 8442 21786
rect 8494 21734 8506 21786
rect 8558 21734 8570 21786
rect 8622 21734 8634 21786
rect 8686 21734 15806 21786
rect 15858 21734 15870 21786
rect 15922 21734 15934 21786
rect 15986 21734 15998 21786
rect 16050 21734 16062 21786
rect 16114 21734 23234 21786
rect 23286 21734 23298 21786
rect 23350 21734 23362 21786
rect 23414 21734 23426 21786
rect 23478 21734 23490 21786
rect 23542 21734 30662 21786
rect 30714 21734 30726 21786
rect 30778 21734 30790 21786
rect 30842 21734 30854 21786
rect 30906 21734 30918 21786
rect 30970 21734 30976 21786
rect 1104 21712 30976 21734
rect 9674 21632 9680 21684
rect 9732 21672 9738 21684
rect 10413 21675 10471 21681
rect 10413 21672 10425 21675
rect 9732 21644 10425 21672
rect 9732 21632 9738 21644
rect 10413 21641 10425 21644
rect 10459 21641 10471 21675
rect 10413 21635 10471 21641
rect 12805 21675 12863 21681
rect 12805 21641 12817 21675
rect 12851 21672 12863 21675
rect 13078 21672 13084 21684
rect 12851 21644 13084 21672
rect 12851 21641 12863 21644
rect 12805 21635 12863 21641
rect 13078 21632 13084 21644
rect 13136 21632 13142 21684
rect 16853 21675 16911 21681
rect 16853 21672 16865 21675
rect 16546 21644 16865 21672
rect 4338 21564 4344 21616
rect 4396 21564 4402 21616
rect 5718 21564 5724 21616
rect 5776 21604 5782 21616
rect 8754 21604 8760 21616
rect 5776 21576 8760 21604
rect 5776 21564 5782 21576
rect 5828 21545 5856 21576
rect 8754 21564 8760 21576
rect 8812 21564 8818 21616
rect 11054 21604 11060 21616
rect 8956 21576 11060 21604
rect 5813 21539 5871 21545
rect 5813 21505 5825 21539
rect 5859 21505 5871 21539
rect 5813 21499 5871 21505
rect 6733 21539 6791 21545
rect 6733 21505 6745 21539
rect 6779 21536 6791 21539
rect 8018 21536 8024 21548
rect 6779 21508 8024 21536
rect 6779 21505 6791 21508
rect 6733 21499 6791 21505
rect 8018 21496 8024 21508
rect 8076 21536 8082 21548
rect 8956 21536 8984 21576
rect 11054 21564 11060 21576
rect 11112 21564 11118 21616
rect 12434 21564 12440 21616
rect 12492 21564 12498 21616
rect 12526 21564 12532 21616
rect 12584 21564 12590 21616
rect 16056 21607 16114 21613
rect 16056 21573 16068 21607
rect 16102 21604 16114 21607
rect 16546 21604 16574 21644
rect 16853 21641 16865 21644
rect 16899 21641 16911 21675
rect 16853 21635 16911 21641
rect 23014 21632 23020 21684
rect 23072 21672 23078 21684
rect 23385 21675 23443 21681
rect 23385 21672 23397 21675
rect 23072 21644 23397 21672
rect 23072 21632 23078 21644
rect 23385 21641 23397 21644
rect 23431 21641 23443 21675
rect 23385 21635 23443 21641
rect 25041 21675 25099 21681
rect 25041 21641 25053 21675
rect 25087 21672 25099 21675
rect 25222 21672 25228 21684
rect 25087 21644 25228 21672
rect 25087 21641 25099 21644
rect 25041 21635 25099 21641
rect 25222 21632 25228 21644
rect 25280 21632 25286 21684
rect 27614 21632 27620 21684
rect 27672 21672 27678 21684
rect 28534 21672 28540 21684
rect 27672 21644 28540 21672
rect 27672 21632 27678 21644
rect 28534 21632 28540 21644
rect 28592 21672 28598 21684
rect 29365 21675 29423 21681
rect 29365 21672 29377 21675
rect 28592 21644 29377 21672
rect 28592 21632 28598 21644
rect 29365 21641 29377 21644
rect 29411 21641 29423 21675
rect 29365 21635 29423 21641
rect 16102 21576 16574 21604
rect 16102 21573 16114 21576
rect 16056 21567 16114 21573
rect 18414 21564 18420 21616
rect 18472 21564 18478 21616
rect 22094 21564 22100 21616
rect 22152 21604 22158 21616
rect 22250 21607 22308 21613
rect 22250 21604 22262 21607
rect 22152 21576 22262 21604
rect 22152 21564 22158 21576
rect 22250 21573 22262 21576
rect 22296 21573 22308 21607
rect 22250 21567 22308 21573
rect 25133 21607 25191 21613
rect 25133 21573 25145 21607
rect 25179 21604 25191 21607
rect 26234 21604 26240 21616
rect 25179 21576 26240 21604
rect 25179 21573 25191 21576
rect 25133 21567 25191 21573
rect 26234 21564 26240 21576
rect 26292 21564 26298 21616
rect 27890 21564 27896 21616
rect 27948 21564 27954 21616
rect 9306 21545 9312 21548
rect 8076 21508 8984 21536
rect 8076 21496 8082 21508
rect 9300 21499 9312 21545
rect 9306 21496 9312 21499
rect 9364 21496 9370 21548
rect 10410 21496 10416 21548
rect 10468 21536 10474 21548
rect 12161 21539 12219 21545
rect 12161 21536 12173 21539
rect 10468 21508 12173 21536
rect 10468 21496 10474 21508
rect 12161 21505 12173 21508
rect 12207 21505 12219 21539
rect 12161 21499 12219 21505
rect 12250 21496 12256 21548
rect 12308 21536 12314 21548
rect 12308 21508 12353 21536
rect 12308 21496 12314 21508
rect 12618 21496 12624 21548
rect 12676 21545 12682 21548
rect 12676 21499 12684 21545
rect 12676 21496 12682 21499
rect 14918 21496 14924 21548
rect 14976 21536 14982 21548
rect 16301 21539 16359 21545
rect 16301 21536 16313 21539
rect 14976 21508 16313 21536
rect 14976 21496 14982 21508
rect 16301 21505 16313 21508
rect 16347 21505 16359 21539
rect 16301 21499 16359 21505
rect 17218 21496 17224 21548
rect 17276 21496 17282 21548
rect 17954 21496 17960 21548
rect 18012 21536 18018 21548
rect 18049 21539 18107 21545
rect 18049 21536 18061 21539
rect 18012 21508 18061 21536
rect 18012 21496 18018 21508
rect 18049 21505 18061 21508
rect 18095 21505 18107 21539
rect 18049 21499 18107 21505
rect 18322 21496 18328 21548
rect 18380 21496 18386 21548
rect 22005 21539 22063 21545
rect 22005 21505 22017 21539
rect 22051 21536 22063 21539
rect 23566 21536 23572 21548
rect 22051 21508 23572 21536
rect 22051 21505 22063 21508
rect 22005 21499 22063 21505
rect 23566 21496 23572 21508
rect 23624 21536 23630 21548
rect 24578 21536 24584 21548
rect 23624 21508 24584 21536
rect 23624 21496 23630 21508
rect 24578 21496 24584 21508
rect 24636 21496 24642 21548
rect 25498 21496 25504 21548
rect 25556 21536 25562 21548
rect 25869 21539 25927 21545
rect 25869 21536 25881 21539
rect 25556 21508 25881 21536
rect 25556 21496 25562 21508
rect 25869 21505 25881 21508
rect 25915 21505 25927 21539
rect 25869 21499 25927 21505
rect 28994 21496 29000 21548
rect 29052 21496 29058 21548
rect 2682 21428 2688 21480
rect 2740 21428 2746 21480
rect 6086 21428 6092 21480
rect 6144 21468 6150 21480
rect 7009 21471 7067 21477
rect 7009 21468 7021 21471
rect 6144 21440 7021 21468
rect 6144 21428 6150 21440
rect 7009 21437 7021 21440
rect 7055 21468 7067 21471
rect 7374 21468 7380 21480
rect 7055 21440 7380 21468
rect 7055 21437 7067 21440
rect 7009 21431 7067 21437
rect 7374 21428 7380 21440
rect 7432 21428 7438 21480
rect 9030 21428 9036 21480
rect 9088 21428 9094 21480
rect 17313 21471 17371 21477
rect 17313 21468 17325 21471
rect 16546 21440 17325 21468
rect 5905 21335 5963 21341
rect 5905 21301 5917 21335
rect 5951 21332 5963 21335
rect 6270 21332 6276 21344
rect 5951 21304 6276 21332
rect 5951 21301 5963 21304
rect 5905 21295 5963 21301
rect 6270 21292 6276 21304
rect 6328 21292 6334 21344
rect 13170 21292 13176 21344
rect 13228 21332 13234 21344
rect 14921 21335 14979 21341
rect 14921 21332 14933 21335
rect 13228 21304 14933 21332
rect 13228 21292 13234 21304
rect 14921 21301 14933 21304
rect 14967 21332 14979 21335
rect 16546 21332 16574 21440
rect 17313 21437 17325 21440
rect 17359 21437 17371 21471
rect 17313 21431 17371 21437
rect 17402 21428 17408 21480
rect 17460 21428 17466 21480
rect 25130 21428 25136 21480
rect 25188 21468 25194 21480
rect 25225 21471 25283 21477
rect 25225 21468 25237 21471
rect 25188 21440 25237 21468
rect 25188 21428 25194 21440
rect 25225 21437 25237 21440
rect 25271 21437 25283 21471
rect 25225 21431 25283 21437
rect 25314 21428 25320 21480
rect 25372 21468 25378 21480
rect 26053 21471 26111 21477
rect 26053 21468 26065 21471
rect 25372 21440 26065 21468
rect 25372 21428 25378 21440
rect 26053 21437 26065 21440
rect 26099 21437 26111 21471
rect 26053 21431 26111 21437
rect 27614 21428 27620 21480
rect 27672 21428 27678 21480
rect 24854 21360 24860 21412
rect 24912 21400 24918 21412
rect 26142 21400 26148 21412
rect 24912 21372 26148 21400
rect 24912 21360 24918 21372
rect 26142 21360 26148 21372
rect 26200 21400 26206 21412
rect 26694 21400 26700 21412
rect 26200 21372 26700 21400
rect 26200 21360 26206 21372
rect 26694 21360 26700 21372
rect 26752 21360 26758 21412
rect 14967 21304 16574 21332
rect 14967 21301 14979 21304
rect 14921 21295 14979 21301
rect 20162 21292 20168 21344
rect 20220 21332 20226 21344
rect 22646 21332 22652 21344
rect 20220 21304 22652 21332
rect 20220 21292 20226 21304
rect 22646 21292 22652 21304
rect 22704 21292 22710 21344
rect 24670 21292 24676 21344
rect 24728 21292 24734 21344
rect 1104 21242 30820 21264
rect 1104 21190 4664 21242
rect 4716 21190 4728 21242
rect 4780 21190 4792 21242
rect 4844 21190 4856 21242
rect 4908 21190 4920 21242
rect 4972 21190 12092 21242
rect 12144 21190 12156 21242
rect 12208 21190 12220 21242
rect 12272 21190 12284 21242
rect 12336 21190 12348 21242
rect 12400 21190 19520 21242
rect 19572 21190 19584 21242
rect 19636 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 26948 21242
rect 27000 21190 27012 21242
rect 27064 21190 27076 21242
rect 27128 21190 27140 21242
rect 27192 21190 27204 21242
rect 27256 21190 30820 21242
rect 1104 21168 30820 21190
rect 2958 21088 2964 21140
rect 3016 21088 3022 21140
rect 3326 21088 3332 21140
rect 3384 21088 3390 21140
rect 13814 21128 13820 21140
rect 4356 21100 13820 21128
rect 2682 20952 2688 21004
rect 2740 20992 2746 21004
rect 4356 21001 4384 21100
rect 13814 21088 13820 21100
rect 13872 21088 13878 21140
rect 14550 21088 14556 21140
rect 14608 21088 14614 21140
rect 15194 21088 15200 21140
rect 15252 21128 15258 21140
rect 16485 21131 16543 21137
rect 16485 21128 16497 21131
rect 15252 21100 16497 21128
rect 15252 21088 15258 21100
rect 16485 21097 16497 21100
rect 16531 21097 16543 21131
rect 16485 21091 16543 21097
rect 17773 21131 17831 21137
rect 17773 21097 17785 21131
rect 17819 21128 17831 21131
rect 18046 21128 18052 21140
rect 17819 21100 18052 21128
rect 17819 21097 17831 21100
rect 17773 21091 17831 21097
rect 18046 21088 18052 21100
rect 18104 21088 18110 21140
rect 22186 21128 22192 21140
rect 18708 21100 22192 21128
rect 7745 21063 7803 21069
rect 7745 21029 7757 21063
rect 7791 21060 7803 21063
rect 8754 21060 8760 21072
rect 7791 21032 8760 21060
rect 7791 21029 7803 21032
rect 7745 21023 7803 21029
rect 8754 21020 8760 21032
rect 8812 21020 8818 21072
rect 9306 21020 9312 21072
rect 9364 21060 9370 21072
rect 9401 21063 9459 21069
rect 9401 21060 9413 21063
rect 9364 21032 9413 21060
rect 9364 21020 9370 21032
rect 9401 21029 9413 21032
rect 9447 21029 9459 21063
rect 9401 21023 9459 21029
rect 12529 21063 12587 21069
rect 12529 21029 12541 21063
rect 12575 21060 12587 21063
rect 12618 21060 12624 21072
rect 12575 21032 12624 21060
rect 12575 21029 12587 21032
rect 12529 21023 12587 21029
rect 12618 21020 12624 21032
rect 12676 21020 12682 21072
rect 18708 21069 18736 21100
rect 22186 21088 22192 21100
rect 22244 21088 22250 21140
rect 24854 21128 24860 21140
rect 24504 21100 24860 21128
rect 18693 21063 18751 21069
rect 18693 21029 18705 21063
rect 18739 21029 18751 21063
rect 18693 21023 18751 21029
rect 20162 21020 20168 21072
rect 20220 21020 20226 21072
rect 4341 20995 4399 21001
rect 2740 20964 4200 20992
rect 2740 20952 2746 20964
rect 3050 20884 3056 20936
rect 3108 20924 3114 20936
rect 3145 20927 3203 20933
rect 3145 20924 3157 20927
rect 3108 20896 3157 20924
rect 3108 20884 3114 20896
rect 3145 20893 3157 20896
rect 3191 20893 3203 20927
rect 3145 20887 3203 20893
rect 3421 20927 3479 20933
rect 3421 20893 3433 20927
rect 3467 20893 3479 20927
rect 3421 20887 3479 20893
rect 3436 20856 3464 20887
rect 3970 20884 3976 20936
rect 4028 20884 4034 20936
rect 4172 20933 4200 20964
rect 4341 20961 4353 20995
rect 4387 20961 4399 20995
rect 4341 20955 4399 20961
rect 5445 20995 5503 21001
rect 5445 20961 5457 20995
rect 5491 20992 5503 20995
rect 5997 20995 6055 21001
rect 5997 20992 6009 20995
rect 5491 20964 6009 20992
rect 5491 20961 5503 20964
rect 5445 20955 5503 20961
rect 5997 20961 6009 20964
rect 6043 20961 6055 20995
rect 5997 20955 6055 20961
rect 6270 20952 6276 21004
rect 6328 20952 6334 21004
rect 9674 20952 9680 21004
rect 9732 20992 9738 21004
rect 9861 20995 9919 21001
rect 9861 20992 9873 20995
rect 9732 20964 9873 20992
rect 9732 20952 9738 20964
rect 9861 20961 9873 20964
rect 9907 20961 9919 20995
rect 9861 20955 9919 20961
rect 9950 20952 9956 21004
rect 10008 20952 10014 21004
rect 14996 20995 15054 21001
rect 14996 20961 15008 20995
rect 15042 20992 15054 20995
rect 18233 20995 18291 21001
rect 15042 20964 17908 20992
rect 15042 20961 15054 20964
rect 14996 20955 15054 20961
rect 4157 20927 4215 20933
rect 4157 20893 4169 20927
rect 4203 20893 4215 20927
rect 4157 20887 4215 20893
rect 5534 20884 5540 20936
rect 5592 20884 5598 20936
rect 10594 20884 10600 20936
rect 10652 20884 10658 20936
rect 10870 20933 10876 20936
rect 10864 20887 10876 20933
rect 10870 20884 10876 20887
rect 10928 20884 10934 20936
rect 12443 20927 12501 20933
rect 12443 20893 12455 20927
rect 12489 20893 12501 20927
rect 12443 20887 12501 20893
rect 12621 20927 12679 20933
rect 12621 20893 12633 20927
rect 12667 20924 12679 20927
rect 12710 20924 12716 20936
rect 12667 20896 12716 20924
rect 12667 20893 12679 20896
rect 12621 20887 12679 20893
rect 3436 20828 4200 20856
rect 4172 20800 4200 20828
rect 7006 20816 7012 20868
rect 7064 20816 7070 20868
rect 9769 20859 9827 20865
rect 9769 20825 9781 20859
rect 9815 20856 9827 20859
rect 11698 20856 11704 20868
rect 9815 20828 11704 20856
rect 9815 20825 9827 20828
rect 9769 20819 9827 20825
rect 11698 20816 11704 20828
rect 11756 20816 11762 20868
rect 12452 20856 12480 20887
rect 12710 20884 12716 20896
rect 12768 20884 12774 20936
rect 14734 20884 14740 20936
rect 14792 20884 14798 20936
rect 15286 20884 15292 20936
rect 15344 20884 15350 20936
rect 15841 20927 15899 20933
rect 15841 20893 15853 20927
rect 15887 20893 15899 20927
rect 15841 20887 15899 20893
rect 16577 20927 16635 20933
rect 16577 20893 16589 20927
rect 16623 20893 16635 20927
rect 16577 20887 16635 20893
rect 15856 20856 15884 20887
rect 16482 20856 16488 20868
rect 11992 20828 12480 20856
rect 15212 20828 16488 20856
rect 4154 20748 4160 20800
rect 4212 20748 4218 20800
rect 11422 20748 11428 20800
rect 11480 20788 11486 20800
rect 11992 20797 12020 20828
rect 15212 20800 15240 20828
rect 16482 20816 16488 20828
rect 16540 20816 16546 20868
rect 16592 20856 16620 20887
rect 17494 20884 17500 20936
rect 17552 20884 17558 20936
rect 17589 20927 17647 20933
rect 17589 20893 17601 20927
rect 17635 20893 17647 20927
rect 17589 20887 17647 20893
rect 17604 20856 17632 20887
rect 17880 20868 17908 20964
rect 18233 20961 18245 20995
rect 18279 20992 18291 20995
rect 18279 20964 21036 20992
rect 18279 20961 18291 20964
rect 18233 20955 18291 20961
rect 18417 20927 18475 20933
rect 18417 20893 18429 20927
rect 18463 20893 18475 20927
rect 18417 20887 18475 20893
rect 16592 20828 17632 20856
rect 11977 20791 12035 20797
rect 11977 20788 11989 20791
rect 11480 20760 11989 20788
rect 11480 20748 11486 20760
rect 11977 20757 11989 20760
rect 12023 20757 12035 20791
rect 11977 20751 12035 20757
rect 14918 20748 14924 20800
rect 14976 20788 14982 20800
rect 15105 20791 15163 20797
rect 15105 20788 15117 20791
rect 14976 20760 15117 20788
rect 14976 20748 14982 20760
rect 15105 20757 15117 20760
rect 15151 20757 15163 20791
rect 15105 20751 15163 20757
rect 15194 20748 15200 20800
rect 15252 20748 15258 20800
rect 17604 20788 17632 20828
rect 17862 20816 17868 20868
rect 17920 20856 17926 20868
rect 18432 20856 18460 20887
rect 18782 20884 18788 20936
rect 18840 20884 18846 20936
rect 19426 20884 19432 20936
rect 19484 20924 19490 20936
rect 19521 20927 19579 20933
rect 19521 20924 19533 20927
rect 19484 20896 19533 20924
rect 19484 20884 19490 20896
rect 19521 20893 19533 20896
rect 19567 20893 19579 20927
rect 19521 20887 19579 20893
rect 19978 20884 19984 20936
rect 20036 20884 20042 20936
rect 20898 20884 20904 20936
rect 20956 20884 20962 20936
rect 21008 20924 21036 20964
rect 24504 20924 24532 21100
rect 24854 21088 24860 21100
rect 24912 21088 24918 21140
rect 25961 21131 26019 21137
rect 25961 21097 25973 21131
rect 26007 21128 26019 21131
rect 26234 21128 26240 21140
rect 26007 21100 26240 21128
rect 26007 21097 26019 21100
rect 25961 21091 26019 21097
rect 26234 21088 26240 21100
rect 26292 21088 26298 21140
rect 26881 21131 26939 21137
rect 26881 21097 26893 21131
rect 26927 21128 26939 21131
rect 27614 21128 27620 21140
rect 26927 21100 27620 21128
rect 26927 21097 26939 21100
rect 26881 21091 26939 21097
rect 27614 21088 27620 21100
rect 27672 21088 27678 21140
rect 29822 21060 29828 21072
rect 26206 21032 29828 21060
rect 21008 20896 24532 20924
rect 24578 20884 24584 20936
rect 24636 20884 24642 20936
rect 24670 20884 24676 20936
rect 24728 20924 24734 20936
rect 24837 20927 24895 20933
rect 24837 20924 24849 20927
rect 24728 20896 24849 20924
rect 24728 20884 24734 20896
rect 24837 20893 24849 20896
rect 24883 20893 24895 20927
rect 24837 20887 24895 20893
rect 17920 20828 18460 20856
rect 21168 20859 21226 20865
rect 17920 20816 17926 20828
rect 21168 20825 21180 20859
rect 21214 20856 21226 20859
rect 21266 20856 21272 20868
rect 21214 20828 21272 20856
rect 21214 20825 21226 20828
rect 21168 20819 21226 20825
rect 21266 20816 21272 20828
rect 21324 20856 21330 20868
rect 22186 20856 22192 20868
rect 21324 20828 22192 20856
rect 21324 20816 21330 20828
rect 22186 20816 22192 20828
rect 22244 20816 22250 20868
rect 26206 20856 26234 21032
rect 29822 21020 29828 21032
rect 29880 21020 29886 21072
rect 28166 20952 28172 21004
rect 28224 20952 28230 21004
rect 28994 20952 29000 21004
rect 29052 20952 29058 21004
rect 26789 20927 26847 20933
rect 26789 20893 26801 20927
rect 26835 20893 26847 20927
rect 26789 20887 26847 20893
rect 22296 20828 26234 20856
rect 17954 20788 17960 20800
rect 17604 20760 17960 20788
rect 17954 20748 17960 20760
rect 18012 20748 18018 20800
rect 22296 20797 22324 20828
rect 22281 20791 22339 20797
rect 22281 20757 22293 20791
rect 22327 20757 22339 20791
rect 22281 20751 22339 20757
rect 22370 20748 22376 20800
rect 22428 20788 22434 20800
rect 23106 20788 23112 20800
rect 22428 20760 23112 20788
rect 22428 20748 22434 20760
rect 23106 20748 23112 20760
rect 23164 20788 23170 20800
rect 26804 20788 26832 20887
rect 28442 20884 28448 20936
rect 28500 20884 28506 20936
rect 23164 20760 26832 20788
rect 23164 20748 23170 20760
rect 1104 20698 30976 20720
rect 1104 20646 8378 20698
rect 8430 20646 8442 20698
rect 8494 20646 8506 20698
rect 8558 20646 8570 20698
rect 8622 20646 8634 20698
rect 8686 20646 15806 20698
rect 15858 20646 15870 20698
rect 15922 20646 15934 20698
rect 15986 20646 15998 20698
rect 16050 20646 16062 20698
rect 16114 20646 23234 20698
rect 23286 20646 23298 20698
rect 23350 20646 23362 20698
rect 23414 20646 23426 20698
rect 23478 20646 23490 20698
rect 23542 20646 30662 20698
rect 30714 20646 30726 20698
rect 30778 20646 30790 20698
rect 30842 20646 30854 20698
rect 30906 20646 30918 20698
rect 30970 20646 30976 20698
rect 1104 20624 30976 20646
rect 5534 20544 5540 20596
rect 5592 20584 5598 20596
rect 8297 20587 8355 20593
rect 8297 20584 8309 20587
rect 5592 20556 8309 20584
rect 5592 20544 5598 20556
rect 4062 20516 4068 20528
rect 4002 20488 4068 20516
rect 4062 20476 4068 20488
rect 4120 20476 4126 20528
rect 5828 20457 5856 20556
rect 8297 20553 8309 20556
rect 8343 20584 8355 20587
rect 10042 20584 10048 20596
rect 8343 20556 10048 20584
rect 8343 20553 8355 20556
rect 8297 20547 8355 20553
rect 10042 20544 10048 20556
rect 10100 20544 10106 20596
rect 10134 20544 10140 20596
rect 10192 20584 10198 20596
rect 10413 20587 10471 20593
rect 10413 20584 10425 20587
rect 10192 20556 10425 20584
rect 10192 20544 10198 20556
rect 10413 20553 10425 20556
rect 10459 20553 10471 20587
rect 10413 20547 10471 20553
rect 15286 20544 15292 20596
rect 15344 20584 15350 20596
rect 15473 20587 15531 20593
rect 15473 20584 15485 20587
rect 15344 20556 15485 20584
rect 15344 20544 15350 20556
rect 15473 20553 15485 20556
rect 15519 20553 15531 20587
rect 15473 20547 15531 20553
rect 15654 20544 15660 20596
rect 15712 20584 15718 20596
rect 18601 20587 18659 20593
rect 15712 20556 18552 20584
rect 15712 20544 15718 20556
rect 5905 20519 5963 20525
rect 5905 20485 5917 20519
rect 5951 20516 5963 20519
rect 6825 20519 6883 20525
rect 6825 20516 6837 20519
rect 5951 20488 6837 20516
rect 5951 20485 5963 20488
rect 5905 20479 5963 20485
rect 6825 20485 6837 20488
rect 6871 20485 6883 20519
rect 6825 20479 6883 20485
rect 7098 20476 7104 20528
rect 7156 20516 7162 20528
rect 7156 20488 7314 20516
rect 8128 20488 9444 20516
rect 7156 20476 7162 20488
rect 4709 20451 4767 20457
rect 4709 20448 4721 20451
rect 4264 20420 4721 20448
rect 2498 20340 2504 20392
rect 2556 20340 2562 20392
rect 2777 20383 2835 20389
rect 2777 20349 2789 20383
rect 2823 20380 2835 20383
rect 3970 20380 3976 20392
rect 2823 20352 3976 20380
rect 2823 20349 2835 20352
rect 2777 20343 2835 20349
rect 3970 20340 3976 20352
rect 4028 20340 4034 20392
rect 4264 20389 4292 20420
rect 4709 20417 4721 20420
rect 4755 20417 4767 20451
rect 4709 20411 4767 20417
rect 5813 20451 5871 20457
rect 5813 20417 5825 20451
rect 5859 20417 5871 20451
rect 5813 20411 5871 20417
rect 4249 20383 4307 20389
rect 4249 20349 4261 20383
rect 4295 20349 4307 20383
rect 4249 20343 4307 20349
rect 6546 20340 6552 20392
rect 6604 20340 6610 20392
rect 7190 20340 7196 20392
rect 7248 20380 7254 20392
rect 8128 20380 8156 20488
rect 9306 20457 9312 20460
rect 9300 20411 9312 20457
rect 9306 20408 9312 20411
rect 9364 20408 9370 20460
rect 9416 20448 9444 20488
rect 9950 20476 9956 20528
rect 10008 20516 10014 20528
rect 15194 20516 15200 20528
rect 10008 20488 12434 20516
rect 10008 20476 10014 20488
rect 12406 20448 12434 20488
rect 14476 20488 15200 20516
rect 14476 20457 14504 20488
rect 15194 20476 15200 20488
rect 15252 20476 15258 20528
rect 15304 20488 18368 20516
rect 14277 20451 14335 20457
rect 14277 20448 14289 20451
rect 9416 20420 10088 20448
rect 12406 20420 14289 20448
rect 7248 20352 8156 20380
rect 9033 20383 9091 20389
rect 7248 20340 7254 20352
rect 9033 20349 9045 20383
rect 9079 20349 9091 20383
rect 10060 20380 10088 20420
rect 14277 20417 14289 20420
rect 14323 20417 14335 20451
rect 14277 20411 14335 20417
rect 14461 20451 14519 20457
rect 14461 20417 14473 20451
rect 14507 20417 14519 20451
rect 14461 20411 14519 20417
rect 14642 20408 14648 20460
rect 14700 20448 14706 20460
rect 15304 20448 15332 20488
rect 14700 20420 15332 20448
rect 14700 20408 14706 20420
rect 15562 20408 15568 20460
rect 15620 20408 15626 20460
rect 16482 20408 16488 20460
rect 16540 20448 16546 20460
rect 16853 20451 16911 20457
rect 16853 20448 16865 20451
rect 16540 20420 16865 20448
rect 16540 20408 16546 20420
rect 16853 20417 16865 20420
rect 16899 20417 16911 20451
rect 16853 20411 16911 20417
rect 17129 20451 17187 20457
rect 17129 20417 17141 20451
rect 17175 20417 17187 20451
rect 17129 20411 17187 20417
rect 17221 20451 17279 20457
rect 17221 20417 17233 20451
rect 17267 20448 17279 20451
rect 17402 20448 17408 20460
rect 17267 20420 17408 20448
rect 17267 20417 17279 20420
rect 17221 20411 17279 20417
rect 17144 20380 17172 20411
rect 17402 20408 17408 20420
rect 17460 20408 17466 20460
rect 18340 20448 18368 20488
rect 18414 20476 18420 20528
rect 18472 20476 18478 20528
rect 18524 20516 18552 20556
rect 18601 20553 18613 20587
rect 18647 20584 18659 20587
rect 18782 20584 18788 20596
rect 18647 20556 18788 20584
rect 18647 20553 18659 20556
rect 18601 20547 18659 20553
rect 18782 20544 18788 20556
rect 18840 20544 18846 20596
rect 19889 20587 19947 20593
rect 19889 20553 19901 20587
rect 19935 20584 19947 20587
rect 20898 20584 20904 20596
rect 19935 20556 20904 20584
rect 19935 20553 19947 20556
rect 19889 20547 19947 20553
rect 20898 20544 20904 20556
rect 20956 20544 20962 20596
rect 23566 20516 23572 20528
rect 18524 20488 23572 20516
rect 23566 20476 23572 20488
rect 23624 20516 23630 20528
rect 23624 20488 24532 20516
rect 23624 20476 23630 20488
rect 19705 20451 19763 20457
rect 19705 20448 19717 20451
rect 18340 20420 19717 20448
rect 19705 20417 19717 20420
rect 19751 20448 19763 20451
rect 19978 20448 19984 20460
rect 19751 20420 19984 20448
rect 19751 20417 19763 20420
rect 19705 20411 19763 20417
rect 19978 20408 19984 20420
rect 20036 20408 20042 20460
rect 20806 20408 20812 20460
rect 20864 20408 20870 20460
rect 21082 20408 21088 20460
rect 21140 20408 21146 20460
rect 22189 20451 22247 20457
rect 22189 20417 22201 20451
rect 22235 20448 22247 20451
rect 22370 20448 22376 20460
rect 22235 20420 22376 20448
rect 22235 20417 22247 20420
rect 22189 20411 22247 20417
rect 22370 20408 22376 20420
rect 22428 20408 22434 20460
rect 24504 20457 24532 20488
rect 24489 20451 24547 20457
rect 24489 20417 24501 20451
rect 24535 20417 24547 20451
rect 24489 20411 24547 20417
rect 24578 20408 24584 20460
rect 24636 20448 24642 20460
rect 24673 20451 24731 20457
rect 24673 20448 24685 20451
rect 24636 20420 24685 20448
rect 24636 20408 24642 20420
rect 24673 20417 24685 20420
rect 24719 20417 24731 20451
rect 24673 20411 24731 20417
rect 10060 20352 12434 20380
rect 17144 20352 17264 20380
rect 9033 20343 9091 20349
rect 3988 20312 4016 20340
rect 4801 20315 4859 20321
rect 4801 20312 4813 20315
rect 3988 20284 4813 20312
rect 4801 20281 4813 20284
rect 4847 20281 4859 20315
rect 4801 20275 4859 20281
rect 9048 20244 9076 20343
rect 9766 20244 9772 20256
rect 9048 20216 9772 20244
rect 9766 20204 9772 20216
rect 9824 20244 9830 20256
rect 10594 20244 10600 20256
rect 9824 20216 10600 20244
rect 9824 20204 9830 20216
rect 10594 20204 10600 20216
rect 10652 20204 10658 20256
rect 12406 20244 12434 20352
rect 17236 20312 17264 20352
rect 17494 20340 17500 20392
rect 17552 20380 17558 20392
rect 17678 20380 17684 20392
rect 17552 20352 17684 20380
rect 17552 20340 17558 20352
rect 17678 20340 17684 20352
rect 17736 20380 17742 20392
rect 19521 20383 19579 20389
rect 19521 20380 19533 20383
rect 17736 20352 19533 20380
rect 17736 20340 17742 20352
rect 19521 20349 19533 20352
rect 19567 20380 19579 20383
rect 19886 20380 19892 20392
rect 19567 20352 19892 20380
rect 19567 20349 19579 20352
rect 19521 20343 19579 20349
rect 19886 20340 19892 20352
rect 19944 20340 19950 20392
rect 21358 20340 21364 20392
rect 21416 20340 21422 20392
rect 17770 20312 17776 20324
rect 17236 20284 17776 20312
rect 17770 20272 17776 20284
rect 17828 20312 17834 20324
rect 18049 20315 18107 20321
rect 18049 20312 18061 20315
rect 17828 20284 18061 20312
rect 17828 20272 17834 20284
rect 18049 20281 18061 20284
rect 18095 20281 18107 20315
rect 18049 20275 18107 20281
rect 15654 20244 15660 20256
rect 12406 20216 15660 20244
rect 15654 20204 15660 20216
rect 15712 20204 15718 20256
rect 18322 20204 18328 20256
rect 18380 20244 18386 20256
rect 18417 20247 18475 20253
rect 18417 20244 18429 20247
rect 18380 20216 18429 20244
rect 18380 20204 18386 20216
rect 18417 20213 18429 20216
rect 18463 20213 18475 20247
rect 18417 20207 18475 20213
rect 22094 20204 22100 20256
rect 22152 20204 22158 20256
rect 24581 20247 24639 20253
rect 24581 20213 24593 20247
rect 24627 20244 24639 20247
rect 25314 20244 25320 20256
rect 24627 20216 25320 20244
rect 24627 20213 24639 20216
rect 24581 20207 24639 20213
rect 25314 20204 25320 20216
rect 25372 20204 25378 20256
rect 1104 20154 30820 20176
rect 1104 20102 4664 20154
rect 4716 20102 4728 20154
rect 4780 20102 4792 20154
rect 4844 20102 4856 20154
rect 4908 20102 4920 20154
rect 4972 20102 12092 20154
rect 12144 20102 12156 20154
rect 12208 20102 12220 20154
rect 12272 20102 12284 20154
rect 12336 20102 12348 20154
rect 12400 20102 19520 20154
rect 19572 20102 19584 20154
rect 19636 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 26948 20154
rect 27000 20102 27012 20154
rect 27064 20102 27076 20154
rect 27128 20102 27140 20154
rect 27192 20102 27204 20154
rect 27256 20102 30820 20154
rect 1104 20080 30820 20102
rect 2498 20000 2504 20052
rect 2556 20040 2562 20052
rect 3145 20043 3203 20049
rect 3145 20040 3157 20043
rect 2556 20012 3157 20040
rect 2556 20000 2562 20012
rect 3145 20009 3157 20012
rect 3191 20009 3203 20043
rect 3145 20003 3203 20009
rect 4062 20000 4068 20052
rect 4120 20000 4126 20052
rect 9306 20000 9312 20052
rect 9364 20040 9370 20052
rect 9493 20043 9551 20049
rect 9493 20040 9505 20043
rect 9364 20012 9505 20040
rect 9364 20000 9370 20012
rect 9493 20009 9505 20012
rect 9539 20009 9551 20043
rect 9493 20003 9551 20009
rect 18506 20000 18512 20052
rect 18564 20040 18570 20052
rect 18877 20043 18935 20049
rect 18877 20040 18889 20043
rect 18564 20012 18889 20040
rect 18564 20000 18570 20012
rect 18877 20009 18889 20012
rect 18923 20040 18935 20043
rect 27982 20040 27988 20052
rect 18923 20012 27988 20040
rect 18923 20009 18935 20012
rect 18877 20003 18935 20009
rect 27982 20000 27988 20012
rect 28040 20000 28046 20052
rect 9950 19932 9956 19984
rect 10008 19972 10014 19984
rect 22189 19975 22247 19981
rect 10008 19944 10088 19972
rect 10008 19932 10014 19944
rect 7098 19864 7104 19916
rect 7156 19864 7162 19916
rect 10060 19913 10088 19944
rect 22189 19941 22201 19975
rect 22235 19972 22247 19975
rect 22370 19972 22376 19984
rect 22235 19944 22376 19972
rect 22235 19941 22247 19944
rect 22189 19935 22247 19941
rect 22370 19932 22376 19944
rect 22428 19932 22434 19984
rect 10045 19907 10103 19913
rect 10045 19873 10057 19907
rect 10091 19873 10103 19907
rect 10045 19867 10103 19873
rect 14734 19864 14740 19916
rect 14792 19904 14798 19916
rect 17497 19907 17555 19913
rect 17497 19904 17509 19907
rect 14792 19876 17509 19904
rect 14792 19864 14798 19876
rect 17497 19873 17509 19876
rect 17543 19873 17555 19907
rect 17497 19867 17555 19873
rect 18966 19864 18972 19916
rect 19024 19904 19030 19916
rect 19889 19907 19947 19913
rect 19024 19876 19748 19904
rect 19024 19864 19030 19876
rect 2593 19839 2651 19845
rect 2593 19805 2605 19839
rect 2639 19836 2651 19839
rect 3237 19839 3295 19845
rect 3237 19836 3249 19839
rect 2639 19808 3249 19836
rect 2639 19805 2651 19808
rect 2593 19799 2651 19805
rect 3237 19805 3249 19808
rect 3283 19836 3295 19839
rect 3878 19836 3884 19848
rect 3283 19808 3884 19836
rect 3283 19805 3295 19808
rect 3237 19799 3295 19805
rect 3878 19796 3884 19808
rect 3936 19796 3942 19848
rect 4154 19796 4160 19848
rect 4212 19796 4218 19848
rect 5258 19796 5264 19848
rect 5316 19796 5322 19848
rect 6086 19796 6092 19848
rect 6144 19796 6150 19848
rect 6454 19796 6460 19848
rect 6512 19796 6518 19848
rect 9858 19796 9864 19848
rect 9916 19796 9922 19848
rect 9953 19839 10011 19845
rect 9953 19805 9965 19839
rect 9999 19836 10011 19839
rect 10134 19836 10140 19848
rect 9999 19808 10140 19836
rect 9999 19805 10011 19808
rect 9953 19799 10011 19805
rect 10134 19796 10140 19808
rect 10192 19796 10198 19848
rect 18322 19796 18328 19848
rect 18380 19836 18386 19848
rect 19426 19836 19432 19848
rect 18380 19808 19432 19836
rect 18380 19796 18386 19808
rect 19426 19796 19432 19808
rect 19484 19836 19490 19848
rect 19720 19845 19748 19876
rect 19889 19873 19901 19907
rect 19935 19904 19947 19907
rect 20346 19904 20352 19916
rect 19935 19876 20352 19904
rect 19935 19873 19947 19876
rect 19889 19867 19947 19873
rect 20346 19864 20352 19876
rect 20404 19864 20410 19916
rect 20717 19907 20775 19913
rect 20717 19873 20729 19907
rect 20763 19904 20775 19907
rect 22094 19904 22100 19916
rect 20763 19876 22100 19904
rect 20763 19873 20775 19876
rect 20717 19867 20775 19873
rect 22094 19864 22100 19876
rect 22152 19864 22158 19916
rect 25317 19907 25375 19913
rect 25317 19873 25329 19907
rect 25363 19904 25375 19907
rect 25406 19904 25412 19916
rect 25363 19876 25412 19904
rect 25363 19873 25375 19876
rect 25317 19867 25375 19873
rect 25406 19864 25412 19876
rect 25464 19864 25470 19916
rect 26694 19864 26700 19916
rect 26752 19904 26758 19916
rect 27249 19907 27307 19913
rect 27249 19904 27261 19907
rect 26752 19876 27261 19904
rect 26752 19864 26758 19876
rect 27249 19873 27261 19876
rect 27295 19873 27307 19907
rect 27249 19867 27307 19873
rect 19521 19839 19579 19845
rect 19521 19836 19533 19839
rect 19484 19808 19533 19836
rect 19484 19796 19490 19808
rect 19521 19805 19533 19808
rect 19567 19805 19579 19839
rect 19521 19799 19579 19805
rect 19705 19839 19763 19845
rect 19705 19805 19717 19839
rect 19751 19805 19763 19839
rect 20441 19839 20499 19845
rect 20441 19836 20453 19839
rect 19705 19799 19763 19805
rect 19812 19808 20453 19836
rect 9876 19768 9904 19796
rect 17218 19768 17224 19780
rect 9876 19740 17224 19768
rect 17218 19728 17224 19740
rect 17276 19768 17282 19780
rect 17586 19768 17592 19780
rect 17276 19740 17592 19768
rect 17276 19728 17282 19740
rect 17586 19728 17592 19740
rect 17644 19728 17650 19780
rect 17764 19771 17822 19777
rect 17764 19737 17776 19771
rect 17810 19768 17822 19771
rect 18414 19768 18420 19780
rect 17810 19740 18420 19768
rect 17810 19737 17822 19740
rect 17764 19731 17822 19737
rect 18414 19728 18420 19740
rect 18472 19728 18478 19780
rect 2130 19660 2136 19712
rect 2188 19700 2194 19712
rect 2501 19703 2559 19709
rect 2501 19700 2513 19703
rect 2188 19672 2513 19700
rect 2188 19660 2194 19672
rect 2501 19669 2513 19672
rect 2547 19669 2559 19703
rect 2501 19663 2559 19669
rect 5445 19703 5503 19709
rect 5445 19669 5457 19703
rect 5491 19700 5503 19703
rect 6178 19700 6184 19712
rect 5491 19672 6184 19700
rect 5491 19669 5503 19672
rect 5445 19663 5503 19669
rect 6178 19660 6184 19672
rect 6236 19660 6242 19712
rect 6546 19660 6552 19712
rect 6604 19700 6610 19712
rect 10870 19700 10876 19712
rect 6604 19672 10876 19700
rect 6604 19660 6610 19672
rect 10870 19660 10876 19672
rect 10928 19700 10934 19712
rect 19812 19700 19840 19808
rect 20441 19805 20453 19808
rect 20487 19805 20499 19839
rect 20441 19799 20499 19805
rect 21358 19728 21364 19780
rect 21416 19728 21422 19780
rect 22002 19728 22008 19780
rect 22060 19768 22066 19780
rect 25041 19771 25099 19777
rect 25041 19768 25053 19771
rect 22060 19740 25053 19768
rect 22060 19728 22066 19740
rect 25041 19737 25053 19740
rect 25087 19737 25099 19771
rect 25041 19731 25099 19737
rect 27516 19771 27574 19777
rect 27516 19737 27528 19771
rect 27562 19768 27574 19771
rect 28442 19768 28448 19780
rect 27562 19740 28448 19768
rect 27562 19737 27574 19740
rect 27516 19731 27574 19737
rect 28442 19728 28448 19740
rect 28500 19728 28506 19780
rect 10928 19672 19840 19700
rect 10928 19660 10934 19672
rect 24670 19660 24676 19712
rect 24728 19660 24734 19712
rect 25133 19703 25191 19709
rect 25133 19669 25145 19703
rect 25179 19700 25191 19703
rect 25866 19700 25872 19712
rect 25179 19672 25872 19700
rect 25179 19669 25191 19672
rect 25133 19663 25191 19669
rect 25866 19660 25872 19672
rect 25924 19660 25930 19712
rect 28626 19660 28632 19712
rect 28684 19660 28690 19712
rect 1104 19610 30976 19632
rect 1104 19558 8378 19610
rect 8430 19558 8442 19610
rect 8494 19558 8506 19610
rect 8558 19558 8570 19610
rect 8622 19558 8634 19610
rect 8686 19558 15806 19610
rect 15858 19558 15870 19610
rect 15922 19558 15934 19610
rect 15986 19558 15998 19610
rect 16050 19558 16062 19610
rect 16114 19558 23234 19610
rect 23286 19558 23298 19610
rect 23350 19558 23362 19610
rect 23414 19558 23426 19610
rect 23478 19558 23490 19610
rect 23542 19558 30662 19610
rect 30714 19558 30726 19610
rect 30778 19558 30790 19610
rect 30842 19558 30854 19610
rect 30906 19558 30918 19610
rect 30970 19558 30976 19610
rect 1104 19536 30976 19558
rect 18414 19456 18420 19508
rect 18472 19456 18478 19508
rect 23661 19499 23719 19505
rect 23661 19465 23673 19499
rect 23707 19496 23719 19499
rect 23707 19468 24808 19496
rect 23707 19465 23719 19468
rect 23661 19459 23719 19465
rect 2130 19388 2136 19440
rect 2188 19388 2194 19440
rect 3878 19388 3884 19440
rect 3936 19388 3942 19440
rect 15194 19428 15200 19440
rect 14844 19400 15200 19428
rect 3234 19320 3240 19372
rect 3292 19320 3298 19372
rect 10594 19320 10600 19372
rect 10652 19360 10658 19372
rect 12894 19360 12900 19372
rect 10652 19332 12900 19360
rect 10652 19320 10658 19332
rect 12894 19320 12900 19332
rect 12952 19320 12958 19372
rect 12986 19320 12992 19372
rect 13044 19360 13050 19372
rect 13153 19363 13211 19369
rect 13153 19360 13165 19363
rect 13044 19332 13165 19360
rect 13044 19320 13050 19332
rect 13153 19329 13165 19332
rect 13199 19329 13211 19363
rect 13153 19323 13211 19329
rect 1854 19252 1860 19304
rect 1912 19252 1918 19304
rect 14844 19301 14872 19400
rect 15194 19388 15200 19400
rect 15252 19388 15258 19440
rect 15378 19388 15384 19440
rect 15436 19388 15442 19440
rect 17586 19388 17592 19440
rect 17644 19428 17650 19440
rect 22002 19428 22008 19440
rect 17644 19400 22008 19428
rect 17644 19388 17650 19400
rect 22002 19388 22008 19400
rect 22060 19388 22066 19440
rect 24397 19431 24455 19437
rect 24397 19397 24409 19431
rect 24443 19428 24455 19431
rect 24670 19428 24676 19440
rect 24443 19400 24676 19428
rect 24443 19397 24455 19400
rect 24397 19391 24455 19397
rect 24670 19388 24676 19400
rect 24728 19388 24734 19440
rect 24780 19428 24808 19468
rect 25866 19456 25872 19508
rect 25924 19496 25930 19508
rect 27430 19496 27436 19508
rect 25924 19468 27436 19496
rect 25924 19456 25930 19468
rect 27430 19456 27436 19468
rect 27488 19496 27494 19508
rect 27801 19499 27859 19505
rect 27801 19496 27813 19499
rect 27488 19468 27813 19496
rect 27488 19456 27494 19468
rect 27801 19465 27813 19468
rect 27847 19465 27859 19499
rect 27801 19459 27859 19465
rect 27893 19499 27951 19505
rect 27893 19465 27905 19499
rect 27939 19496 27951 19499
rect 28626 19496 28632 19508
rect 27939 19468 28632 19496
rect 27939 19465 27951 19468
rect 27893 19459 27951 19465
rect 28626 19456 28632 19468
rect 28684 19456 28690 19508
rect 24780 19400 24886 19428
rect 27982 19388 27988 19440
rect 28040 19388 28046 19440
rect 29914 19428 29920 19440
rect 28920 19400 29920 19428
rect 15105 19363 15163 19369
rect 15105 19329 15117 19363
rect 15151 19360 15163 19363
rect 15396 19360 15424 19388
rect 15151 19332 15424 19360
rect 15151 19329 15163 19332
rect 15105 19323 15163 19329
rect 15654 19320 15660 19372
rect 15712 19360 15718 19372
rect 15749 19363 15807 19369
rect 15749 19360 15761 19363
rect 15712 19332 15761 19360
rect 15712 19320 15718 19332
rect 15749 19329 15761 19332
rect 15795 19329 15807 19363
rect 15749 19323 15807 19329
rect 18506 19320 18512 19372
rect 18564 19320 18570 19372
rect 23477 19363 23535 19369
rect 23477 19329 23489 19363
rect 23523 19360 23535 19363
rect 23566 19360 23572 19372
rect 23523 19332 23572 19360
rect 23523 19329 23535 19332
rect 23477 19323 23535 19329
rect 23566 19320 23572 19332
rect 23624 19320 23630 19372
rect 23658 19320 23664 19372
rect 23716 19360 23722 19372
rect 28920 19369 28948 19400
rect 29914 19388 29920 19400
rect 29972 19388 29978 19440
rect 24121 19363 24179 19369
rect 24121 19360 24133 19363
rect 23716 19332 24133 19360
rect 23716 19320 23722 19332
rect 24121 19329 24133 19332
rect 24167 19329 24179 19363
rect 24121 19323 24179 19329
rect 28905 19363 28963 19369
rect 28905 19329 28917 19363
rect 28951 19329 28963 19363
rect 28905 19323 28963 19329
rect 28994 19320 29000 19372
rect 29052 19320 29058 19372
rect 29178 19320 29184 19372
rect 29236 19320 29242 19372
rect 14829 19295 14887 19301
rect 14829 19261 14841 19295
rect 14875 19261 14887 19295
rect 14829 19255 14887 19261
rect 15381 19295 15439 19301
rect 15381 19261 15393 19295
rect 15427 19261 15439 19295
rect 15381 19255 15439 19261
rect 16117 19295 16175 19301
rect 16117 19261 16129 19295
rect 16163 19292 16175 19295
rect 16206 19292 16212 19304
rect 16163 19264 16212 19292
rect 16163 19261 16175 19264
rect 16117 19255 16175 19261
rect 14458 19184 14464 19236
rect 14516 19224 14522 19236
rect 15286 19224 15292 19236
rect 14516 19196 15292 19224
rect 14516 19184 14522 19196
rect 15286 19184 15292 19196
rect 15344 19224 15350 19236
rect 15396 19224 15424 19255
rect 15344 19196 15424 19224
rect 15344 19184 15350 19196
rect 14274 19116 14280 19168
rect 14332 19156 14338 19168
rect 16132 19156 16160 19255
rect 16206 19252 16212 19264
rect 16264 19252 16270 19304
rect 29362 19252 29368 19304
rect 29420 19252 29426 19304
rect 27617 19227 27675 19233
rect 27617 19193 27629 19227
rect 27663 19224 27675 19227
rect 27706 19224 27712 19236
rect 27663 19196 27712 19224
rect 27663 19193 27675 19196
rect 27617 19187 27675 19193
rect 27706 19184 27712 19196
rect 27764 19184 27770 19236
rect 14332 19128 16160 19156
rect 28169 19159 28227 19165
rect 14332 19116 14338 19128
rect 28169 19125 28181 19159
rect 28215 19156 28227 19159
rect 29178 19156 29184 19168
rect 28215 19128 29184 19156
rect 28215 19125 28227 19128
rect 28169 19119 28227 19125
rect 29178 19116 29184 19128
rect 29236 19116 29242 19168
rect 1104 19066 30820 19088
rect 1104 19014 4664 19066
rect 4716 19014 4728 19066
rect 4780 19014 4792 19066
rect 4844 19014 4856 19066
rect 4908 19014 4920 19066
rect 4972 19014 12092 19066
rect 12144 19014 12156 19066
rect 12208 19014 12220 19066
rect 12272 19014 12284 19066
rect 12336 19014 12348 19066
rect 12400 19014 19520 19066
rect 19572 19014 19584 19066
rect 19636 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 26948 19066
rect 27000 19014 27012 19066
rect 27064 19014 27076 19066
rect 27128 19014 27140 19066
rect 27192 19014 27204 19066
rect 27256 19014 30820 19066
rect 1104 18992 30820 19014
rect 1854 18912 1860 18964
rect 1912 18952 1918 18964
rect 2409 18955 2467 18961
rect 2409 18952 2421 18955
rect 1912 18924 2421 18952
rect 1912 18912 1918 18924
rect 2409 18921 2421 18924
rect 2455 18921 2467 18955
rect 2409 18915 2467 18921
rect 3234 18912 3240 18964
rect 3292 18952 3298 18964
rect 3329 18955 3387 18961
rect 3329 18952 3341 18955
rect 3292 18924 3341 18952
rect 3292 18912 3298 18924
rect 3329 18921 3341 18924
rect 3375 18921 3387 18955
rect 3329 18915 3387 18921
rect 12986 18912 12992 18964
rect 13044 18912 13050 18964
rect 20073 18955 20131 18961
rect 20073 18921 20085 18955
rect 20119 18952 20131 18955
rect 25406 18952 25412 18964
rect 20119 18924 25412 18952
rect 20119 18921 20131 18924
rect 20073 18915 20131 18921
rect 25406 18912 25412 18924
rect 25464 18912 25470 18964
rect 28442 18912 28448 18964
rect 28500 18912 28506 18964
rect 28994 18912 29000 18964
rect 29052 18952 29058 18964
rect 29181 18955 29239 18961
rect 29181 18952 29193 18955
rect 29052 18924 29193 18952
rect 29052 18912 29058 18924
rect 29181 18921 29193 18924
rect 29227 18921 29239 18955
rect 29181 18915 29239 18921
rect 27982 18884 27988 18896
rect 27632 18856 27988 18884
rect 7760 18788 9168 18816
rect 2498 18708 2504 18760
rect 2556 18708 2562 18760
rect 3418 18708 3424 18760
rect 3476 18748 3482 18760
rect 4062 18748 4068 18760
rect 3476 18720 4068 18748
rect 3476 18708 3482 18720
rect 4062 18708 4068 18720
rect 4120 18748 4126 18760
rect 7760 18757 7788 18788
rect 9140 18757 9168 18788
rect 12342 18776 12348 18828
rect 12400 18816 12406 18828
rect 13541 18819 13599 18825
rect 13541 18816 13553 18819
rect 12400 18788 13553 18816
rect 12400 18776 12406 18788
rect 13541 18785 13553 18788
rect 13587 18816 13599 18819
rect 14366 18816 14372 18828
rect 13587 18788 14372 18816
rect 13587 18785 13599 18788
rect 13541 18779 13599 18785
rect 14366 18776 14372 18788
rect 14424 18776 14430 18828
rect 17126 18776 17132 18828
rect 17184 18816 17190 18828
rect 21269 18819 21327 18825
rect 17184 18788 18000 18816
rect 17184 18776 17190 18788
rect 7745 18751 7803 18757
rect 4120 18720 5764 18748
rect 4120 18708 4126 18720
rect 5736 18692 5764 18720
rect 7745 18717 7757 18751
rect 7791 18717 7803 18751
rect 7745 18711 7803 18717
rect 8205 18751 8263 18757
rect 8205 18717 8217 18751
rect 8251 18717 8263 18751
rect 8205 18711 8263 18717
rect 9125 18751 9183 18757
rect 9125 18717 9137 18751
rect 9171 18748 9183 18751
rect 9214 18748 9220 18760
rect 9171 18720 9220 18748
rect 9171 18717 9183 18720
rect 9125 18711 9183 18717
rect 5718 18640 5724 18692
rect 5776 18680 5782 18692
rect 8220 18680 8248 18711
rect 9214 18708 9220 18720
rect 9272 18708 9278 18760
rect 11146 18708 11152 18760
rect 11204 18748 11210 18760
rect 13357 18751 13415 18757
rect 13357 18748 13369 18751
rect 11204 18720 13369 18748
rect 11204 18708 11210 18720
rect 13357 18717 13369 18720
rect 13403 18717 13415 18751
rect 13357 18711 13415 18717
rect 13814 18708 13820 18760
rect 13872 18748 13878 18760
rect 15105 18751 15163 18757
rect 15105 18748 15117 18751
rect 13872 18720 15117 18748
rect 13872 18708 13878 18720
rect 15105 18717 15117 18720
rect 15151 18717 15163 18751
rect 15105 18711 15163 18717
rect 15286 18708 15292 18760
rect 15344 18748 15350 18760
rect 16298 18748 16304 18760
rect 15344 18720 16304 18748
rect 15344 18708 15350 18720
rect 16298 18708 16304 18720
rect 16356 18748 16362 18760
rect 17972 18757 18000 18788
rect 21269 18785 21281 18819
rect 21315 18816 21327 18819
rect 22922 18816 22928 18828
rect 21315 18788 22928 18816
rect 21315 18785 21327 18788
rect 21269 18779 21327 18785
rect 22922 18776 22928 18788
rect 22980 18776 22986 18828
rect 23658 18776 23664 18828
rect 23716 18816 23722 18828
rect 24578 18816 24584 18828
rect 23716 18788 24584 18816
rect 23716 18776 23722 18788
rect 24578 18776 24584 18788
rect 24636 18776 24642 18828
rect 17865 18751 17923 18757
rect 17865 18748 17877 18751
rect 16356 18720 17877 18748
rect 16356 18708 16362 18720
rect 17865 18717 17877 18720
rect 17911 18717 17923 18751
rect 17865 18711 17923 18717
rect 17957 18751 18015 18757
rect 17957 18717 17969 18751
rect 18003 18748 18015 18751
rect 18414 18748 18420 18760
rect 18003 18720 18420 18748
rect 18003 18717 18015 18720
rect 17957 18711 18015 18717
rect 18414 18708 18420 18720
rect 18472 18708 18478 18760
rect 19426 18708 19432 18760
rect 19484 18708 19490 18760
rect 19886 18708 19892 18760
rect 19944 18708 19950 18760
rect 20990 18708 20996 18760
rect 21048 18748 21054 18760
rect 21085 18751 21143 18757
rect 21085 18748 21097 18751
rect 21048 18720 21097 18748
rect 21048 18708 21054 18720
rect 21085 18717 21097 18720
rect 21131 18717 21143 18751
rect 21085 18711 21143 18717
rect 27430 18708 27436 18760
rect 27488 18708 27494 18760
rect 27632 18757 27660 18856
rect 27982 18844 27988 18856
rect 28040 18844 28046 18896
rect 29196 18884 29224 18915
rect 29196 18856 30144 18884
rect 27709 18819 27767 18825
rect 27709 18785 27721 18819
rect 27755 18816 27767 18819
rect 29733 18819 29791 18825
rect 27755 18788 29040 18816
rect 27755 18785 27767 18788
rect 27709 18779 27767 18785
rect 27617 18751 27675 18757
rect 27617 18717 27629 18751
rect 27663 18717 27675 18751
rect 27617 18711 27675 18717
rect 27837 18751 27895 18757
rect 27837 18717 27849 18751
rect 27883 18748 27895 18751
rect 28537 18751 28595 18757
rect 28537 18748 28549 18751
rect 27883 18720 28549 18748
rect 27883 18717 27895 18720
rect 27837 18711 27895 18717
rect 28537 18717 28549 18720
rect 28583 18748 28595 18751
rect 28626 18748 28632 18760
rect 28583 18720 28632 18748
rect 28583 18717 28595 18720
rect 28537 18711 28595 18717
rect 28626 18708 28632 18720
rect 28684 18708 28690 18760
rect 29012 18757 29040 18788
rect 29733 18785 29745 18819
rect 29779 18816 29791 18819
rect 29822 18816 29828 18828
rect 29779 18788 29828 18816
rect 29779 18785 29791 18788
rect 29733 18779 29791 18785
rect 29822 18776 29828 18788
rect 29880 18776 29886 18828
rect 29914 18776 29920 18828
rect 29972 18816 29978 18828
rect 30009 18819 30067 18825
rect 30009 18816 30021 18819
rect 29972 18788 30021 18816
rect 29972 18776 29978 18788
rect 30009 18785 30021 18788
rect 30055 18785 30067 18819
rect 30009 18779 30067 18785
rect 28997 18751 29055 18757
rect 28997 18717 29009 18751
rect 29043 18717 29055 18751
rect 28997 18711 29055 18717
rect 29178 18708 29184 18760
rect 29236 18708 29242 18760
rect 30116 18757 30144 18856
rect 30101 18751 30159 18757
rect 30101 18717 30113 18751
rect 30147 18717 30159 18751
rect 30101 18711 30159 18717
rect 5776 18652 8248 18680
rect 13449 18683 13507 18689
rect 5776 18640 5782 18652
rect 13449 18649 13461 18683
rect 13495 18680 13507 18683
rect 14274 18680 14280 18692
rect 13495 18652 14280 18680
rect 13495 18649 13507 18652
rect 13449 18643 13507 18649
rect 14274 18640 14280 18652
rect 14332 18640 14338 18692
rect 17402 18640 17408 18692
rect 17460 18640 17466 18692
rect 17494 18640 17500 18692
rect 17552 18640 17558 18692
rect 18046 18640 18052 18692
rect 18104 18640 18110 18692
rect 24854 18640 24860 18692
rect 24912 18640 24918 18692
rect 25314 18640 25320 18692
rect 25372 18640 25378 18692
rect 27706 18640 27712 18692
rect 27764 18640 27770 18692
rect 7466 18572 7472 18624
rect 7524 18612 7530 18624
rect 7653 18615 7711 18621
rect 7653 18612 7665 18615
rect 7524 18584 7665 18612
rect 7524 18572 7530 18584
rect 7653 18581 7665 18584
rect 7699 18581 7711 18615
rect 7653 18575 7711 18581
rect 8297 18615 8355 18621
rect 8297 18581 8309 18615
rect 8343 18612 8355 18615
rect 8754 18612 8760 18624
rect 8343 18584 8760 18612
rect 8343 18581 8355 18584
rect 8297 18575 8355 18581
rect 8754 18572 8760 18584
rect 8812 18572 8818 18624
rect 9122 18572 9128 18624
rect 9180 18612 9186 18624
rect 9217 18615 9275 18621
rect 9217 18612 9229 18615
rect 9180 18584 9229 18612
rect 9180 18572 9186 18584
rect 9217 18581 9229 18584
rect 9263 18581 9275 18615
rect 9217 18575 9275 18581
rect 15194 18572 15200 18624
rect 15252 18612 15258 18624
rect 15470 18612 15476 18624
rect 15252 18584 15476 18612
rect 15252 18572 15258 18584
rect 15470 18572 15476 18584
rect 15528 18572 15534 18624
rect 16390 18572 16396 18624
rect 16448 18572 16454 18624
rect 17512 18612 17540 18640
rect 18322 18612 18328 18624
rect 17512 18584 18328 18612
rect 18322 18572 18328 18584
rect 18380 18572 18386 18624
rect 20622 18572 20628 18624
rect 20680 18572 20686 18624
rect 20993 18615 21051 18621
rect 20993 18581 21005 18615
rect 21039 18612 21051 18615
rect 22462 18612 22468 18624
rect 21039 18584 22468 18612
rect 21039 18581 21051 18584
rect 20993 18575 21051 18581
rect 22462 18572 22468 18584
rect 22520 18572 22526 18624
rect 26326 18572 26332 18624
rect 26384 18612 26390 18624
rect 27724 18612 27752 18640
rect 26384 18584 27752 18612
rect 26384 18572 26390 18584
rect 1104 18522 30976 18544
rect 1104 18470 8378 18522
rect 8430 18470 8442 18522
rect 8494 18470 8506 18522
rect 8558 18470 8570 18522
rect 8622 18470 8634 18522
rect 8686 18470 15806 18522
rect 15858 18470 15870 18522
rect 15922 18470 15934 18522
rect 15986 18470 15998 18522
rect 16050 18470 16062 18522
rect 16114 18470 23234 18522
rect 23286 18470 23298 18522
rect 23350 18470 23362 18522
rect 23414 18470 23426 18522
rect 23478 18470 23490 18522
rect 23542 18470 30662 18522
rect 30714 18470 30726 18522
rect 30778 18470 30790 18522
rect 30842 18470 30854 18522
rect 30906 18470 30918 18522
rect 30970 18470 30976 18522
rect 1104 18448 30976 18470
rect 2498 18368 2504 18420
rect 2556 18408 2562 18420
rect 2556 18380 4108 18408
rect 2556 18368 2562 18380
rect 2774 18300 2780 18352
rect 2832 18300 2838 18352
rect 4080 18349 4108 18380
rect 6546 18368 6552 18420
rect 6604 18368 6610 18420
rect 12345 18411 12403 18417
rect 12345 18377 12357 18411
rect 12391 18408 12403 18411
rect 14553 18411 14611 18417
rect 12391 18380 12425 18408
rect 12391 18377 12403 18380
rect 12345 18371 12403 18377
rect 14553 18377 14565 18411
rect 14599 18377 14611 18411
rect 14553 18371 14611 18377
rect 4065 18343 4123 18349
rect 4065 18309 4077 18343
rect 4111 18309 4123 18343
rect 6564 18340 6592 18368
rect 4065 18303 4123 18309
rect 5276 18312 6592 18340
rect 5276 18281 5304 18312
rect 7466 18300 7472 18352
rect 7524 18300 7530 18352
rect 8754 18340 8760 18352
rect 8694 18312 8760 18340
rect 8754 18300 8760 18312
rect 8812 18300 8818 18352
rect 9214 18300 9220 18352
rect 9272 18300 9278 18352
rect 11698 18300 11704 18352
rect 11756 18340 11762 18352
rect 12360 18340 12388 18371
rect 14568 18340 14596 18371
rect 15470 18368 15476 18420
rect 15528 18408 15534 18420
rect 17126 18408 17132 18420
rect 15528 18380 17132 18408
rect 15528 18368 15534 18380
rect 17126 18368 17132 18380
rect 17184 18368 17190 18420
rect 17221 18411 17279 18417
rect 17221 18377 17233 18411
rect 17267 18408 17279 18411
rect 18046 18408 18052 18420
rect 17267 18380 18052 18408
rect 17267 18377 17279 18380
rect 17221 18371 17279 18377
rect 14734 18340 14740 18352
rect 11756 18312 14412 18340
rect 14568 18312 14740 18340
rect 11756 18300 11762 18312
rect 5261 18275 5319 18281
rect 5261 18241 5273 18275
rect 5307 18241 5319 18275
rect 5261 18235 5319 18241
rect 5718 18232 5724 18284
rect 5776 18272 5782 18284
rect 5905 18275 5963 18281
rect 5905 18272 5917 18275
rect 5776 18244 5917 18272
rect 5776 18232 5782 18244
rect 5905 18241 5917 18244
rect 5951 18241 5963 18275
rect 5905 18235 5963 18241
rect 6549 18275 6607 18281
rect 6549 18241 6561 18275
rect 6595 18272 6607 18275
rect 6730 18272 6736 18284
rect 6595 18244 6736 18272
rect 6595 18241 6607 18244
rect 6549 18235 6607 18241
rect 6730 18232 6736 18244
rect 6788 18232 6794 18284
rect 9861 18275 9919 18281
rect 9861 18241 9873 18275
rect 9907 18272 9919 18275
rect 10870 18272 10876 18284
rect 9907 18244 10876 18272
rect 9907 18241 9919 18244
rect 9861 18235 9919 18241
rect 10870 18232 10876 18244
rect 10928 18232 10934 18284
rect 12894 18232 12900 18284
rect 12952 18272 12958 18284
rect 13173 18275 13231 18281
rect 13173 18272 13185 18275
rect 12952 18244 13185 18272
rect 12952 18232 12958 18244
rect 13173 18241 13185 18244
rect 13219 18241 13231 18275
rect 13173 18235 13231 18241
rect 13440 18275 13498 18281
rect 13440 18241 13452 18275
rect 13486 18272 13498 18275
rect 14274 18272 14280 18284
rect 13486 18244 14280 18272
rect 13486 18241 13498 18244
rect 13440 18235 13498 18241
rect 14274 18232 14280 18244
rect 14332 18232 14338 18284
rect 14384 18272 14412 18312
rect 14734 18300 14740 18312
rect 14792 18340 14798 18352
rect 15381 18343 15439 18349
rect 15381 18340 15393 18343
rect 14792 18312 15393 18340
rect 14792 18300 14798 18312
rect 15381 18309 15393 18312
rect 15427 18340 15439 18343
rect 15654 18340 15660 18352
rect 15427 18312 15660 18340
rect 15427 18309 15439 18312
rect 15381 18303 15439 18309
rect 15654 18300 15660 18312
rect 15712 18340 15718 18352
rect 17313 18343 17371 18349
rect 17313 18340 17325 18343
rect 15712 18312 17325 18340
rect 15712 18300 15718 18312
rect 17313 18309 17325 18312
rect 17359 18340 17371 18343
rect 17402 18340 17408 18352
rect 17359 18312 17408 18340
rect 17359 18309 17371 18312
rect 17313 18303 17371 18309
rect 17402 18300 17408 18312
rect 17460 18300 17466 18352
rect 15194 18272 15200 18284
rect 14384 18244 15200 18272
rect 15194 18232 15200 18244
rect 15252 18232 15258 18284
rect 15286 18232 15292 18284
rect 15344 18272 15350 18284
rect 15473 18275 15531 18281
rect 15473 18272 15485 18275
rect 15344 18244 15485 18272
rect 15344 18232 15350 18244
rect 15473 18241 15485 18244
rect 15519 18241 15531 18275
rect 15473 18235 15531 18241
rect 15565 18275 15623 18281
rect 15565 18241 15577 18275
rect 15611 18241 15623 18275
rect 15565 18235 15623 18241
rect 16025 18275 16083 18281
rect 16025 18241 16037 18275
rect 16071 18272 16083 18275
rect 16206 18272 16212 18284
rect 16071 18244 16212 18272
rect 16071 18241 16083 18244
rect 16025 18235 16083 18241
rect 2038 18164 2044 18216
rect 2096 18164 2102 18216
rect 2314 18164 2320 18216
rect 2372 18164 2378 18216
rect 6641 18207 6699 18213
rect 6641 18173 6653 18207
rect 6687 18204 6699 18207
rect 7193 18207 7251 18213
rect 7193 18204 7205 18207
rect 6687 18176 7205 18204
rect 6687 18173 6699 18176
rect 6641 18167 6699 18173
rect 7193 18173 7205 18176
rect 7239 18173 7251 18207
rect 7193 18167 7251 18173
rect 12434 18164 12440 18216
rect 12492 18164 12498 18216
rect 12529 18207 12587 18213
rect 12529 18173 12541 18207
rect 12575 18173 12587 18207
rect 12529 18167 12587 18173
rect 5169 18139 5227 18145
rect 5169 18105 5181 18139
rect 5215 18136 5227 18139
rect 5994 18136 6000 18148
rect 5215 18108 6000 18136
rect 5215 18105 5227 18108
rect 5169 18099 5227 18105
rect 5994 18096 6000 18108
rect 6052 18096 6058 18148
rect 11882 18096 11888 18148
rect 11940 18136 11946 18148
rect 12342 18136 12348 18148
rect 11940 18108 12348 18136
rect 11940 18096 11946 18108
rect 12342 18096 12348 18108
rect 12400 18136 12406 18148
rect 12544 18136 12572 18167
rect 15378 18164 15384 18216
rect 15436 18204 15442 18216
rect 15580 18204 15608 18235
rect 16206 18232 16212 18244
rect 16264 18272 16270 18284
rect 16264 18244 17356 18272
rect 16264 18232 16270 18244
rect 15436 18176 15608 18204
rect 15933 18207 15991 18213
rect 15436 18164 15442 18176
rect 15933 18173 15945 18207
rect 15979 18204 15991 18207
rect 16482 18204 16488 18216
rect 15979 18176 16488 18204
rect 15979 18173 15991 18176
rect 15933 18167 15991 18173
rect 16482 18164 16488 18176
rect 16540 18164 16546 18216
rect 16945 18207 17003 18213
rect 16945 18173 16957 18207
rect 16991 18173 17003 18207
rect 17328 18204 17356 18244
rect 17604 18204 17632 18380
rect 18046 18368 18052 18380
rect 18104 18368 18110 18420
rect 22186 18368 22192 18420
rect 22244 18408 22250 18420
rect 22373 18411 22431 18417
rect 22373 18408 22385 18411
rect 22244 18380 22385 18408
rect 22244 18368 22250 18380
rect 22373 18377 22385 18380
rect 22419 18377 22431 18411
rect 22373 18371 22431 18377
rect 24854 18368 24860 18420
rect 24912 18368 24918 18420
rect 25317 18411 25375 18417
rect 25317 18377 25329 18411
rect 25363 18408 25375 18411
rect 26326 18408 26332 18420
rect 25363 18380 26332 18408
rect 25363 18377 25375 18380
rect 25317 18371 25375 18377
rect 26326 18368 26332 18380
rect 26384 18368 26390 18420
rect 17678 18300 17684 18352
rect 17736 18340 17742 18352
rect 18322 18340 18328 18352
rect 17736 18312 18328 18340
rect 17736 18300 17742 18312
rect 18322 18300 18328 18312
rect 18380 18340 18386 18352
rect 19972 18343 20030 18349
rect 18380 18312 19104 18340
rect 18380 18300 18386 18312
rect 18966 18232 18972 18284
rect 19024 18232 19030 18284
rect 19076 18281 19104 18312
rect 19972 18309 19984 18343
rect 20018 18340 20030 18343
rect 20622 18340 20628 18352
rect 20018 18312 20628 18340
rect 20018 18309 20030 18312
rect 19972 18303 20030 18309
rect 20622 18300 20628 18312
rect 20680 18300 20686 18352
rect 21376 18312 22692 18340
rect 19061 18275 19119 18281
rect 19061 18241 19073 18275
rect 19107 18241 19119 18275
rect 19061 18235 19119 18241
rect 19245 18275 19303 18281
rect 19245 18241 19257 18275
rect 19291 18272 19303 18275
rect 21376 18272 21404 18312
rect 19291 18244 21404 18272
rect 19291 18241 19303 18244
rect 19245 18235 19303 18241
rect 17328 18176 17632 18204
rect 16945 18167 17003 18173
rect 12400 18108 12572 18136
rect 12400 18096 12406 18108
rect 5810 18028 5816 18080
rect 5868 18028 5874 18080
rect 9766 18028 9772 18080
rect 9824 18028 9830 18080
rect 11974 18028 11980 18080
rect 12032 18028 12038 18080
rect 16298 18028 16304 18080
rect 16356 18068 16362 18080
rect 16960 18068 16988 18167
rect 18230 18164 18236 18216
rect 18288 18204 18294 18216
rect 18984 18204 19012 18232
rect 18288 18176 19012 18204
rect 19705 18207 19763 18213
rect 18288 18164 18294 18176
rect 19705 18173 19717 18207
rect 19751 18173 19763 18207
rect 19705 18167 19763 18173
rect 16356 18040 16988 18068
rect 19720 18068 19748 18167
rect 21450 18164 21456 18216
rect 21508 18204 21514 18216
rect 22664 18213 22692 18312
rect 25222 18232 25228 18284
rect 25280 18232 25286 18284
rect 29822 18232 29828 18284
rect 29880 18232 29886 18284
rect 22465 18207 22523 18213
rect 22465 18204 22477 18207
rect 21508 18176 22477 18204
rect 21508 18164 21514 18176
rect 22465 18173 22477 18176
rect 22511 18173 22523 18207
rect 22465 18167 22523 18173
rect 22649 18207 22707 18213
rect 22649 18173 22661 18207
rect 22695 18204 22707 18207
rect 22922 18204 22928 18216
rect 22695 18176 22928 18204
rect 22695 18173 22707 18176
rect 22649 18167 22707 18173
rect 22922 18164 22928 18176
rect 22980 18164 22986 18216
rect 25406 18164 25412 18216
rect 25464 18164 25470 18216
rect 30101 18207 30159 18213
rect 30101 18173 30113 18207
rect 30147 18204 30159 18207
rect 31018 18204 31024 18216
rect 30147 18176 31024 18204
rect 30147 18173 30159 18176
rect 30101 18167 30159 18173
rect 31018 18164 31024 18176
rect 31076 18164 31082 18216
rect 20070 18068 20076 18080
rect 19720 18040 20076 18068
rect 16356 18028 16362 18040
rect 20070 18028 20076 18040
rect 20128 18028 20134 18080
rect 20990 18028 20996 18080
rect 21048 18068 21054 18080
rect 21085 18071 21143 18077
rect 21085 18068 21097 18071
rect 21048 18040 21097 18068
rect 21048 18028 21054 18040
rect 21085 18037 21097 18040
rect 21131 18037 21143 18071
rect 21085 18031 21143 18037
rect 22002 18028 22008 18080
rect 22060 18028 22066 18080
rect 1104 17978 30820 18000
rect 1104 17926 4664 17978
rect 4716 17926 4728 17978
rect 4780 17926 4792 17978
rect 4844 17926 4856 17978
rect 4908 17926 4920 17978
rect 4972 17926 12092 17978
rect 12144 17926 12156 17978
rect 12208 17926 12220 17978
rect 12272 17926 12284 17978
rect 12336 17926 12348 17978
rect 12400 17926 19520 17978
rect 19572 17926 19584 17978
rect 19636 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 26948 17978
rect 27000 17926 27012 17978
rect 27064 17926 27076 17978
rect 27128 17926 27140 17978
rect 27192 17926 27204 17978
rect 27256 17926 30820 17978
rect 1104 17904 30820 17926
rect 2041 17867 2099 17873
rect 2041 17833 2053 17867
rect 2087 17864 2099 17867
rect 2314 17864 2320 17876
rect 2087 17836 2320 17864
rect 2087 17833 2099 17836
rect 2041 17827 2099 17833
rect 2314 17824 2320 17836
rect 2372 17824 2378 17876
rect 2685 17867 2743 17873
rect 2685 17833 2697 17867
rect 2731 17864 2743 17867
rect 2774 17864 2780 17876
rect 2731 17836 2780 17864
rect 2731 17833 2743 17836
rect 2685 17827 2743 17833
rect 2774 17824 2780 17836
rect 2832 17824 2838 17876
rect 11054 17864 11060 17876
rect 8404 17836 11060 17864
rect 8404 17737 8432 17836
rect 11054 17824 11060 17836
rect 11112 17824 11118 17876
rect 12434 17824 12440 17876
rect 12492 17864 12498 17876
rect 13173 17867 13231 17873
rect 13173 17864 13185 17867
rect 12492 17836 13185 17864
rect 12492 17824 12498 17836
rect 13173 17833 13185 17836
rect 13219 17833 13231 17867
rect 13173 17827 13231 17833
rect 10870 17756 10876 17808
rect 10928 17756 10934 17808
rect 8389 17731 8447 17737
rect 8389 17697 8401 17731
rect 8435 17697 8447 17731
rect 8389 17691 8447 17697
rect 9122 17688 9128 17740
rect 9180 17688 9186 17740
rect 9401 17731 9459 17737
rect 9401 17697 9413 17731
rect 9447 17728 9459 17731
rect 9766 17728 9772 17740
rect 9447 17700 9772 17728
rect 9447 17697 9459 17700
rect 9401 17691 9459 17697
rect 9766 17688 9772 17700
rect 9824 17688 9830 17740
rect 11974 17688 11980 17740
rect 12032 17728 12038 17740
rect 12069 17731 12127 17737
rect 12069 17728 12081 17731
rect 12032 17700 12081 17728
rect 12032 17688 12038 17700
rect 12069 17697 12081 17700
rect 12115 17697 12127 17731
rect 12069 17691 12127 17697
rect 2133 17663 2191 17669
rect 2133 17629 2145 17663
rect 2179 17660 2191 17663
rect 2498 17660 2504 17672
rect 2179 17632 2504 17660
rect 2179 17629 2191 17632
rect 2133 17623 2191 17629
rect 2498 17620 2504 17632
rect 2556 17620 2562 17672
rect 2593 17663 2651 17669
rect 2593 17629 2605 17663
rect 2639 17660 2651 17663
rect 3326 17660 3332 17672
rect 2639 17632 3332 17660
rect 2639 17629 2651 17632
rect 2593 17623 2651 17629
rect 3326 17620 3332 17632
rect 3384 17620 3390 17672
rect 3421 17663 3479 17669
rect 3421 17629 3433 17663
rect 3467 17660 3479 17663
rect 3970 17660 3976 17672
rect 3467 17632 3976 17660
rect 3467 17629 3479 17632
rect 3421 17623 3479 17629
rect 3970 17620 3976 17632
rect 4028 17620 4034 17672
rect 5074 17620 5080 17672
rect 5132 17620 5138 17672
rect 5718 17620 5724 17672
rect 5776 17620 5782 17672
rect 5813 17663 5871 17669
rect 5813 17629 5825 17663
rect 5859 17660 5871 17663
rect 6546 17660 6552 17672
rect 5859 17632 6552 17660
rect 5859 17629 5871 17632
rect 5813 17623 5871 17629
rect 6546 17620 6552 17632
rect 6604 17620 6610 17672
rect 11793 17663 11851 17669
rect 11793 17629 11805 17663
rect 11839 17660 11851 17663
rect 12434 17660 12440 17672
rect 11839 17632 12440 17660
rect 11839 17629 11851 17632
rect 11793 17623 11851 17629
rect 12434 17620 12440 17632
rect 12492 17660 12498 17672
rect 12894 17660 12900 17672
rect 12492 17632 12900 17660
rect 12492 17620 12498 17632
rect 12894 17620 12900 17632
rect 12952 17620 12958 17672
rect 13188 17660 13216 17827
rect 14274 17824 14280 17876
rect 14332 17824 14338 17876
rect 21450 17824 21456 17876
rect 21508 17824 21514 17876
rect 14366 17756 14372 17808
rect 14424 17796 14430 17808
rect 14424 17768 14872 17796
rect 14424 17756 14430 17768
rect 14734 17688 14740 17740
rect 14792 17688 14798 17740
rect 14844 17737 14872 17768
rect 14829 17731 14887 17737
rect 14829 17697 14841 17731
rect 14875 17697 14887 17731
rect 14829 17691 14887 17697
rect 16298 17688 16304 17740
rect 16356 17728 16362 17740
rect 16356 17700 18552 17728
rect 16356 17688 16362 17700
rect 15194 17660 15200 17672
rect 13188 17632 15200 17660
rect 15194 17620 15200 17632
rect 15252 17620 15258 17672
rect 15654 17620 15660 17672
rect 15712 17660 15718 17672
rect 16390 17660 16396 17672
rect 15712 17632 16396 17660
rect 15712 17620 15718 17632
rect 16390 17620 16396 17632
rect 16448 17620 16454 17672
rect 17957 17663 18015 17669
rect 17957 17660 17969 17663
rect 17236 17632 17969 17660
rect 6365 17595 6423 17601
rect 6365 17561 6377 17595
rect 6411 17592 6423 17595
rect 6730 17592 6736 17604
rect 6411 17564 6736 17592
rect 6411 17561 6423 17564
rect 6365 17555 6423 17561
rect 6730 17552 6736 17564
rect 6788 17552 6794 17604
rect 7466 17552 7472 17604
rect 7524 17552 7530 17604
rect 8113 17595 8171 17601
rect 8113 17561 8125 17595
rect 8159 17561 8171 17595
rect 10962 17592 10968 17604
rect 10626 17564 10968 17592
rect 8113 17555 8171 17561
rect 3326 17484 3332 17536
rect 3384 17484 3390 17536
rect 6822 17484 6828 17536
rect 6880 17524 6886 17536
rect 8128 17524 8156 17555
rect 10962 17552 10968 17564
rect 11020 17552 11026 17604
rect 14645 17595 14703 17601
rect 14645 17561 14657 17595
rect 14691 17592 14703 17595
rect 15102 17592 15108 17604
rect 14691 17564 15108 17592
rect 14691 17561 14703 17564
rect 14645 17555 14703 17561
rect 15102 17552 15108 17564
rect 15160 17552 15166 17604
rect 15470 17552 15476 17604
rect 15528 17592 15534 17604
rect 17236 17592 17264 17632
rect 17957 17629 17969 17632
rect 18003 17629 18015 17663
rect 17957 17623 18015 17629
rect 18414 17620 18420 17672
rect 18472 17620 18478 17672
rect 18524 17669 18552 17700
rect 20070 17688 20076 17740
rect 20128 17688 20134 17740
rect 18509 17663 18567 17669
rect 18509 17629 18521 17663
rect 18555 17629 18567 17663
rect 18509 17623 18567 17629
rect 15528 17564 17264 17592
rect 17405 17595 17463 17601
rect 15528 17552 15534 17564
rect 17405 17561 17417 17595
rect 17451 17592 17463 17595
rect 17862 17592 17868 17604
rect 17451 17564 17868 17592
rect 17451 17561 17463 17564
rect 17405 17555 17463 17561
rect 17862 17552 17868 17564
rect 17920 17552 17926 17604
rect 18049 17595 18107 17601
rect 18049 17561 18061 17595
rect 18095 17561 18107 17595
rect 18049 17555 18107 17561
rect 6880 17496 8156 17524
rect 6880 17484 6886 17496
rect 17954 17484 17960 17536
rect 18012 17524 18018 17536
rect 18064 17524 18092 17555
rect 18138 17552 18144 17604
rect 18196 17592 18202 17604
rect 18601 17595 18659 17601
rect 18601 17592 18613 17595
rect 18196 17564 18613 17592
rect 18196 17552 18202 17564
rect 18601 17561 18613 17564
rect 18647 17561 18659 17595
rect 20088 17592 20116 17688
rect 20340 17663 20398 17669
rect 20340 17629 20352 17663
rect 20386 17660 20398 17663
rect 22002 17660 22008 17672
rect 20386 17632 22008 17660
rect 20386 17629 20398 17632
rect 20340 17623 20398 17629
rect 22002 17620 22008 17632
rect 22060 17620 22066 17672
rect 22189 17663 22247 17669
rect 22189 17629 22201 17663
rect 22235 17660 22247 17663
rect 22235 17632 22692 17660
rect 22235 17629 22247 17632
rect 22189 17623 22247 17629
rect 22204 17592 22232 17623
rect 22462 17601 22468 17604
rect 20088 17564 22232 17592
rect 18601 17555 18659 17561
rect 22456 17555 22468 17601
rect 22462 17552 22468 17555
rect 22520 17552 22526 17604
rect 22664 17592 22692 17632
rect 22738 17620 22744 17672
rect 22796 17660 22802 17672
rect 25222 17660 25228 17672
rect 22796 17632 25228 17660
rect 22796 17620 22802 17632
rect 25222 17620 25228 17632
rect 25280 17620 25286 17672
rect 26605 17663 26663 17669
rect 26605 17629 26617 17663
rect 26651 17660 26663 17663
rect 27614 17660 27620 17672
rect 26651 17632 27620 17660
rect 26651 17629 26663 17632
rect 26605 17623 26663 17629
rect 27614 17620 27620 17632
rect 27672 17620 27678 17672
rect 23658 17592 23664 17604
rect 22664 17564 23664 17592
rect 23658 17552 23664 17564
rect 23716 17552 23722 17604
rect 18012 17496 18092 17524
rect 18012 17484 18018 17496
rect 23566 17484 23572 17536
rect 23624 17484 23630 17536
rect 26418 17484 26424 17536
rect 26476 17524 26482 17536
rect 26513 17527 26571 17533
rect 26513 17524 26525 17527
rect 26476 17496 26525 17524
rect 26476 17484 26482 17496
rect 26513 17493 26525 17496
rect 26559 17493 26571 17527
rect 26513 17487 26571 17493
rect 1104 17434 30976 17456
rect 1104 17382 8378 17434
rect 8430 17382 8442 17434
rect 8494 17382 8506 17434
rect 8558 17382 8570 17434
rect 8622 17382 8634 17434
rect 8686 17382 15806 17434
rect 15858 17382 15870 17434
rect 15922 17382 15934 17434
rect 15986 17382 15998 17434
rect 16050 17382 16062 17434
rect 16114 17382 23234 17434
rect 23286 17382 23298 17434
rect 23350 17382 23362 17434
rect 23414 17382 23426 17434
rect 23478 17382 23490 17434
rect 23542 17382 30662 17434
rect 30714 17382 30726 17434
rect 30778 17382 30790 17434
rect 30842 17382 30854 17434
rect 30906 17382 30918 17434
rect 30970 17382 30976 17434
rect 1104 17360 30976 17382
rect 5718 17280 5724 17332
rect 5776 17320 5782 17332
rect 5776 17292 5948 17320
rect 5776 17280 5782 17292
rect 3970 17212 3976 17264
rect 4028 17212 4034 17264
rect 5810 17252 5816 17264
rect 5290 17224 5816 17252
rect 5810 17212 5816 17224
rect 5868 17212 5874 17264
rect 5920 17252 5948 17292
rect 6822 17280 6828 17332
rect 6880 17280 6886 17332
rect 7466 17280 7472 17332
rect 7524 17280 7530 17332
rect 13814 17320 13820 17332
rect 13648 17292 13820 17320
rect 12434 17252 12440 17264
rect 5920 17224 7420 17252
rect 2866 17144 2872 17196
rect 2924 17144 2930 17196
rect 3329 17187 3387 17193
rect 3329 17153 3341 17187
rect 3375 17184 3387 17187
rect 3418 17184 3424 17196
rect 3375 17156 3424 17184
rect 3375 17153 3387 17156
rect 3329 17147 3387 17153
rect 3418 17144 3424 17156
rect 3476 17144 3482 17196
rect 5994 17144 6000 17196
rect 6052 17144 6058 17196
rect 6730 17144 6736 17196
rect 6788 17144 6794 17196
rect 7392 17193 7420 17224
rect 11716 17224 12440 17252
rect 11716 17193 11744 17224
rect 12434 17212 12440 17224
rect 12492 17212 12498 17264
rect 13648 17261 13676 17292
rect 13814 17280 13820 17292
rect 13872 17320 13878 17332
rect 14642 17320 14648 17332
rect 13872 17292 14648 17320
rect 13872 17280 13878 17292
rect 14642 17280 14648 17292
rect 14700 17280 14706 17332
rect 16758 17280 16764 17332
rect 16816 17320 16822 17332
rect 17770 17320 17776 17332
rect 16816 17292 17776 17320
rect 16816 17280 16822 17292
rect 17770 17280 17776 17292
rect 17828 17320 17834 17332
rect 19426 17320 19432 17332
rect 17828 17292 19432 17320
rect 17828 17280 17834 17292
rect 13633 17255 13691 17261
rect 13633 17221 13645 17255
rect 13679 17221 13691 17255
rect 13633 17215 13691 17221
rect 13998 17212 14004 17264
rect 14056 17212 14062 17264
rect 14185 17255 14243 17261
rect 14185 17221 14197 17255
rect 14231 17252 14243 17255
rect 15286 17252 15292 17264
rect 14231 17224 15292 17252
rect 14231 17221 14243 17224
rect 14185 17215 14243 17221
rect 15286 17212 15292 17224
rect 15344 17212 15350 17264
rect 15378 17212 15384 17264
rect 15436 17252 15442 17264
rect 15436 17224 15976 17252
rect 15436 17212 15442 17224
rect 7377 17187 7435 17193
rect 7377 17153 7389 17187
rect 7423 17153 7435 17187
rect 7377 17147 7435 17153
rect 11701 17187 11759 17193
rect 11701 17153 11713 17187
rect 11747 17153 11759 17187
rect 11701 17147 11759 17153
rect 11790 17144 11796 17196
rect 11848 17184 11854 17196
rect 11957 17187 12015 17193
rect 11957 17184 11969 17187
rect 11848 17156 11969 17184
rect 11848 17144 11854 17156
rect 11957 17153 11969 17156
rect 12003 17153 12015 17187
rect 11957 17147 12015 17153
rect 14093 17187 14151 17193
rect 14093 17153 14105 17187
rect 14139 17153 14151 17187
rect 14093 17147 14151 17153
rect 5718 17076 5724 17128
rect 5776 17076 5782 17128
rect 13078 17008 13084 17060
rect 13136 17048 13142 17060
rect 14108 17048 14136 17147
rect 15194 17144 15200 17196
rect 15252 17144 15258 17196
rect 15470 17144 15476 17196
rect 15528 17144 15534 17196
rect 15948 17193 15976 17224
rect 16206 17212 16212 17264
rect 16264 17252 16270 17264
rect 18138 17252 18144 17264
rect 16264 17224 18144 17252
rect 16264 17212 16270 17224
rect 18138 17212 18144 17224
rect 18196 17252 18202 17264
rect 18196 17224 18552 17252
rect 18196 17212 18202 17224
rect 15933 17187 15991 17193
rect 15933 17153 15945 17187
rect 15979 17184 15991 17187
rect 16114 17184 16120 17196
rect 15979 17156 16120 17184
rect 15979 17153 15991 17156
rect 15933 17147 15991 17153
rect 16114 17144 16120 17156
rect 16172 17144 16178 17196
rect 16758 17144 16764 17196
rect 16816 17184 16822 17196
rect 16853 17187 16911 17193
rect 16853 17184 16865 17187
rect 16816 17156 16865 17184
rect 16816 17144 16822 17156
rect 16853 17153 16865 17156
rect 16899 17153 16911 17187
rect 16853 17147 16911 17153
rect 17494 17144 17500 17196
rect 17552 17144 17558 17196
rect 18230 17144 18236 17196
rect 18288 17144 18294 17196
rect 18322 17144 18328 17196
rect 18380 17144 18386 17196
rect 18417 17187 18475 17193
rect 18417 17153 18429 17187
rect 18463 17153 18475 17187
rect 18524 17184 18552 17224
rect 19352 17193 19380 17292
rect 19426 17280 19432 17292
rect 19484 17280 19490 17332
rect 22373 17323 22431 17329
rect 22373 17289 22385 17323
rect 22419 17320 22431 17323
rect 22462 17320 22468 17332
rect 22419 17292 22468 17320
rect 22419 17289 22431 17292
rect 22373 17283 22431 17289
rect 22462 17280 22468 17292
rect 22520 17280 22526 17332
rect 27614 17320 27620 17332
rect 26206 17292 27620 17320
rect 26206 17252 26234 17292
rect 27614 17280 27620 17292
rect 27672 17280 27678 17332
rect 20916 17224 26234 17252
rect 20916 17193 20944 17224
rect 27430 17212 27436 17264
rect 27488 17212 27494 17264
rect 18601 17187 18659 17193
rect 18601 17184 18613 17187
rect 18524 17156 18613 17184
rect 18417 17147 18475 17153
rect 18601 17153 18613 17156
rect 18647 17153 18659 17187
rect 18601 17147 18659 17153
rect 19061 17187 19119 17193
rect 19061 17153 19073 17187
rect 19107 17153 19119 17187
rect 19061 17147 19119 17153
rect 19337 17187 19395 17193
rect 19337 17153 19349 17187
rect 19383 17153 19395 17187
rect 19337 17147 19395 17153
rect 20901 17187 20959 17193
rect 20901 17153 20913 17187
rect 20947 17153 20959 17187
rect 20901 17147 20959 17153
rect 14274 17076 14280 17128
rect 14332 17116 14338 17128
rect 14369 17119 14427 17125
rect 14369 17116 14381 17119
rect 14332 17088 14381 17116
rect 14332 17076 14338 17088
rect 14369 17085 14381 17088
rect 14415 17085 14427 17119
rect 15488 17116 15516 17144
rect 14369 17079 14427 17085
rect 14476 17088 15516 17116
rect 14476 17048 14504 17088
rect 15746 17076 15752 17128
rect 15804 17116 15810 17128
rect 16298 17116 16304 17128
rect 15804 17088 16304 17116
rect 15804 17076 15810 17088
rect 16298 17076 16304 17088
rect 16356 17076 16362 17128
rect 16574 17076 16580 17128
rect 16632 17116 16638 17128
rect 17221 17119 17279 17125
rect 17221 17116 17233 17119
rect 16632 17088 17233 17116
rect 16632 17076 16638 17088
rect 17221 17085 17233 17088
rect 17267 17085 17279 17119
rect 17221 17079 17279 17085
rect 13136 17020 14504 17048
rect 13136 17008 13142 17020
rect 15378 17008 15384 17060
rect 15436 17048 15442 17060
rect 15562 17048 15568 17060
rect 15436 17020 15568 17048
rect 15436 17008 15442 17020
rect 15562 17008 15568 17020
rect 15620 17048 15626 17060
rect 18248 17048 18276 17144
rect 18432 17116 18460 17147
rect 19076 17116 19104 17147
rect 22738 17144 22744 17196
rect 22796 17144 22802 17196
rect 22833 17187 22891 17193
rect 22833 17153 22845 17187
rect 22879 17184 22891 17187
rect 23566 17184 23572 17196
rect 22879 17156 23572 17184
rect 22879 17153 22891 17156
rect 22833 17147 22891 17153
rect 23566 17144 23572 17156
rect 23624 17184 23630 17196
rect 23845 17187 23903 17193
rect 23624 17156 23796 17184
rect 23624 17144 23630 17156
rect 18432 17088 19104 17116
rect 18432 17060 18460 17088
rect 19426 17076 19432 17128
rect 19484 17076 19490 17128
rect 20990 17076 20996 17128
rect 21048 17076 21054 17128
rect 22922 17076 22928 17128
rect 22980 17076 22986 17128
rect 23768 17125 23796 17156
rect 23845 17153 23857 17187
rect 23891 17184 23903 17187
rect 26053 17187 26111 17193
rect 26053 17184 26065 17187
rect 23891 17156 26065 17184
rect 23891 17153 23903 17156
rect 23845 17147 23903 17153
rect 26053 17153 26065 17156
rect 26099 17184 26111 17187
rect 28350 17184 28356 17196
rect 26099 17156 26234 17184
rect 28106 17156 28356 17184
rect 26099 17153 26111 17156
rect 26053 17147 26111 17153
rect 23753 17119 23811 17125
rect 23753 17085 23765 17119
rect 23799 17085 23811 17119
rect 26206 17116 26234 17156
rect 28350 17144 28356 17156
rect 28408 17184 28414 17196
rect 28408 17156 28934 17184
rect 28408 17144 28414 17156
rect 27890 17116 27896 17128
rect 26206 17088 27896 17116
rect 23753 17079 23811 17085
rect 27890 17076 27896 17088
rect 27948 17076 27954 17128
rect 27982 17076 27988 17128
rect 28040 17116 28046 17128
rect 28997 17119 29055 17125
rect 28997 17116 29009 17119
rect 28040 17088 29009 17116
rect 28040 17076 28046 17088
rect 28997 17085 29009 17088
rect 29043 17085 29055 17119
rect 28997 17079 29055 17085
rect 29730 17076 29736 17128
rect 29788 17076 29794 17128
rect 15620 17020 18276 17048
rect 15620 17008 15626 17020
rect 18414 17008 18420 17060
rect 18472 17008 18478 17060
rect 2777 16983 2835 16989
rect 2777 16949 2789 16983
rect 2823 16980 2835 16983
rect 2958 16980 2964 16992
rect 2823 16952 2964 16980
rect 2823 16949 2835 16952
rect 2777 16943 2835 16949
rect 2958 16940 2964 16952
rect 3016 16940 3022 16992
rect 3418 16940 3424 16992
rect 3476 16940 3482 16992
rect 14274 16940 14280 16992
rect 14332 16980 14338 16992
rect 15746 16980 15752 16992
rect 14332 16952 15752 16980
rect 14332 16940 14338 16952
rect 15746 16940 15752 16952
rect 15804 16940 15810 16992
rect 18046 16940 18052 16992
rect 18104 16940 18110 16992
rect 21266 16940 21272 16992
rect 21324 16940 21330 16992
rect 24213 16983 24271 16989
rect 24213 16949 24225 16983
rect 24259 16980 24271 16983
rect 24946 16980 24952 16992
rect 24259 16952 24952 16980
rect 24259 16949 24271 16952
rect 24213 16943 24271 16949
rect 24946 16940 24952 16952
rect 25004 16940 25010 16992
rect 26142 16940 26148 16992
rect 26200 16940 26206 16992
rect 1104 16890 30820 16912
rect 1104 16838 4664 16890
rect 4716 16838 4728 16890
rect 4780 16838 4792 16890
rect 4844 16838 4856 16890
rect 4908 16838 4920 16890
rect 4972 16838 12092 16890
rect 12144 16838 12156 16890
rect 12208 16838 12220 16890
rect 12272 16838 12284 16890
rect 12336 16838 12348 16890
rect 12400 16838 19520 16890
rect 19572 16838 19584 16890
rect 19636 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 26948 16890
rect 27000 16838 27012 16890
rect 27064 16838 27076 16890
rect 27128 16838 27140 16890
rect 27192 16838 27204 16890
rect 27256 16838 30820 16890
rect 1104 16816 30820 16838
rect 11790 16736 11796 16788
rect 11848 16736 11854 16788
rect 11882 16736 11888 16788
rect 11940 16776 11946 16788
rect 12342 16776 12348 16788
rect 11940 16748 12348 16776
rect 11940 16736 11946 16748
rect 12342 16736 12348 16748
rect 12400 16736 12406 16788
rect 14366 16736 14372 16788
rect 14424 16736 14430 16788
rect 18414 16776 18420 16788
rect 16868 16748 18420 16776
rect 2866 16668 2872 16720
rect 2924 16708 2930 16720
rect 4706 16708 4712 16720
rect 2924 16680 4712 16708
rect 2924 16668 2930 16680
rect 4706 16668 4712 16680
rect 4764 16668 4770 16720
rect 9784 16680 13400 16708
rect 2884 16640 2912 16668
rect 2792 16612 2912 16640
rect 2038 16532 2044 16584
rect 2096 16572 2102 16584
rect 2792 16581 2820 16612
rect 3970 16600 3976 16652
rect 4028 16640 4034 16652
rect 4028 16612 4568 16640
rect 4028 16600 4034 16612
rect 4540 16581 4568 16612
rect 9582 16600 9588 16652
rect 9640 16640 9646 16652
rect 9784 16649 9812 16680
rect 9769 16643 9827 16649
rect 9769 16640 9781 16643
rect 9640 16612 9781 16640
rect 9640 16600 9646 16612
rect 9769 16609 9781 16612
rect 9815 16609 9827 16643
rect 9769 16603 9827 16609
rect 12253 16643 12311 16649
rect 12253 16609 12265 16643
rect 12299 16609 12311 16643
rect 12253 16603 12311 16609
rect 2685 16575 2743 16581
rect 2685 16572 2697 16575
rect 2096 16544 2697 16572
rect 2096 16532 2102 16544
rect 2685 16541 2697 16544
rect 2731 16541 2743 16575
rect 2685 16535 2743 16541
rect 2777 16575 2835 16581
rect 2777 16541 2789 16575
rect 2823 16541 2835 16575
rect 2777 16535 2835 16541
rect 4525 16575 4583 16581
rect 4525 16541 4537 16575
rect 4571 16541 4583 16575
rect 4525 16535 4583 16541
rect 4617 16575 4675 16581
rect 4617 16541 4629 16575
rect 4663 16572 4675 16575
rect 5718 16572 5724 16584
rect 4663 16544 5724 16572
rect 4663 16541 4675 16544
rect 4617 16535 4675 16541
rect 5718 16532 5724 16544
rect 5776 16532 5782 16584
rect 6178 16532 6184 16584
rect 6236 16532 6242 16584
rect 12268 16572 12296 16603
rect 12342 16600 12348 16652
rect 12400 16600 12406 16652
rect 13078 16640 13084 16652
rect 12452 16612 13084 16640
rect 12452 16572 12480 16612
rect 13078 16600 13084 16612
rect 13136 16600 13142 16652
rect 13372 16649 13400 16680
rect 15562 16668 15568 16720
rect 15620 16708 15626 16720
rect 16482 16708 16488 16720
rect 15620 16680 16488 16708
rect 15620 16668 15626 16680
rect 16482 16668 16488 16680
rect 16540 16708 16546 16720
rect 16868 16708 16896 16748
rect 18414 16736 18420 16748
rect 18472 16736 18478 16788
rect 27614 16736 27620 16788
rect 27672 16776 27678 16788
rect 27893 16779 27951 16785
rect 27893 16776 27905 16779
rect 27672 16748 27905 16776
rect 27672 16736 27678 16748
rect 27893 16745 27905 16748
rect 27939 16745 27951 16779
rect 27893 16739 27951 16745
rect 16540 16680 16896 16708
rect 16540 16668 16546 16680
rect 13357 16643 13415 16649
rect 13357 16609 13369 16643
rect 13403 16609 13415 16643
rect 13814 16640 13820 16652
rect 13357 16603 13415 16609
rect 13740 16612 13820 16640
rect 12268 16544 12480 16572
rect 13538 16532 13544 16584
rect 13596 16532 13602 16584
rect 13740 16581 13768 16612
rect 13814 16600 13820 16612
rect 13872 16600 13878 16652
rect 14274 16600 14280 16652
rect 14332 16640 14338 16652
rect 14461 16643 14519 16649
rect 14461 16640 14473 16643
rect 14332 16612 14473 16640
rect 14332 16600 14338 16612
rect 14461 16609 14473 16612
rect 14507 16640 14519 16643
rect 14507 16612 15148 16640
rect 14507 16609 14519 16612
rect 14461 16603 14519 16609
rect 13725 16575 13783 16581
rect 13725 16541 13737 16575
rect 13771 16572 13783 16575
rect 14737 16575 14795 16581
rect 13771 16544 13805 16572
rect 13771 16541 13783 16544
rect 13725 16535 13783 16541
rect 14737 16541 14749 16575
rect 14783 16541 14795 16575
rect 14737 16535 14795 16541
rect 6454 16464 6460 16516
rect 6512 16464 6518 16516
rect 8294 16464 8300 16516
rect 8352 16504 8358 16516
rect 9585 16507 9643 16513
rect 9585 16504 9597 16507
rect 8352 16476 9597 16504
rect 8352 16464 8358 16476
rect 9585 16473 9597 16476
rect 9631 16473 9643 16507
rect 9585 16467 9643 16473
rect 9122 16396 9128 16448
rect 9180 16396 9186 16448
rect 9490 16396 9496 16448
rect 9548 16436 9554 16448
rect 12161 16439 12219 16445
rect 12161 16436 12173 16439
rect 9548 16408 12173 16436
rect 9548 16396 9554 16408
rect 12161 16405 12173 16408
rect 12207 16405 12219 16439
rect 14752 16436 14780 16535
rect 15120 16504 15148 16612
rect 15194 16600 15200 16652
rect 15252 16640 15258 16652
rect 16301 16643 16359 16649
rect 15252 16612 15976 16640
rect 15252 16600 15258 16612
rect 15470 16532 15476 16584
rect 15528 16572 15534 16584
rect 15841 16575 15899 16581
rect 15841 16572 15853 16575
rect 15528 16544 15853 16572
rect 15528 16532 15534 16544
rect 15841 16541 15853 16544
rect 15887 16541 15899 16575
rect 15841 16535 15899 16541
rect 15948 16513 15976 16612
rect 16301 16609 16313 16643
rect 16347 16640 16359 16643
rect 16758 16640 16764 16652
rect 16347 16612 16764 16640
rect 16347 16609 16359 16612
rect 16301 16603 16359 16609
rect 16758 16600 16764 16612
rect 16816 16600 16822 16652
rect 16868 16581 16896 16680
rect 17034 16668 17040 16720
rect 17092 16668 17098 16720
rect 17954 16708 17960 16720
rect 17144 16680 17960 16708
rect 17144 16581 17172 16680
rect 17954 16668 17960 16680
rect 18012 16668 18018 16720
rect 19426 16600 19432 16652
rect 19484 16640 19490 16652
rect 19978 16640 19984 16652
rect 19484 16612 19984 16640
rect 19484 16600 19490 16612
rect 19978 16600 19984 16612
rect 20036 16600 20042 16652
rect 26142 16600 26148 16652
rect 26200 16600 26206 16652
rect 26418 16600 26424 16652
rect 26476 16600 26482 16652
rect 16853 16575 16911 16581
rect 16853 16541 16865 16575
rect 16899 16541 16911 16575
rect 16853 16535 16911 16541
rect 17129 16575 17187 16581
rect 17129 16541 17141 16575
rect 17175 16541 17187 16575
rect 17129 16535 17187 16541
rect 17589 16575 17647 16581
rect 17589 16541 17601 16575
rect 17635 16541 17647 16575
rect 17589 16535 17647 16541
rect 15565 16507 15623 16513
rect 15565 16504 15577 16507
rect 15120 16476 15577 16504
rect 15565 16473 15577 16476
rect 15611 16473 15623 16507
rect 15565 16467 15623 16473
rect 15933 16507 15991 16513
rect 15933 16473 15945 16507
rect 15979 16504 15991 16507
rect 16206 16504 16212 16516
rect 15979 16476 16212 16504
rect 15979 16473 15991 16476
rect 15933 16467 15991 16473
rect 16206 16464 16212 16476
rect 16264 16464 16270 16516
rect 16482 16464 16488 16516
rect 16540 16504 16546 16516
rect 17604 16504 17632 16535
rect 17862 16532 17868 16584
rect 17920 16532 17926 16584
rect 18009 16575 18067 16581
rect 18009 16541 18021 16575
rect 18055 16572 18067 16575
rect 22002 16572 22008 16584
rect 18055 16544 22008 16572
rect 18055 16541 18067 16544
rect 18009 16535 18067 16541
rect 22002 16532 22008 16544
rect 22060 16532 22066 16584
rect 27890 16532 27896 16584
rect 27948 16572 27954 16584
rect 28258 16572 28264 16584
rect 27948 16544 28264 16572
rect 27948 16532 27954 16544
rect 28258 16532 28264 16544
rect 28316 16572 28322 16584
rect 28537 16575 28595 16581
rect 28537 16572 28549 16575
rect 28316 16544 28549 16572
rect 28316 16532 28322 16544
rect 28537 16541 28549 16544
rect 28583 16541 28595 16575
rect 28537 16535 28595 16541
rect 29638 16532 29644 16584
rect 29696 16572 29702 16584
rect 29733 16575 29791 16581
rect 29733 16572 29745 16575
rect 29696 16544 29745 16572
rect 29696 16532 29702 16544
rect 29733 16541 29745 16544
rect 29779 16541 29791 16575
rect 29733 16535 29791 16541
rect 16540 16476 17632 16504
rect 17773 16507 17831 16513
rect 16540 16464 16546 16476
rect 17773 16473 17785 16507
rect 17819 16504 17831 16507
rect 18158 16507 18216 16513
rect 17819 16476 18092 16504
rect 17819 16473 17831 16476
rect 17773 16467 17831 16473
rect 18064 16448 18092 16476
rect 18158 16473 18170 16507
rect 18204 16504 18216 16507
rect 23106 16504 23112 16516
rect 18204 16476 23112 16504
rect 18204 16473 18216 16476
rect 18158 16467 18216 16473
rect 23106 16464 23112 16476
rect 23164 16464 23170 16516
rect 27430 16464 27436 16516
rect 27488 16464 27494 16516
rect 15286 16436 15292 16448
rect 14752 16408 15292 16436
rect 12161 16399 12219 16405
rect 15286 16396 15292 16408
rect 15344 16436 15350 16448
rect 15749 16439 15807 16445
rect 15749 16436 15761 16439
rect 15344 16408 15761 16436
rect 15344 16396 15350 16408
rect 15749 16405 15761 16408
rect 15795 16436 15807 16439
rect 16114 16436 16120 16448
rect 15795 16408 16120 16436
rect 15795 16405 15807 16408
rect 15749 16399 15807 16405
rect 16114 16396 16120 16408
rect 16172 16396 16178 16448
rect 18046 16396 18052 16448
rect 18104 16396 18110 16448
rect 19426 16396 19432 16448
rect 19484 16396 19490 16448
rect 19518 16396 19524 16448
rect 19576 16436 19582 16448
rect 19797 16439 19855 16445
rect 19797 16436 19809 16439
rect 19576 16408 19809 16436
rect 19576 16396 19582 16408
rect 19797 16405 19809 16408
rect 19843 16405 19855 16439
rect 19797 16399 19855 16405
rect 19886 16396 19892 16448
rect 19944 16396 19950 16448
rect 28629 16439 28687 16445
rect 28629 16405 28641 16439
rect 28675 16436 28687 16439
rect 28718 16436 28724 16448
rect 28675 16408 28724 16436
rect 28675 16405 28687 16408
rect 28629 16399 28687 16405
rect 28718 16396 28724 16408
rect 28776 16396 28782 16448
rect 29825 16439 29883 16445
rect 29825 16405 29837 16439
rect 29871 16436 29883 16439
rect 30006 16436 30012 16448
rect 29871 16408 30012 16436
rect 29871 16405 29883 16408
rect 29825 16399 29883 16405
rect 30006 16396 30012 16408
rect 30064 16396 30070 16448
rect 1104 16346 30976 16368
rect 1104 16294 8378 16346
rect 8430 16294 8442 16346
rect 8494 16294 8506 16346
rect 8558 16294 8570 16346
rect 8622 16294 8634 16346
rect 8686 16294 15806 16346
rect 15858 16294 15870 16346
rect 15922 16294 15934 16346
rect 15986 16294 15998 16346
rect 16050 16294 16062 16346
rect 16114 16294 23234 16346
rect 23286 16294 23298 16346
rect 23350 16294 23362 16346
rect 23414 16294 23426 16346
rect 23478 16294 23490 16346
rect 23542 16294 30662 16346
rect 30714 16294 30726 16346
rect 30778 16294 30790 16346
rect 30842 16294 30854 16346
rect 30906 16294 30918 16346
rect 30970 16294 30976 16346
rect 1104 16272 30976 16294
rect 7469 16235 7527 16241
rect 7469 16201 7481 16235
rect 7515 16232 7527 16235
rect 7515 16204 10916 16232
rect 7515 16201 7527 16204
rect 7469 16195 7527 16201
rect 2958 16124 2964 16176
rect 3016 16124 3022 16176
rect 3418 16124 3424 16176
rect 3476 16124 3482 16176
rect 4706 16124 4712 16176
rect 4764 16124 4770 16176
rect 9122 16124 9128 16176
rect 9180 16164 9186 16176
rect 9410 16167 9468 16173
rect 9410 16164 9422 16167
rect 9180 16136 9422 16164
rect 9180 16124 9186 16136
rect 9410 16133 9422 16136
rect 9456 16133 9468 16167
rect 10888 16164 10916 16204
rect 10962 16192 10968 16244
rect 11020 16192 11026 16244
rect 13538 16192 13544 16244
rect 13596 16232 13602 16244
rect 15562 16232 15568 16244
rect 13596 16204 15568 16232
rect 13596 16192 13602 16204
rect 15562 16192 15568 16204
rect 15620 16192 15626 16244
rect 28258 16192 28264 16244
rect 28316 16192 28322 16244
rect 11146 16164 11152 16176
rect 10888 16136 11152 16164
rect 9410 16127 9468 16133
rect 11146 16124 11152 16136
rect 11204 16124 11210 16176
rect 14737 16167 14795 16173
rect 14737 16133 14749 16167
rect 14783 16164 14795 16167
rect 15654 16164 15660 16176
rect 14783 16136 15660 16164
rect 14783 16133 14795 16136
rect 14737 16127 14795 16133
rect 15654 16124 15660 16136
rect 15712 16124 15718 16176
rect 18684 16167 18742 16173
rect 18684 16133 18696 16167
rect 18730 16164 18742 16167
rect 19426 16164 19432 16176
rect 18730 16136 19432 16164
rect 18730 16133 18742 16136
rect 18684 16127 18742 16133
rect 19426 16124 19432 16136
rect 19484 16124 19490 16176
rect 29730 16164 29736 16176
rect 29302 16136 29736 16164
rect 29730 16124 29736 16136
rect 29788 16124 29794 16176
rect 9582 16096 9588 16108
rect 7760 16068 9588 16096
rect 2685 16031 2743 16037
rect 2685 15997 2697 16031
rect 2731 16028 2743 16031
rect 3326 16028 3332 16040
rect 2731 16000 3332 16028
rect 2731 15997 2743 16000
rect 2685 15991 2743 15997
rect 3326 15988 3332 16000
rect 3384 15988 3390 16040
rect 6178 15988 6184 16040
rect 6236 16028 6242 16040
rect 7760 16037 7788 16068
rect 9582 16056 9588 16068
rect 9640 16056 9646 16108
rect 10137 16099 10195 16105
rect 10137 16096 10149 16099
rect 9692 16068 10149 16096
rect 9692 16037 9720 16068
rect 10137 16065 10149 16068
rect 10183 16096 10195 16099
rect 10873 16099 10931 16105
rect 10873 16096 10885 16099
rect 10183 16068 10885 16096
rect 10183 16065 10195 16068
rect 10137 16059 10195 16065
rect 10873 16065 10885 16068
rect 10919 16065 10931 16099
rect 10873 16059 10931 16065
rect 7561 16031 7619 16037
rect 7561 16028 7573 16031
rect 6236 16000 7573 16028
rect 6236 15988 6242 16000
rect 7561 15997 7573 16000
rect 7607 15997 7619 16031
rect 7561 15991 7619 15997
rect 7745 16031 7803 16037
rect 7745 15997 7757 16031
rect 7791 15997 7803 16031
rect 7745 15991 7803 15997
rect 9677 16031 9735 16037
rect 9677 15997 9689 16031
rect 9723 15997 9735 16031
rect 10888 16028 10916 16059
rect 11606 16056 11612 16108
rect 11664 16096 11670 16108
rect 12161 16099 12219 16105
rect 12161 16096 12173 16099
rect 11664 16068 12173 16096
rect 11664 16056 11670 16068
rect 12161 16065 12173 16068
rect 12207 16096 12219 16099
rect 12989 16099 13047 16105
rect 12989 16096 13001 16099
rect 12207 16068 13001 16096
rect 12207 16065 12219 16068
rect 12161 16059 12219 16065
rect 12989 16065 13001 16068
rect 13035 16065 13047 16099
rect 12989 16059 13047 16065
rect 15378 16056 15384 16108
rect 15436 16056 15442 16108
rect 15562 16056 15568 16108
rect 15620 16056 15626 16108
rect 16206 16056 16212 16108
rect 16264 16056 16270 16108
rect 23750 16056 23756 16108
rect 23808 16056 23814 16108
rect 24394 16056 24400 16108
rect 24452 16096 24458 16108
rect 24581 16099 24639 16105
rect 24581 16096 24593 16099
rect 24452 16068 24593 16096
rect 24452 16056 24458 16068
rect 24581 16065 24593 16068
rect 24627 16096 24639 16099
rect 24762 16096 24768 16108
rect 24627 16068 24768 16096
rect 24627 16065 24639 16068
rect 24581 16059 24639 16065
rect 24762 16056 24768 16068
rect 24820 16056 24826 16108
rect 30006 16056 30012 16108
rect 30064 16056 30070 16108
rect 11790 16028 11796 16040
rect 10888 16000 11796 16028
rect 9677 15991 9735 15997
rect 7101 15895 7159 15901
rect 7101 15861 7113 15895
rect 7147 15892 7159 15895
rect 7282 15892 7288 15904
rect 7147 15864 7288 15892
rect 7147 15861 7159 15864
rect 7101 15855 7159 15861
rect 7282 15852 7288 15864
rect 7340 15852 7346 15904
rect 8294 15852 8300 15904
rect 8352 15852 8358 15904
rect 9306 15852 9312 15904
rect 9364 15892 9370 15904
rect 9692 15892 9720 15991
rect 11790 15988 11796 16000
rect 11848 15988 11854 16040
rect 15102 15988 15108 16040
rect 15160 16028 15166 16040
rect 15197 16031 15255 16037
rect 15197 16028 15209 16031
rect 15160 16000 15209 16028
rect 15160 15988 15166 16000
rect 15197 15997 15209 16000
rect 15243 15997 15255 16031
rect 15197 15991 15255 15997
rect 16482 15988 16488 16040
rect 16540 16028 16546 16040
rect 18417 16031 18475 16037
rect 18417 16028 18429 16031
rect 16540 16000 18429 16028
rect 16540 15988 16546 16000
rect 18417 15997 18429 16000
rect 18463 15997 18475 16031
rect 18417 15991 18475 15997
rect 23569 16031 23627 16037
rect 23569 15997 23581 16031
rect 23615 16028 23627 16031
rect 23658 16028 23664 16040
rect 23615 16000 23664 16028
rect 23615 15997 23627 16000
rect 23569 15991 23627 15997
rect 23658 15988 23664 16000
rect 23716 15988 23722 16040
rect 24302 15988 24308 16040
rect 24360 15988 24366 16040
rect 24489 16031 24547 16037
rect 24489 15997 24501 16031
rect 24535 16028 24547 16031
rect 25958 16028 25964 16040
rect 24535 16000 25964 16028
rect 24535 15997 24547 16000
rect 24489 15991 24547 15997
rect 25958 15988 25964 16000
rect 26016 15988 26022 16040
rect 28718 15988 28724 16040
rect 28776 16028 28782 16040
rect 29733 16031 29791 16037
rect 29733 16028 29745 16031
rect 28776 16000 29745 16028
rect 28776 15988 28782 16000
rect 29733 15997 29745 16000
rect 29779 15997 29791 16031
rect 29733 15991 29791 15997
rect 10321 15963 10379 15969
rect 10321 15929 10333 15963
rect 10367 15960 10379 15963
rect 10367 15932 13768 15960
rect 10367 15929 10379 15932
rect 10321 15923 10379 15929
rect 9364 15864 9720 15892
rect 9364 15852 9370 15864
rect 11882 15852 11888 15904
rect 11940 15892 11946 15904
rect 12069 15895 12127 15901
rect 12069 15892 12081 15895
rect 11940 15864 12081 15892
rect 11940 15852 11946 15864
rect 12069 15861 12081 15864
rect 12115 15861 12127 15895
rect 13740 15892 13768 15932
rect 13814 15920 13820 15972
rect 13872 15960 13878 15972
rect 13998 15960 14004 15972
rect 13872 15932 14004 15960
rect 13872 15920 13878 15932
rect 13998 15920 14004 15932
rect 14056 15960 14062 15972
rect 16117 15963 16175 15969
rect 16117 15960 16129 15963
rect 14056 15932 16129 15960
rect 14056 15920 14062 15932
rect 16117 15929 16129 15932
rect 16163 15929 16175 15963
rect 16117 15923 16175 15929
rect 14090 15892 14096 15904
rect 13740 15864 14096 15892
rect 12069 15855 12127 15861
rect 14090 15852 14096 15864
rect 14148 15852 14154 15904
rect 19797 15895 19855 15901
rect 19797 15861 19809 15895
rect 19843 15892 19855 15895
rect 19886 15892 19892 15904
rect 19843 15864 19892 15892
rect 19843 15861 19855 15864
rect 19797 15855 19855 15861
rect 19886 15852 19892 15864
rect 19944 15852 19950 15904
rect 24854 15852 24860 15904
rect 24912 15892 24918 15904
rect 24949 15895 25007 15901
rect 24949 15892 24961 15895
rect 24912 15864 24961 15892
rect 24912 15852 24918 15864
rect 24949 15861 24961 15864
rect 24995 15861 25007 15895
rect 24949 15855 25007 15861
rect 1104 15802 30820 15824
rect 1104 15750 4664 15802
rect 4716 15750 4728 15802
rect 4780 15750 4792 15802
rect 4844 15750 4856 15802
rect 4908 15750 4920 15802
rect 4972 15750 12092 15802
rect 12144 15750 12156 15802
rect 12208 15750 12220 15802
rect 12272 15750 12284 15802
rect 12336 15750 12348 15802
rect 12400 15750 19520 15802
rect 19572 15750 19584 15802
rect 19636 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 26948 15802
rect 27000 15750 27012 15802
rect 27064 15750 27076 15802
rect 27128 15750 27140 15802
rect 27192 15750 27204 15802
rect 27256 15750 30820 15802
rect 1104 15728 30820 15750
rect 6178 15648 6184 15700
rect 6236 15648 6242 15700
rect 6454 15648 6460 15700
rect 6512 15688 6518 15700
rect 6822 15688 6828 15700
rect 6512 15660 6828 15688
rect 6512 15648 6518 15660
rect 6822 15648 6828 15660
rect 6880 15688 6886 15700
rect 9122 15688 9128 15700
rect 6880 15660 9128 15688
rect 6880 15648 6886 15660
rect 7576 15561 7604 15660
rect 9122 15648 9128 15660
rect 9180 15688 9186 15700
rect 9306 15688 9312 15700
rect 9180 15660 9312 15688
rect 9180 15648 9186 15660
rect 9306 15648 9312 15660
rect 9364 15648 9370 15700
rect 25958 15648 25964 15700
rect 26016 15648 26022 15700
rect 11146 15580 11152 15632
rect 11204 15620 11210 15632
rect 12618 15620 12624 15632
rect 11204 15592 12624 15620
rect 11204 15580 11210 15592
rect 12618 15580 12624 15592
rect 12676 15580 12682 15632
rect 15378 15620 15384 15632
rect 13280 15592 15384 15620
rect 7561 15555 7619 15561
rect 7561 15521 7573 15555
rect 7607 15521 7619 15555
rect 12710 15552 12716 15564
rect 7561 15515 7619 15521
rect 12406 15524 12716 15552
rect 5166 15444 5172 15496
rect 5224 15484 5230 15496
rect 5261 15487 5319 15493
rect 5261 15484 5273 15487
rect 5224 15456 5273 15484
rect 5224 15444 5230 15456
rect 5261 15453 5273 15456
rect 5307 15453 5319 15487
rect 5261 15447 5319 15453
rect 7282 15444 7288 15496
rect 7340 15493 7346 15496
rect 7340 15484 7352 15493
rect 7340 15456 7385 15484
rect 7340 15447 7352 15456
rect 7340 15444 7346 15447
rect 9030 15444 9036 15496
rect 9088 15484 9094 15496
rect 9309 15487 9367 15493
rect 9309 15484 9321 15487
rect 9088 15456 9321 15484
rect 9088 15444 9094 15456
rect 9309 15453 9321 15456
rect 9355 15484 9367 15487
rect 12406 15484 12434 15524
rect 12710 15512 12716 15524
rect 12768 15512 12774 15564
rect 12802 15512 12808 15564
rect 12860 15552 12866 15564
rect 13280 15561 13308 15592
rect 15378 15580 15384 15592
rect 15436 15620 15442 15632
rect 16574 15620 16580 15632
rect 15436 15592 16580 15620
rect 15436 15580 15442 15592
rect 16574 15580 16580 15592
rect 16632 15580 16638 15632
rect 19978 15580 19984 15632
rect 20036 15620 20042 15632
rect 24302 15620 24308 15632
rect 20036 15592 24308 15620
rect 20036 15580 20042 15592
rect 23860 15561 23888 15592
rect 24302 15580 24308 15592
rect 24360 15580 24366 15632
rect 13265 15555 13323 15561
rect 13265 15552 13277 15555
rect 12860 15524 13277 15552
rect 12860 15512 12866 15524
rect 13265 15521 13277 15524
rect 13311 15521 13323 15555
rect 23845 15555 23903 15561
rect 13265 15515 13323 15521
rect 21468 15524 22140 15552
rect 21468 15496 21496 15524
rect 9355 15456 12434 15484
rect 12529 15487 12587 15493
rect 9355 15453 9367 15456
rect 9309 15447 9367 15453
rect 12529 15453 12541 15487
rect 12575 15453 12587 15487
rect 12529 15447 12587 15453
rect 9576 15419 9634 15425
rect 9576 15385 9588 15419
rect 9622 15416 9634 15419
rect 9766 15416 9772 15428
rect 9622 15388 9772 15416
rect 9622 15385 9634 15388
rect 9576 15379 9634 15385
rect 9766 15376 9772 15388
rect 9824 15376 9830 15428
rect 11974 15376 11980 15428
rect 12032 15416 12038 15428
rect 12253 15419 12311 15425
rect 12253 15416 12265 15419
rect 12032 15388 12265 15416
rect 12032 15376 12038 15388
rect 12253 15385 12265 15388
rect 12299 15385 12311 15419
rect 12544 15416 12572 15447
rect 13538 15444 13544 15496
rect 13596 15484 13602 15496
rect 13725 15487 13783 15493
rect 13725 15484 13737 15487
rect 13596 15456 13737 15484
rect 13596 15444 13602 15456
rect 13725 15453 13737 15456
rect 13771 15453 13783 15487
rect 13725 15447 13783 15453
rect 16206 15444 16212 15496
rect 16264 15484 16270 15496
rect 16482 15484 16488 15496
rect 16264 15456 16488 15484
rect 16264 15444 16270 15456
rect 16482 15444 16488 15456
rect 16540 15484 16546 15496
rect 16577 15487 16635 15493
rect 16577 15484 16589 15487
rect 16540 15456 16589 15484
rect 16540 15444 16546 15456
rect 16577 15453 16589 15456
rect 16623 15453 16635 15487
rect 16577 15447 16635 15453
rect 18598 15444 18604 15496
rect 18656 15484 18662 15496
rect 19429 15487 19487 15493
rect 19429 15484 19441 15487
rect 18656 15456 19441 15484
rect 18656 15444 18662 15456
rect 19429 15453 19441 15456
rect 19475 15453 19487 15487
rect 19429 15447 19487 15453
rect 19613 15487 19671 15493
rect 19613 15453 19625 15487
rect 19659 15453 19671 15487
rect 19613 15447 19671 15453
rect 13446 15416 13452 15428
rect 12544 15388 13452 15416
rect 12253 15379 12311 15385
rect 13446 15376 13452 15388
rect 13504 15376 13510 15428
rect 13633 15419 13691 15425
rect 13633 15385 13645 15419
rect 13679 15416 13691 15419
rect 13814 15416 13820 15428
rect 13679 15388 13820 15416
rect 13679 15385 13691 15388
rect 13633 15379 13691 15385
rect 13814 15376 13820 15388
rect 13872 15376 13878 15428
rect 16850 15425 16856 15428
rect 16844 15379 16856 15425
rect 16850 15376 16856 15379
rect 16908 15376 16914 15428
rect 18782 15376 18788 15428
rect 18840 15416 18846 15428
rect 19628 15416 19656 15447
rect 21450 15444 21456 15496
rect 21508 15444 21514 15496
rect 22112 15493 22140 15524
rect 23845 15521 23857 15555
rect 23891 15521 23903 15555
rect 29638 15552 29644 15564
rect 23845 15515 23903 15521
rect 27448 15524 29644 15552
rect 21913 15487 21971 15493
rect 21913 15453 21925 15487
rect 21959 15453 21971 15487
rect 21913 15447 21971 15453
rect 22097 15487 22155 15493
rect 22097 15453 22109 15487
rect 22143 15453 22155 15487
rect 22097 15447 22155 15453
rect 18840 15388 19656 15416
rect 21269 15419 21327 15425
rect 18840 15376 18846 15388
rect 21269 15385 21281 15419
rect 21315 15416 21327 15419
rect 21928 15416 21956 15447
rect 22738 15444 22744 15496
rect 22796 15484 22802 15496
rect 23661 15487 23719 15493
rect 23661 15484 23673 15487
rect 22796 15456 23673 15484
rect 22796 15444 22802 15456
rect 23661 15453 23673 15456
rect 23707 15453 23719 15487
rect 23661 15447 23719 15453
rect 23750 15444 23756 15496
rect 23808 15484 23814 15496
rect 24854 15493 24860 15496
rect 24581 15487 24639 15493
rect 24581 15484 24593 15487
rect 23808 15456 24593 15484
rect 23808 15444 23814 15456
rect 24581 15453 24593 15456
rect 24627 15453 24639 15487
rect 24848 15484 24860 15493
rect 24815 15456 24860 15484
rect 24581 15447 24639 15453
rect 24848 15447 24860 15456
rect 24854 15444 24860 15447
rect 24912 15444 24918 15496
rect 27448 15493 27476 15524
rect 29638 15512 29644 15524
rect 29696 15512 29702 15564
rect 27433 15487 27491 15493
rect 27433 15484 27445 15487
rect 26206 15456 27445 15484
rect 26206 15416 26234 15456
rect 27433 15453 27445 15456
rect 27479 15453 27491 15487
rect 27433 15447 27491 15453
rect 27982 15444 27988 15496
rect 28040 15484 28046 15496
rect 28169 15487 28227 15493
rect 28169 15484 28181 15487
rect 28040 15456 28181 15484
rect 28040 15444 28046 15456
rect 28169 15453 28181 15456
rect 28215 15453 28227 15487
rect 28169 15447 28227 15453
rect 28350 15444 28356 15496
rect 28408 15444 28414 15496
rect 21315 15388 26234 15416
rect 21315 15385 21327 15388
rect 21269 15379 21327 15385
rect 29178 15376 29184 15428
rect 29236 15376 29242 15428
rect 4430 15308 4436 15360
rect 4488 15348 4494 15360
rect 5169 15351 5227 15357
rect 5169 15348 5181 15351
rect 4488 15320 5181 15348
rect 4488 15308 4494 15320
rect 5169 15317 5181 15320
rect 5215 15317 5227 15351
rect 5169 15311 5227 15317
rect 10226 15308 10232 15360
rect 10284 15348 10290 15360
rect 10689 15351 10747 15357
rect 10689 15348 10701 15351
rect 10284 15320 10701 15348
rect 10284 15308 10290 15320
rect 10689 15317 10701 15320
rect 10735 15317 10747 15351
rect 10689 15311 10747 15317
rect 12434 15308 12440 15360
rect 12492 15348 12498 15360
rect 13541 15351 13599 15357
rect 13541 15348 13553 15351
rect 12492 15320 13553 15348
rect 12492 15308 12498 15320
rect 13541 15317 13553 15320
rect 13587 15317 13599 15351
rect 13541 15311 13599 15317
rect 17957 15351 18015 15357
rect 17957 15317 17969 15351
rect 18003 15348 18015 15351
rect 18598 15348 18604 15360
rect 18003 15320 18604 15348
rect 18003 15317 18015 15320
rect 17957 15311 18015 15317
rect 18598 15308 18604 15320
rect 18656 15308 18662 15360
rect 19613 15351 19671 15357
rect 19613 15317 19625 15351
rect 19659 15348 19671 15351
rect 20714 15348 20720 15360
rect 19659 15320 20720 15348
rect 19659 15317 19671 15320
rect 19613 15311 19671 15317
rect 20714 15308 20720 15320
rect 20772 15308 20778 15360
rect 21082 15308 21088 15360
rect 21140 15308 21146 15360
rect 21174 15308 21180 15360
rect 21232 15348 21238 15360
rect 21913 15351 21971 15357
rect 21913 15348 21925 15351
rect 21232 15320 21925 15348
rect 21232 15308 21238 15320
rect 21913 15317 21925 15320
rect 21959 15317 21971 15351
rect 21913 15311 21971 15317
rect 23293 15351 23351 15357
rect 23293 15317 23305 15351
rect 23339 15348 23351 15351
rect 23566 15348 23572 15360
rect 23339 15320 23572 15348
rect 23339 15317 23351 15320
rect 23293 15311 23351 15317
rect 23566 15308 23572 15320
rect 23624 15308 23630 15360
rect 23753 15351 23811 15357
rect 23753 15317 23765 15351
rect 23799 15348 23811 15351
rect 24578 15348 24584 15360
rect 23799 15320 24584 15348
rect 23799 15317 23811 15320
rect 23753 15311 23811 15317
rect 24578 15308 24584 15320
rect 24636 15308 24642 15360
rect 27525 15351 27583 15357
rect 27525 15317 27537 15351
rect 27571 15348 27583 15351
rect 28166 15348 28172 15360
rect 27571 15320 28172 15348
rect 27571 15317 27583 15320
rect 27525 15311 27583 15317
rect 28166 15308 28172 15320
rect 28224 15308 28230 15360
rect 1104 15258 30976 15280
rect 1104 15206 8378 15258
rect 8430 15206 8442 15258
rect 8494 15206 8506 15258
rect 8558 15206 8570 15258
rect 8622 15206 8634 15258
rect 8686 15206 15806 15258
rect 15858 15206 15870 15258
rect 15922 15206 15934 15258
rect 15986 15206 15998 15258
rect 16050 15206 16062 15258
rect 16114 15206 23234 15258
rect 23286 15206 23298 15258
rect 23350 15206 23362 15258
rect 23414 15206 23426 15258
rect 23478 15206 23490 15258
rect 23542 15206 30662 15258
rect 30714 15206 30726 15258
rect 30778 15206 30790 15258
rect 30842 15206 30854 15258
rect 30906 15206 30918 15258
rect 30970 15206 30976 15258
rect 1104 15184 30976 15206
rect 8018 15104 8024 15156
rect 8076 15104 8082 15156
rect 9766 15104 9772 15156
rect 9824 15104 9830 15156
rect 10226 15104 10232 15156
rect 10284 15104 10290 15156
rect 11054 15104 11060 15156
rect 11112 15104 11118 15156
rect 11974 15104 11980 15156
rect 12032 15104 12038 15156
rect 16850 15104 16856 15156
rect 16908 15104 16914 15156
rect 22002 15104 22008 15156
rect 22060 15144 22066 15156
rect 22097 15147 22155 15153
rect 22097 15144 22109 15147
rect 22060 15116 22109 15144
rect 22060 15104 22066 15116
rect 22097 15113 22109 15116
rect 22143 15113 22155 15147
rect 22097 15107 22155 15113
rect 24578 15104 24584 15156
rect 24636 15104 24642 15156
rect 29638 15104 29644 15156
rect 29696 15104 29702 15156
rect 11992 15076 12020 15104
rect 11164 15048 12020 15076
rect 5258 14968 5264 15020
rect 5316 14968 5322 15020
rect 6546 14968 6552 15020
rect 6604 14968 6610 15020
rect 11164 15017 11192 15048
rect 13170 15036 13176 15088
rect 13228 15036 13234 15088
rect 14734 15036 14740 15088
rect 14792 15076 14798 15088
rect 15013 15079 15071 15085
rect 15013 15076 15025 15079
rect 14792 15048 15025 15076
rect 14792 15036 14798 15048
rect 15013 15045 15025 15048
rect 15059 15076 15071 15079
rect 17126 15076 17132 15088
rect 15059 15048 17132 15076
rect 15059 15045 15071 15048
rect 15013 15039 15071 15045
rect 17126 15036 17132 15048
rect 17184 15036 17190 15088
rect 17313 15079 17371 15085
rect 17313 15045 17325 15079
rect 17359 15076 17371 15079
rect 18598 15076 18604 15088
rect 17359 15048 18604 15076
rect 17359 15045 17371 15048
rect 17313 15039 17371 15045
rect 18598 15036 18604 15048
rect 18656 15036 18662 15088
rect 18969 15079 19027 15085
rect 18969 15045 18981 15079
rect 19015 15076 19027 15079
rect 19015 15048 20576 15076
rect 19015 15045 19027 15048
rect 18969 15039 19027 15045
rect 10137 15011 10195 15017
rect 10137 14977 10149 15011
rect 10183 15008 10195 15011
rect 11149 15011 11207 15017
rect 10183 14980 11100 15008
rect 10183 14977 10195 14980
rect 10137 14971 10195 14977
rect 5350 14900 5356 14952
rect 5408 14900 5414 14952
rect 5902 14900 5908 14952
rect 5960 14900 5966 14952
rect 9582 14900 9588 14952
rect 9640 14940 9646 14952
rect 10321 14943 10379 14949
rect 10321 14940 10333 14943
rect 9640 14912 10333 14940
rect 9640 14900 9646 14912
rect 10321 14909 10333 14912
rect 10367 14909 10379 14943
rect 10321 14903 10379 14909
rect 11072 14804 11100 14980
rect 11149 14977 11161 15011
rect 11195 14977 11207 15011
rect 11149 14971 11207 14977
rect 11882 14968 11888 15020
rect 11940 14968 11946 15020
rect 13446 14968 13452 15020
rect 13504 15008 13510 15020
rect 13504 14980 13952 15008
rect 13504 14968 13510 14980
rect 12161 14943 12219 14949
rect 12161 14909 12173 14943
rect 12207 14940 12219 14943
rect 13814 14940 13820 14952
rect 12207 14912 13820 14940
rect 12207 14909 12219 14912
rect 12161 14903 12219 14909
rect 13814 14900 13820 14912
rect 13872 14900 13878 14952
rect 13924 14949 13952 14980
rect 17218 14968 17224 15020
rect 17276 15008 17282 15020
rect 17494 15008 17500 15020
rect 17276 14980 17500 15008
rect 17276 14968 17282 14980
rect 17494 14968 17500 14980
rect 17552 14968 17558 15020
rect 18782 15008 18788 15020
rect 18616 14980 18788 15008
rect 18616 14952 18644 14980
rect 18782 14968 18788 14980
rect 18840 14968 18846 15020
rect 20548 15017 20576 15048
rect 20714 15036 20720 15088
rect 20772 15036 20778 15088
rect 20809 15079 20867 15085
rect 20809 15045 20821 15079
rect 20855 15076 20867 15079
rect 21082 15076 21088 15088
rect 20855 15048 21088 15076
rect 20855 15045 20867 15048
rect 20809 15039 20867 15045
rect 21082 15036 21088 15048
rect 21140 15036 21146 15088
rect 23468 15079 23526 15085
rect 23468 15045 23480 15079
rect 23514 15076 23526 15079
rect 23566 15076 23572 15088
rect 23514 15048 23572 15076
rect 23514 15045 23526 15048
rect 23468 15039 23526 15045
rect 23566 15036 23572 15048
rect 23624 15036 23630 15088
rect 23658 15036 23664 15088
rect 23716 15036 23722 15088
rect 28166 15036 28172 15088
rect 28224 15036 28230 15088
rect 29178 15036 29184 15088
rect 29236 15036 29242 15088
rect 19613 15011 19671 15017
rect 19613 14977 19625 15011
rect 19659 14977 19671 15011
rect 20441 15011 20499 15017
rect 20441 15008 20453 15011
rect 19613 14971 19671 14977
rect 19996 14980 20453 15008
rect 13909 14943 13967 14949
rect 13909 14909 13921 14943
rect 13955 14940 13967 14943
rect 15194 14940 15200 14952
rect 13955 14912 15200 14940
rect 13955 14909 13967 14912
rect 13909 14903 13967 14909
rect 15194 14900 15200 14912
rect 15252 14900 15258 14952
rect 17034 14900 17040 14952
rect 17092 14940 17098 14952
rect 17402 14940 17408 14952
rect 17092 14912 17408 14940
rect 17092 14900 17098 14912
rect 17402 14900 17408 14912
rect 17460 14900 17466 14952
rect 18598 14900 18604 14952
rect 18656 14900 18662 14952
rect 19628 14872 19656 14971
rect 19705 14943 19763 14949
rect 19705 14909 19717 14943
rect 19751 14940 19763 14943
rect 19886 14940 19892 14952
rect 19751 14912 19892 14940
rect 19751 14909 19763 14912
rect 19705 14903 19763 14909
rect 19886 14900 19892 14912
rect 19944 14900 19950 14952
rect 19996 14949 20024 14980
rect 20441 14977 20453 14980
rect 20487 14977 20499 15011
rect 20441 14971 20499 14977
rect 20534 15011 20592 15017
rect 20534 14977 20546 15011
rect 20580 14977 20592 15011
rect 20534 14971 20592 14977
rect 20947 15011 21005 15017
rect 20947 14977 20959 15011
rect 20993 15008 21005 15011
rect 21174 15008 21180 15020
rect 20993 14980 21180 15008
rect 20993 14977 21005 14980
rect 20947 14971 21005 14977
rect 21174 14968 21180 14980
rect 21232 14968 21238 15020
rect 21910 14968 21916 15020
rect 21968 15008 21974 15020
rect 22005 15011 22063 15017
rect 22005 15008 22017 15011
rect 21968 14980 22017 15008
rect 21968 14968 21974 14980
rect 22005 14977 22017 14980
rect 22051 14977 22063 15011
rect 22005 14971 22063 14977
rect 22281 15011 22339 15017
rect 22281 14977 22293 15011
rect 22327 14977 22339 15011
rect 22281 14971 22339 14977
rect 23201 15011 23259 15017
rect 23201 14977 23213 15011
rect 23247 15008 23259 15011
rect 23676 15008 23704 15036
rect 23247 14980 23704 15008
rect 25317 15011 25375 15017
rect 23247 14977 23259 14980
rect 23201 14971 23259 14977
rect 25317 14977 25329 15011
rect 25363 15008 25375 15011
rect 27798 15008 27804 15020
rect 25363 14980 27804 15008
rect 25363 14977 25375 14980
rect 25317 14971 25375 14977
rect 19981 14943 20039 14949
rect 19981 14909 19993 14943
rect 20027 14909 20039 14943
rect 22296 14940 22324 14971
rect 27798 14968 27804 14980
rect 27856 14968 27862 15020
rect 19981 14903 20039 14909
rect 21100 14912 22324 14940
rect 20990 14872 20996 14884
rect 14844 14844 16574 14872
rect 19628 14844 20996 14872
rect 11698 14804 11704 14816
rect 11072 14776 11704 14804
rect 11698 14764 11704 14776
rect 11756 14804 11762 14816
rect 14642 14804 14648 14816
rect 11756 14776 14648 14804
rect 11756 14764 11762 14776
rect 14642 14764 14648 14776
rect 14700 14804 14706 14816
rect 14844 14804 14872 14844
rect 14700 14776 14872 14804
rect 14700 14764 14706 14776
rect 14918 14764 14924 14816
rect 14976 14804 14982 14816
rect 15289 14807 15347 14813
rect 15289 14804 15301 14807
rect 14976 14776 15301 14804
rect 14976 14764 14982 14776
rect 15289 14773 15301 14776
rect 15335 14804 15347 14807
rect 16206 14804 16212 14816
rect 15335 14776 16212 14804
rect 15335 14773 15347 14776
rect 15289 14767 15347 14773
rect 16206 14764 16212 14776
rect 16264 14764 16270 14816
rect 16546 14804 16574 14844
rect 20990 14832 20996 14844
rect 21048 14832 21054 14884
rect 21100 14881 21128 14912
rect 22462 14900 22468 14952
rect 22520 14900 22526 14952
rect 25409 14943 25467 14949
rect 25409 14909 25421 14943
rect 25455 14940 25467 14943
rect 25958 14940 25964 14952
rect 25455 14912 25964 14940
rect 25455 14909 25467 14912
rect 25409 14903 25467 14909
rect 25958 14900 25964 14912
rect 26016 14900 26022 14952
rect 27890 14900 27896 14952
rect 27948 14900 27954 14952
rect 21085 14875 21143 14881
rect 21085 14841 21097 14875
rect 21131 14841 21143 14875
rect 21085 14835 21143 14841
rect 17218 14804 17224 14816
rect 16546 14776 17224 14804
rect 17218 14764 17224 14776
rect 17276 14804 17282 14816
rect 22738 14804 22744 14816
rect 17276 14776 22744 14804
rect 17276 14764 17282 14776
rect 22738 14764 22744 14776
rect 22796 14764 22802 14816
rect 25685 14807 25743 14813
rect 25685 14773 25697 14807
rect 25731 14804 25743 14807
rect 25866 14804 25872 14816
rect 25731 14776 25872 14804
rect 25731 14773 25743 14776
rect 25685 14767 25743 14773
rect 25866 14764 25872 14776
rect 25924 14764 25930 14816
rect 1104 14714 30820 14736
rect 1104 14662 4664 14714
rect 4716 14662 4728 14714
rect 4780 14662 4792 14714
rect 4844 14662 4856 14714
rect 4908 14662 4920 14714
rect 4972 14662 12092 14714
rect 12144 14662 12156 14714
rect 12208 14662 12220 14714
rect 12272 14662 12284 14714
rect 12336 14662 12348 14714
rect 12400 14662 19520 14714
rect 19572 14662 19584 14714
rect 19636 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 26948 14714
rect 27000 14662 27012 14714
rect 27064 14662 27076 14714
rect 27128 14662 27140 14714
rect 27192 14662 27204 14714
rect 27256 14662 30820 14714
rect 1104 14640 30820 14662
rect 6546 14560 6552 14612
rect 6604 14600 6610 14612
rect 18506 14600 18512 14612
rect 6604 14572 18512 14600
rect 6604 14560 6610 14572
rect 18506 14560 18512 14572
rect 18564 14600 18570 14612
rect 20898 14600 20904 14612
rect 18564 14572 20904 14600
rect 18564 14560 18570 14572
rect 20898 14560 20904 14572
rect 20956 14560 20962 14612
rect 21266 14560 21272 14612
rect 21324 14600 21330 14612
rect 21453 14603 21511 14609
rect 21453 14600 21465 14603
rect 21324 14572 21465 14600
rect 21324 14560 21330 14572
rect 21453 14569 21465 14572
rect 21499 14569 21511 14603
rect 21453 14563 21511 14569
rect 21910 14560 21916 14612
rect 21968 14560 21974 14612
rect 27890 14560 27896 14612
rect 27948 14600 27954 14612
rect 27985 14603 28043 14609
rect 27985 14600 27997 14603
rect 27948 14572 27997 14600
rect 27948 14560 27954 14572
rect 27985 14569 27997 14572
rect 28031 14569 28043 14603
rect 27985 14563 28043 14569
rect 10226 14532 10232 14544
rect 9508 14504 10232 14532
rect 9508 14473 9536 14504
rect 10226 14492 10232 14504
rect 10284 14492 10290 14544
rect 10962 14492 10968 14544
rect 11020 14532 11026 14544
rect 13081 14535 13139 14541
rect 11020 14504 12020 14532
rect 11020 14492 11026 14504
rect 4525 14467 4583 14473
rect 4525 14433 4537 14467
rect 4571 14464 4583 14467
rect 5077 14467 5135 14473
rect 5077 14464 5089 14467
rect 4571 14436 5089 14464
rect 4571 14433 4583 14436
rect 4525 14427 4583 14433
rect 5077 14433 5089 14436
rect 5123 14433 5135 14467
rect 5077 14427 5135 14433
rect 5353 14467 5411 14473
rect 5353 14433 5365 14467
rect 5399 14464 5411 14467
rect 7653 14467 7711 14473
rect 7653 14464 7665 14467
rect 5399 14436 7665 14464
rect 5399 14433 5411 14436
rect 5353 14427 5411 14433
rect 7653 14433 7665 14436
rect 7699 14433 7711 14467
rect 7653 14427 7711 14433
rect 9493 14467 9551 14473
rect 9493 14433 9505 14467
rect 9539 14433 9551 14467
rect 9493 14427 9551 14433
rect 9769 14467 9827 14473
rect 9769 14433 9781 14467
rect 9815 14464 9827 14467
rect 10686 14464 10692 14476
rect 9815 14436 10692 14464
rect 9815 14433 9827 14436
rect 9769 14427 9827 14433
rect 10686 14424 10692 14436
rect 10744 14424 10750 14476
rect 11992 14473 12020 14504
rect 13081 14501 13093 14535
rect 13127 14532 13139 14535
rect 13170 14532 13176 14544
rect 13127 14504 13176 14532
rect 13127 14501 13139 14504
rect 13081 14495 13139 14501
rect 13170 14492 13176 14504
rect 13228 14492 13234 14544
rect 13814 14492 13820 14544
rect 13872 14532 13878 14544
rect 14369 14535 14427 14541
rect 14369 14532 14381 14535
rect 13872 14504 14381 14532
rect 13872 14492 13878 14504
rect 14369 14501 14381 14504
rect 14415 14501 14427 14535
rect 14369 14495 14427 14501
rect 20990 14492 20996 14544
rect 21048 14532 21054 14544
rect 21048 14504 26234 14532
rect 21048 14492 21054 14504
rect 10873 14467 10931 14473
rect 10873 14433 10885 14467
rect 10919 14464 10931 14467
rect 11701 14467 11759 14473
rect 11701 14464 11713 14467
rect 10919 14436 11713 14464
rect 10919 14433 10931 14436
rect 10873 14427 10931 14433
rect 11701 14433 11713 14436
rect 11747 14433 11759 14467
rect 11701 14427 11759 14433
rect 11977 14467 12035 14473
rect 11977 14433 11989 14467
rect 12023 14433 12035 14467
rect 11977 14427 12035 14433
rect 14918 14424 14924 14476
rect 14976 14424 14982 14476
rect 17126 14424 17132 14476
rect 17184 14464 17190 14476
rect 19613 14467 19671 14473
rect 19613 14464 19625 14467
rect 17184 14436 19625 14464
rect 17184 14424 17190 14436
rect 19613 14433 19625 14436
rect 19659 14433 19671 14467
rect 19613 14427 19671 14433
rect 4614 14356 4620 14408
rect 4672 14356 4678 14408
rect 7561 14399 7619 14405
rect 7561 14365 7573 14399
rect 7607 14365 7619 14399
rect 7561 14359 7619 14365
rect 5902 14288 5908 14340
rect 5960 14288 5966 14340
rect 6730 14288 6736 14340
rect 6788 14328 6794 14340
rect 7101 14331 7159 14337
rect 7101 14328 7113 14331
rect 6788 14300 7113 14328
rect 6788 14288 6794 14300
rect 7101 14297 7113 14300
rect 7147 14328 7159 14331
rect 7576 14328 7604 14359
rect 9398 14356 9404 14408
rect 9456 14356 9462 14408
rect 10965 14399 11023 14405
rect 10965 14365 10977 14399
rect 11011 14396 11023 14399
rect 11606 14396 11612 14408
rect 11011 14368 11612 14396
rect 11011 14365 11023 14368
rect 10965 14359 11023 14365
rect 11606 14356 11612 14368
rect 11664 14356 11670 14408
rect 11790 14356 11796 14408
rect 11848 14356 11854 14408
rect 11885 14399 11943 14405
rect 11885 14365 11897 14399
rect 11931 14365 11943 14399
rect 11885 14359 11943 14365
rect 12161 14399 12219 14405
rect 12161 14365 12173 14399
rect 12207 14396 12219 14399
rect 12434 14396 12440 14408
rect 12207 14368 12440 14396
rect 12207 14365 12219 14368
rect 12161 14359 12219 14365
rect 7147 14300 7604 14328
rect 7147 14297 7159 14300
rect 7101 14291 7159 14297
rect 11514 14220 11520 14272
rect 11572 14220 11578 14272
rect 11900 14260 11928 14359
rect 12434 14356 12440 14368
rect 12492 14356 12498 14408
rect 13265 14399 13323 14405
rect 13265 14365 13277 14399
rect 13311 14396 13323 14399
rect 14182 14396 14188 14408
rect 13311 14368 14188 14396
rect 13311 14365 13323 14368
rect 13265 14359 13323 14365
rect 14182 14356 14188 14368
rect 14240 14356 14246 14408
rect 14461 14399 14519 14405
rect 14461 14365 14473 14399
rect 14507 14365 14519 14399
rect 19628 14396 19656 14427
rect 20898 14424 20904 14476
rect 20956 14464 20962 14476
rect 24394 14464 24400 14476
rect 20956 14436 24400 14464
rect 20956 14424 20962 14436
rect 24394 14424 24400 14436
rect 24452 14424 24458 14476
rect 24578 14424 24584 14476
rect 24636 14464 24642 14476
rect 24673 14467 24731 14473
rect 24673 14464 24685 14467
rect 24636 14436 24685 14464
rect 24636 14424 24642 14436
rect 24673 14433 24685 14436
rect 24719 14433 24731 14467
rect 24673 14427 24731 14433
rect 25133 14467 25191 14473
rect 25133 14433 25145 14467
rect 25179 14464 25191 14467
rect 25590 14464 25596 14476
rect 25179 14436 25596 14464
rect 25179 14433 25191 14436
rect 25133 14427 25191 14433
rect 25590 14424 25596 14436
rect 25648 14424 25654 14476
rect 21637 14399 21695 14405
rect 14461 14359 14519 14365
rect 15028 14368 16574 14396
rect 19628 14368 20116 14396
rect 12066 14288 12072 14340
rect 12124 14328 12130 14340
rect 14476 14328 14504 14359
rect 15028 14328 15056 14368
rect 12124 14300 15056 14328
rect 15188 14331 15246 14337
rect 12124 14288 12130 14300
rect 15188 14297 15200 14331
rect 15234 14328 15246 14331
rect 15562 14328 15568 14340
rect 15234 14300 15568 14328
rect 15234 14297 15246 14300
rect 15188 14291 15246 14297
rect 15562 14288 15568 14300
rect 15620 14288 15626 14340
rect 16546 14328 16574 14368
rect 16758 14328 16764 14340
rect 16546 14300 16764 14328
rect 16758 14288 16764 14300
rect 16816 14288 16822 14340
rect 19880 14331 19938 14337
rect 19880 14297 19892 14331
rect 19926 14328 19938 14331
rect 19978 14328 19984 14340
rect 19926 14300 19984 14328
rect 19926 14297 19938 14300
rect 19880 14291 19938 14297
rect 19978 14288 19984 14300
rect 20036 14288 20042 14340
rect 20088 14328 20116 14368
rect 21637 14365 21649 14399
rect 21683 14365 21695 14399
rect 21637 14359 21695 14365
rect 20088 14300 21404 14328
rect 12434 14260 12440 14272
rect 11900 14232 12440 14260
rect 12434 14220 12440 14232
rect 12492 14220 12498 14272
rect 16298 14220 16304 14272
rect 16356 14220 16362 14272
rect 16482 14220 16488 14272
rect 16540 14260 16546 14272
rect 20898 14260 20904 14272
rect 16540 14232 20904 14260
rect 16540 14220 16546 14232
rect 20898 14220 20904 14232
rect 20956 14220 20962 14272
rect 20990 14220 20996 14272
rect 21048 14220 21054 14272
rect 21376 14260 21404 14300
rect 21450 14288 21456 14340
rect 21508 14288 21514 14340
rect 21542 14288 21548 14340
rect 21600 14328 21606 14340
rect 21652 14328 21680 14359
rect 21726 14356 21732 14408
rect 21784 14356 21790 14408
rect 21600 14300 21680 14328
rect 24412 14328 24440 14424
rect 24762 14356 24768 14408
rect 24820 14356 24826 14408
rect 26206 14396 26234 14504
rect 27448 14436 28764 14464
rect 27448 14405 27476 14436
rect 28736 14408 28764 14436
rect 27433 14399 27491 14405
rect 27433 14396 27445 14399
rect 26206 14368 27445 14396
rect 27433 14365 27445 14368
rect 27479 14365 27491 14399
rect 27433 14359 27491 14365
rect 27798 14356 27804 14408
rect 27856 14396 27862 14408
rect 28077 14399 28135 14405
rect 28077 14396 28089 14399
rect 27856 14368 28089 14396
rect 27856 14356 27862 14368
rect 28077 14365 28089 14368
rect 28123 14365 28135 14399
rect 28077 14359 28135 14365
rect 25682 14328 25688 14340
rect 24412 14300 25688 14328
rect 21600 14288 21606 14300
rect 25682 14288 25688 14300
rect 25740 14288 25746 14340
rect 28092 14328 28120 14359
rect 28718 14356 28724 14408
rect 28776 14356 28782 14408
rect 30282 14356 30288 14408
rect 30340 14356 30346 14408
rect 29638 14328 29644 14340
rect 28092 14300 29644 14328
rect 29638 14288 29644 14300
rect 29696 14288 29702 14340
rect 30009 14331 30067 14337
rect 30009 14297 30021 14331
rect 30055 14328 30067 14331
rect 31018 14328 31024 14340
rect 30055 14300 31024 14328
rect 30055 14297 30067 14300
rect 30009 14291 30067 14297
rect 31018 14288 31024 14300
rect 31076 14288 31082 14340
rect 23750 14260 23756 14272
rect 21376 14232 23756 14260
rect 23750 14220 23756 14232
rect 23808 14220 23814 14272
rect 27341 14263 27399 14269
rect 27341 14229 27353 14263
rect 27387 14260 27399 14263
rect 27522 14260 27528 14272
rect 27387 14232 27528 14260
rect 27387 14229 27399 14232
rect 27341 14223 27399 14229
rect 27522 14220 27528 14232
rect 27580 14220 27586 14272
rect 28626 14220 28632 14272
rect 28684 14220 28690 14272
rect 1104 14170 30976 14192
rect 1104 14118 8378 14170
rect 8430 14118 8442 14170
rect 8494 14118 8506 14170
rect 8558 14118 8570 14170
rect 8622 14118 8634 14170
rect 8686 14118 15806 14170
rect 15858 14118 15870 14170
rect 15922 14118 15934 14170
rect 15986 14118 15998 14170
rect 16050 14118 16062 14170
rect 16114 14118 23234 14170
rect 23286 14118 23298 14170
rect 23350 14118 23362 14170
rect 23414 14118 23426 14170
rect 23478 14118 23490 14170
rect 23542 14118 30662 14170
rect 30714 14118 30726 14170
rect 30778 14118 30790 14170
rect 30842 14118 30854 14170
rect 30906 14118 30918 14170
rect 30970 14118 30976 14170
rect 1104 14096 30976 14118
rect 4614 14016 4620 14068
rect 4672 14056 4678 14068
rect 5166 14056 5172 14068
rect 4672 14028 5172 14056
rect 4672 14016 4678 14028
rect 5166 14016 5172 14028
rect 5224 14056 5230 14068
rect 5905 14059 5963 14065
rect 5905 14056 5917 14059
rect 5224 14028 5917 14056
rect 5224 14016 5230 14028
rect 5905 14025 5917 14028
rect 5951 14056 5963 14059
rect 9398 14056 9404 14068
rect 5951 14028 9404 14056
rect 5951 14025 5963 14028
rect 5905 14019 5963 14025
rect 9398 14016 9404 14028
rect 9456 14016 9462 14068
rect 14182 14016 14188 14068
rect 14240 14016 14246 14068
rect 15562 14016 15568 14068
rect 15620 14016 15626 14068
rect 16025 14059 16083 14065
rect 16025 14025 16037 14059
rect 16071 14056 16083 14059
rect 16298 14056 16304 14068
rect 16071 14028 16304 14056
rect 16071 14025 16083 14028
rect 16025 14019 16083 14025
rect 16298 14016 16304 14028
rect 16356 14016 16362 14068
rect 16390 14016 16396 14068
rect 16448 14056 16454 14068
rect 16853 14059 16911 14065
rect 16853 14056 16865 14059
rect 16448 14028 16865 14056
rect 16448 14016 16454 14028
rect 16853 14025 16865 14028
rect 16899 14025 16911 14059
rect 16853 14019 16911 14025
rect 17218 14016 17224 14068
rect 17276 14016 17282 14068
rect 19978 14016 19984 14068
rect 20036 14016 20042 14068
rect 20441 14059 20499 14065
rect 20441 14025 20453 14059
rect 20487 14056 20499 14059
rect 20990 14056 20996 14068
rect 20487 14028 20996 14056
rect 20487 14025 20499 14028
rect 20441 14019 20499 14025
rect 20990 14016 20996 14028
rect 21048 14016 21054 14068
rect 22462 14016 22468 14068
rect 22520 14056 22526 14068
rect 26053 14059 26111 14065
rect 26053 14056 26065 14059
rect 22520 14028 26065 14056
rect 22520 14016 22526 14028
rect 26053 14025 26065 14028
rect 26099 14025 26111 14059
rect 26053 14019 26111 14025
rect 29638 14016 29644 14068
rect 29696 14056 29702 14068
rect 30101 14059 30159 14065
rect 30101 14056 30113 14059
rect 29696 14028 30113 14056
rect 29696 14016 29702 14028
rect 30101 14025 30113 14028
rect 30147 14025 30159 14059
rect 30101 14019 30159 14025
rect 4430 13948 4436 14000
rect 4488 13948 4494 14000
rect 5810 13988 5816 14000
rect 5658 13960 5816 13988
rect 5810 13948 5816 13960
rect 5868 13948 5874 14000
rect 16316 13988 16344 14016
rect 16316 13960 22508 13988
rect 6730 13880 6736 13932
rect 6788 13880 6794 13932
rect 11882 13880 11888 13932
rect 11940 13920 11946 13932
rect 12526 13929 12532 13932
rect 12253 13923 12311 13929
rect 12253 13920 12265 13923
rect 11940 13892 12265 13920
rect 11940 13880 11946 13892
rect 12253 13889 12265 13892
rect 12299 13889 12311 13923
rect 12253 13883 12311 13889
rect 12520 13883 12532 13929
rect 12526 13880 12532 13883
rect 12584 13880 12590 13932
rect 14090 13880 14096 13932
rect 14148 13880 14154 13932
rect 14918 13880 14924 13932
rect 14976 13920 14982 13932
rect 15933 13923 15991 13929
rect 15933 13920 15945 13923
rect 14976 13892 15945 13920
rect 14976 13880 14982 13892
rect 15933 13889 15945 13892
rect 15979 13920 15991 13923
rect 16482 13920 16488 13932
rect 15979 13892 16488 13920
rect 15979 13889 15991 13892
rect 15933 13883 15991 13889
rect 16482 13880 16488 13892
rect 16540 13880 16546 13932
rect 17494 13880 17500 13932
rect 17552 13920 17558 13932
rect 20349 13923 20407 13929
rect 20349 13920 20361 13923
rect 17552 13892 20361 13920
rect 17552 13880 17558 13892
rect 20349 13889 20361 13892
rect 20395 13889 20407 13923
rect 20349 13883 20407 13889
rect 20438 13880 20444 13932
rect 20496 13920 20502 13932
rect 21726 13920 21732 13932
rect 20496 13892 21732 13920
rect 20496 13880 20502 13892
rect 21726 13880 21732 13892
rect 21784 13880 21790 13932
rect 4154 13812 4160 13864
rect 4212 13812 4218 13864
rect 6178 13812 6184 13864
rect 6236 13852 6242 13864
rect 6641 13855 6699 13861
rect 6641 13852 6653 13855
rect 6236 13824 6653 13852
rect 6236 13812 6242 13824
rect 6641 13821 6653 13824
rect 6687 13821 6699 13855
rect 6641 13815 6699 13821
rect 7101 13855 7159 13861
rect 7101 13821 7113 13855
rect 7147 13852 7159 13855
rect 7190 13852 7196 13864
rect 7147 13824 7196 13852
rect 7147 13821 7159 13824
rect 7101 13815 7159 13821
rect 7190 13812 7196 13824
rect 7248 13812 7254 13864
rect 16209 13855 16267 13861
rect 16209 13821 16221 13855
rect 16255 13821 16267 13855
rect 16209 13815 16267 13821
rect 16224 13784 16252 13815
rect 17310 13812 17316 13864
rect 17368 13812 17374 13864
rect 17402 13812 17408 13864
rect 17460 13812 17466 13864
rect 22480 13861 22508 13960
rect 23106 13948 23112 14000
rect 23164 13988 23170 14000
rect 23385 13991 23443 13997
rect 23385 13988 23397 13991
rect 23164 13960 23397 13988
rect 23164 13948 23170 13960
rect 23385 13957 23397 13960
rect 23431 13957 23443 13991
rect 23385 13951 23443 13957
rect 25590 13948 25596 14000
rect 25648 13948 25654 14000
rect 28626 13988 28632 14000
rect 28368 13960 28632 13988
rect 22557 13923 22615 13929
rect 22557 13889 22569 13923
rect 22603 13920 22615 13923
rect 23014 13920 23020 13932
rect 22603 13892 23020 13920
rect 22603 13889 22615 13892
rect 22557 13883 22615 13889
rect 23014 13880 23020 13892
rect 23072 13880 23078 13932
rect 25866 13880 25872 13932
rect 25924 13880 25930 13932
rect 26510 13920 26516 13932
rect 26206 13892 26516 13920
rect 20533 13855 20591 13861
rect 20533 13821 20545 13855
rect 20579 13821 20591 13855
rect 20533 13815 20591 13821
rect 22465 13855 22523 13861
rect 22465 13821 22477 13855
rect 22511 13821 22523 13855
rect 22465 13815 22523 13821
rect 22925 13855 22983 13861
rect 22925 13821 22937 13855
rect 22971 13852 22983 13855
rect 25685 13855 25743 13861
rect 25685 13852 25697 13855
rect 22971 13824 25697 13852
rect 22971 13821 22983 13824
rect 22925 13815 22983 13821
rect 25685 13821 25697 13824
rect 25731 13821 25743 13855
rect 25685 13815 25743 13821
rect 16224 13756 16574 13784
rect 13170 13676 13176 13728
rect 13228 13716 13234 13728
rect 13633 13719 13691 13725
rect 13633 13716 13645 13719
rect 13228 13688 13645 13716
rect 13228 13676 13234 13688
rect 13633 13685 13645 13688
rect 13679 13685 13691 13719
rect 16546 13716 16574 13756
rect 17420 13716 17448 13812
rect 20070 13744 20076 13796
rect 20128 13784 20134 13796
rect 20548 13784 20576 13815
rect 20128 13756 20576 13784
rect 20128 13744 20134 13756
rect 24762 13744 24768 13796
rect 24820 13784 24826 13796
rect 26206 13784 26234 13892
rect 26510 13880 26516 13892
rect 26568 13920 26574 13932
rect 28368 13929 28396 13960
rect 28626 13948 28632 13960
rect 28684 13948 28690 14000
rect 27157 13923 27215 13929
rect 27157 13920 27169 13923
rect 26568 13892 27169 13920
rect 26568 13880 26574 13892
rect 27157 13889 27169 13892
rect 27203 13889 27215 13923
rect 27157 13883 27215 13889
rect 28353 13923 28411 13929
rect 28353 13889 28365 13923
rect 28399 13889 28411 13923
rect 28353 13883 28411 13889
rect 29730 13880 29736 13932
rect 29788 13880 29794 13932
rect 28626 13812 28632 13864
rect 28684 13812 28690 13864
rect 24820 13756 26234 13784
rect 24820 13744 24826 13756
rect 16546 13688 17448 13716
rect 13633 13679 13691 13685
rect 24578 13676 24584 13728
rect 24636 13716 24642 13728
rect 24673 13719 24731 13725
rect 24673 13716 24685 13719
rect 24636 13688 24685 13716
rect 24636 13676 24642 13688
rect 24673 13685 24685 13688
rect 24719 13685 24731 13719
rect 24673 13679 24731 13685
rect 24946 13676 24952 13728
rect 25004 13716 25010 13728
rect 25593 13719 25651 13725
rect 25593 13716 25605 13719
rect 25004 13688 25605 13716
rect 25004 13676 25010 13688
rect 25593 13685 25605 13688
rect 25639 13685 25651 13719
rect 25593 13679 25651 13685
rect 27249 13719 27307 13725
rect 27249 13685 27261 13719
rect 27295 13716 27307 13719
rect 27338 13716 27344 13728
rect 27295 13688 27344 13716
rect 27295 13685 27307 13688
rect 27249 13679 27307 13685
rect 27338 13676 27344 13688
rect 27396 13676 27402 13728
rect 1104 13626 30820 13648
rect 1104 13574 4664 13626
rect 4716 13574 4728 13626
rect 4780 13574 4792 13626
rect 4844 13574 4856 13626
rect 4908 13574 4920 13626
rect 4972 13574 12092 13626
rect 12144 13574 12156 13626
rect 12208 13574 12220 13626
rect 12272 13574 12284 13626
rect 12336 13574 12348 13626
rect 12400 13574 19520 13626
rect 19572 13574 19584 13626
rect 19636 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 26948 13626
rect 27000 13574 27012 13626
rect 27064 13574 27076 13626
rect 27128 13574 27140 13626
rect 27192 13574 27204 13626
rect 27256 13574 30820 13626
rect 1104 13552 30820 13574
rect 4154 13472 4160 13524
rect 4212 13512 4218 13524
rect 4801 13515 4859 13521
rect 4801 13512 4813 13515
rect 4212 13484 4813 13512
rect 4212 13472 4218 13484
rect 4801 13481 4813 13484
rect 4847 13481 4859 13515
rect 4801 13475 4859 13481
rect 12526 13472 12532 13524
rect 12584 13512 12590 13524
rect 12713 13515 12771 13521
rect 12713 13512 12725 13515
rect 12584 13484 12725 13512
rect 12584 13472 12590 13484
rect 12713 13481 12725 13484
rect 12759 13481 12771 13515
rect 12713 13475 12771 13481
rect 18601 13515 18659 13521
rect 18601 13481 18613 13515
rect 18647 13512 18659 13515
rect 20438 13512 20444 13524
rect 18647 13484 20444 13512
rect 18647 13481 18659 13484
rect 18601 13475 18659 13481
rect 20438 13472 20444 13484
rect 20496 13472 20502 13524
rect 21085 13515 21143 13521
rect 21085 13481 21097 13515
rect 21131 13512 21143 13515
rect 21542 13512 21548 13524
rect 21131 13484 21548 13512
rect 21131 13481 21143 13484
rect 21085 13475 21143 13481
rect 21542 13472 21548 13484
rect 21600 13472 21606 13524
rect 28626 13472 28632 13524
rect 28684 13512 28690 13524
rect 29825 13515 29883 13521
rect 29825 13512 29837 13515
rect 28684 13484 29837 13512
rect 28684 13472 28690 13484
rect 29825 13481 29837 13484
rect 29871 13481 29883 13515
rect 29825 13475 29883 13481
rect 28718 13404 28724 13456
rect 28776 13404 28782 13456
rect 5258 13336 5264 13388
rect 5316 13376 5322 13388
rect 5721 13379 5779 13385
rect 5721 13376 5733 13379
rect 5316 13348 5733 13376
rect 5316 13336 5322 13348
rect 5721 13345 5733 13348
rect 5767 13345 5779 13379
rect 5721 13339 5779 13345
rect 9122 13336 9128 13388
rect 9180 13336 9186 13388
rect 13170 13336 13176 13388
rect 13228 13336 13234 13388
rect 13262 13336 13268 13388
rect 13320 13376 13326 13388
rect 13357 13379 13415 13385
rect 13357 13376 13369 13379
rect 13320 13348 13369 13376
rect 13320 13336 13326 13348
rect 13357 13345 13369 13348
rect 13403 13376 13415 13379
rect 15102 13376 15108 13388
rect 13403 13348 15108 13376
rect 13403 13345 13415 13348
rect 13357 13339 13415 13345
rect 15102 13336 15108 13348
rect 15160 13336 15166 13388
rect 17310 13336 17316 13388
rect 17368 13376 17374 13388
rect 18141 13379 18199 13385
rect 18141 13376 18153 13379
rect 17368 13348 18153 13376
rect 17368 13336 17374 13348
rect 18141 13345 18153 13348
rect 18187 13345 18199 13379
rect 18141 13339 18199 13345
rect 20809 13379 20867 13385
rect 20809 13345 20821 13379
rect 20855 13376 20867 13379
rect 20990 13376 20996 13388
rect 20855 13348 20996 13376
rect 20855 13345 20867 13348
rect 20809 13339 20867 13345
rect 20990 13336 20996 13348
rect 21048 13336 21054 13388
rect 26973 13379 27031 13385
rect 26973 13345 26985 13379
rect 27019 13376 27031 13379
rect 27338 13376 27344 13388
rect 27019 13348 27344 13376
rect 27019 13345 27031 13348
rect 26973 13339 27031 13345
rect 27338 13336 27344 13348
rect 27396 13336 27402 13388
rect 4893 13311 4951 13317
rect 4893 13277 4905 13311
rect 4939 13308 4951 13311
rect 4982 13308 4988 13320
rect 4939 13280 4988 13308
rect 4939 13277 4951 13280
rect 4893 13271 4951 13277
rect 4982 13268 4988 13280
rect 5040 13268 5046 13320
rect 6825 13311 6883 13317
rect 6825 13277 6837 13311
rect 6871 13308 6883 13311
rect 8018 13308 8024 13320
rect 6871 13280 8024 13308
rect 6871 13277 6883 13280
rect 6825 13271 6883 13277
rect 8018 13268 8024 13280
rect 8076 13308 8082 13320
rect 8076 13280 13400 13308
rect 8076 13268 8082 13280
rect 13372 13252 13400 13280
rect 16206 13268 16212 13320
rect 16264 13268 16270 13320
rect 18230 13268 18236 13320
rect 18288 13268 18294 13320
rect 20717 13311 20775 13317
rect 20717 13277 20729 13311
rect 20763 13308 20775 13311
rect 22922 13308 22928 13320
rect 20763 13280 22928 13308
rect 20763 13277 20775 13280
rect 20717 13271 20775 13277
rect 22922 13268 22928 13280
rect 22980 13268 22986 13320
rect 24029 13311 24087 13317
rect 24029 13277 24041 13311
rect 24075 13308 24087 13311
rect 24762 13308 24768 13320
rect 24075 13280 24768 13308
rect 24075 13277 24087 13280
rect 24029 13271 24087 13277
rect 24762 13268 24768 13280
rect 24820 13268 24826 13320
rect 29638 13268 29644 13320
rect 29696 13308 29702 13320
rect 29917 13311 29975 13317
rect 29917 13308 29929 13311
rect 29696 13280 29929 13308
rect 29696 13268 29702 13280
rect 29917 13277 29929 13280
rect 29963 13277 29975 13311
rect 29917 13271 29975 13277
rect 9214 13200 9220 13252
rect 9272 13240 9278 13252
rect 9370 13243 9428 13249
rect 9370 13240 9382 13243
rect 9272 13212 9382 13240
rect 9272 13200 9278 13212
rect 9370 13209 9382 13212
rect 9416 13209 9428 13243
rect 9370 13203 9428 13209
rect 9490 13200 9496 13252
rect 9548 13240 9554 13252
rect 9548 13212 12434 13240
rect 9548 13200 9554 13212
rect 9582 13132 9588 13184
rect 9640 13172 9646 13184
rect 10505 13175 10563 13181
rect 10505 13172 10517 13175
rect 9640 13144 10517 13172
rect 9640 13132 9646 13144
rect 10505 13141 10517 13144
rect 10551 13141 10563 13175
rect 12406 13172 12434 13212
rect 13354 13200 13360 13252
rect 13412 13200 13418 13252
rect 16476 13243 16534 13249
rect 16476 13209 16488 13243
rect 16522 13240 16534 13243
rect 16850 13240 16856 13252
rect 16522 13212 16856 13240
rect 16522 13209 16534 13212
rect 16476 13203 16534 13209
rect 16850 13200 16856 13212
rect 16908 13200 16914 13252
rect 24578 13200 24584 13252
rect 24636 13200 24642 13252
rect 27249 13243 27307 13249
rect 27249 13209 27261 13243
rect 27295 13240 27307 13243
rect 27522 13240 27528 13252
rect 27295 13212 27528 13240
rect 27295 13209 27307 13212
rect 27249 13203 27307 13209
rect 27522 13200 27528 13212
rect 27580 13200 27586 13252
rect 28258 13200 28264 13252
rect 28316 13200 28322 13252
rect 13081 13175 13139 13181
rect 13081 13172 13093 13175
rect 12406 13144 13093 13172
rect 10505 13135 10563 13141
rect 13081 13141 13093 13144
rect 13127 13172 13139 13175
rect 17494 13172 17500 13184
rect 13127 13144 17500 13172
rect 13127 13141 13139 13144
rect 13081 13135 13139 13141
rect 17494 13132 17500 13144
rect 17552 13132 17558 13184
rect 17586 13132 17592 13184
rect 17644 13132 17650 13184
rect 23937 13175 23995 13181
rect 23937 13141 23949 13175
rect 23983 13172 23995 13175
rect 25038 13172 25044 13184
rect 23983 13144 25044 13172
rect 23983 13141 23995 13144
rect 23937 13135 23995 13141
rect 25038 13132 25044 13144
rect 25096 13132 25102 13184
rect 26050 13132 26056 13184
rect 26108 13132 26114 13184
rect 1104 13082 30976 13104
rect 1104 13030 8378 13082
rect 8430 13030 8442 13082
rect 8494 13030 8506 13082
rect 8558 13030 8570 13082
rect 8622 13030 8634 13082
rect 8686 13030 15806 13082
rect 15858 13030 15870 13082
rect 15922 13030 15934 13082
rect 15986 13030 15998 13082
rect 16050 13030 16062 13082
rect 16114 13030 23234 13082
rect 23286 13030 23298 13082
rect 23350 13030 23362 13082
rect 23414 13030 23426 13082
rect 23478 13030 23490 13082
rect 23542 13030 30662 13082
rect 30714 13030 30726 13082
rect 30778 13030 30790 13082
rect 30842 13030 30854 13082
rect 30906 13030 30918 13082
rect 30970 13030 30976 13082
rect 1104 13008 30976 13030
rect 5810 12928 5816 12980
rect 5868 12928 5874 12980
rect 9214 12928 9220 12980
rect 9272 12928 9278 12980
rect 9582 12928 9588 12980
rect 9640 12968 9646 12980
rect 9677 12971 9735 12977
rect 9677 12968 9689 12971
rect 9640 12940 9689 12968
rect 9640 12928 9646 12940
rect 9677 12937 9689 12940
rect 9723 12937 9735 12971
rect 9677 12931 9735 12937
rect 14737 12971 14795 12977
rect 14737 12937 14749 12971
rect 14783 12937 14795 12971
rect 14737 12931 14795 12937
rect 6914 12860 6920 12912
rect 6972 12900 6978 12912
rect 7469 12903 7527 12909
rect 7469 12900 7481 12903
rect 6972 12872 7481 12900
rect 6972 12860 6978 12872
rect 7469 12869 7481 12872
rect 7515 12869 7527 12903
rect 13164 12903 13222 12909
rect 7469 12863 7527 12869
rect 7576 12872 12434 12900
rect 5169 12835 5227 12841
rect 5169 12801 5181 12835
rect 5215 12832 5227 12835
rect 5258 12832 5264 12844
rect 5215 12804 5264 12832
rect 5215 12801 5227 12804
rect 5169 12795 5227 12801
rect 5258 12792 5264 12804
rect 5316 12792 5322 12844
rect 5350 12792 5356 12844
rect 5408 12792 5414 12844
rect 7098 12792 7104 12844
rect 7156 12832 7162 12844
rect 7285 12835 7343 12841
rect 7285 12832 7297 12835
rect 7156 12804 7297 12832
rect 7156 12792 7162 12804
rect 7285 12801 7297 12804
rect 7331 12832 7343 12835
rect 7576 12832 7604 12872
rect 7331 12804 7604 12832
rect 7331 12801 7343 12804
rect 7285 12795 7343 12801
rect 7650 12792 7656 12844
rect 7708 12832 7714 12844
rect 8389 12835 8447 12841
rect 8389 12832 8401 12835
rect 7708 12804 8401 12832
rect 7708 12792 7714 12804
rect 8389 12801 8401 12804
rect 8435 12801 8447 12835
rect 8389 12795 8447 12801
rect 9490 12792 9496 12844
rect 9548 12832 9554 12844
rect 9585 12835 9643 12841
rect 9585 12832 9597 12835
rect 9548 12804 9597 12832
rect 9548 12792 9554 12804
rect 9585 12801 9597 12804
rect 9631 12801 9643 12835
rect 12406 12832 12434 12872
rect 13164 12869 13176 12903
rect 13210 12900 13222 12903
rect 14752 12900 14780 12931
rect 16850 12928 16856 12980
rect 16908 12928 16914 12980
rect 26050 12928 26056 12980
rect 26108 12968 26114 12980
rect 26108 12940 28120 12968
rect 26108 12928 26114 12940
rect 13210 12872 14780 12900
rect 13210 12869 13222 12872
rect 13164 12863 13222 12869
rect 25038 12860 25044 12912
rect 25096 12860 25102 12912
rect 12406 12804 14320 12832
rect 9585 12795 9643 12801
rect 5276 12764 5304 12792
rect 5442 12764 5448 12776
rect 5276 12736 5448 12764
rect 5442 12724 5448 12736
rect 5500 12724 5506 12776
rect 8294 12724 8300 12776
rect 8352 12724 8358 12776
rect 9861 12767 9919 12773
rect 9861 12733 9873 12767
rect 9907 12733 9919 12767
rect 9861 12727 9919 12733
rect 9122 12656 9128 12708
rect 9180 12696 9186 12708
rect 9876 12696 9904 12727
rect 11882 12724 11888 12776
rect 11940 12764 11946 12776
rect 12897 12767 12955 12773
rect 12897 12764 12909 12767
rect 11940 12736 12909 12764
rect 11940 12724 11946 12736
rect 12897 12733 12909 12736
rect 12943 12733 12955 12767
rect 12897 12727 12955 12733
rect 14292 12764 14320 12804
rect 14918 12792 14924 12844
rect 14976 12832 14982 12844
rect 15105 12835 15163 12841
rect 15105 12832 15117 12835
rect 14976 12804 15117 12832
rect 14976 12792 14982 12804
rect 15105 12801 15117 12804
rect 15151 12801 15163 12835
rect 15105 12795 15163 12801
rect 17221 12835 17279 12841
rect 17221 12801 17233 12835
rect 17267 12801 17279 12835
rect 17221 12795 17279 12801
rect 17313 12835 17371 12841
rect 17313 12801 17325 12835
rect 17359 12832 17371 12835
rect 17586 12832 17592 12844
rect 17359 12804 17592 12832
rect 17359 12801 17371 12804
rect 17313 12795 17371 12801
rect 15197 12767 15255 12773
rect 15197 12764 15209 12767
rect 14292 12736 15209 12764
rect 12802 12696 12808 12708
rect 9180 12668 12808 12696
rect 9180 12656 9186 12668
rect 12802 12656 12808 12668
rect 12860 12656 12866 12708
rect 14292 12705 14320 12736
rect 15197 12733 15209 12736
rect 15243 12733 15255 12767
rect 15197 12727 15255 12733
rect 15289 12767 15347 12773
rect 15289 12733 15301 12767
rect 15335 12733 15347 12767
rect 17236 12764 17264 12795
rect 17586 12792 17592 12804
rect 17644 12832 17650 12844
rect 19613 12835 19671 12841
rect 17644 12804 19564 12832
rect 17644 12792 17650 12804
rect 17236 12736 17356 12764
rect 15289 12727 15347 12733
rect 14277 12699 14335 12705
rect 14277 12665 14289 12699
rect 14323 12665 14335 12699
rect 14277 12659 14335 12665
rect 15102 12656 15108 12708
rect 15160 12696 15166 12708
rect 15304 12696 15332 12727
rect 15160 12668 15332 12696
rect 17328 12696 17356 12736
rect 17402 12724 17408 12776
rect 17460 12724 17466 12776
rect 19536 12773 19564 12804
rect 19613 12801 19625 12835
rect 19659 12832 19671 12835
rect 19886 12832 19892 12844
rect 19659 12804 19892 12832
rect 19659 12801 19671 12804
rect 19613 12795 19671 12801
rect 19886 12792 19892 12804
rect 19944 12792 19950 12844
rect 22922 12792 22928 12844
rect 22980 12792 22986 12844
rect 23106 12792 23112 12844
rect 23164 12832 23170 12844
rect 23385 12835 23443 12841
rect 23385 12832 23397 12835
rect 23164 12804 23397 12832
rect 23164 12792 23170 12804
rect 23385 12801 23397 12804
rect 23431 12801 23443 12835
rect 23385 12795 23443 12801
rect 24121 12835 24179 12841
rect 24121 12801 24133 12835
rect 24167 12801 24179 12835
rect 24121 12795 24179 12801
rect 19521 12767 19579 12773
rect 19521 12733 19533 12767
rect 19567 12733 19579 12767
rect 19521 12727 19579 12733
rect 19981 12767 20039 12773
rect 19981 12733 19993 12767
rect 20027 12764 20039 12767
rect 21450 12764 21456 12776
rect 20027 12736 21456 12764
rect 20027 12733 20039 12736
rect 19981 12727 20039 12733
rect 21450 12724 21456 12736
rect 21508 12724 21514 12776
rect 22940 12764 22968 12792
rect 23934 12764 23940 12776
rect 22940 12736 23940 12764
rect 23934 12724 23940 12736
rect 23992 12764 23998 12776
rect 24136 12764 24164 12795
rect 26142 12792 26148 12844
rect 26200 12792 26206 12844
rect 27430 12792 27436 12844
rect 27488 12792 27494 12844
rect 28092 12832 28120 12940
rect 28169 12903 28227 12909
rect 28169 12869 28181 12903
rect 28215 12900 28227 12903
rect 28258 12900 28264 12912
rect 28215 12872 28264 12900
rect 28215 12869 28227 12872
rect 28169 12863 28227 12869
rect 28258 12860 28264 12872
rect 28316 12860 28322 12912
rect 29730 12860 29736 12912
rect 29788 12860 29794 12912
rect 28350 12832 28356 12844
rect 28092 12818 28356 12832
rect 28106 12804 28356 12818
rect 28350 12792 28356 12804
rect 28408 12832 28414 12844
rect 28408 12804 29118 12832
rect 28408 12792 28414 12804
rect 23992 12736 24164 12764
rect 24213 12767 24271 12773
rect 23992 12724 23998 12736
rect 24213 12733 24225 12767
rect 24259 12764 24271 12767
rect 24765 12767 24823 12773
rect 24765 12764 24777 12767
rect 24259 12736 24777 12764
rect 24259 12733 24271 12736
rect 24213 12727 24271 12733
rect 24765 12733 24777 12736
rect 24811 12733 24823 12767
rect 24765 12727 24823 12733
rect 26510 12724 26516 12776
rect 26568 12724 26574 12776
rect 27448 12764 27476 12792
rect 27982 12764 27988 12776
rect 27448 12736 27988 12764
rect 27982 12724 27988 12736
rect 28040 12764 28046 12776
rect 29181 12767 29239 12773
rect 29181 12764 29193 12767
rect 28040 12736 29193 12764
rect 28040 12724 28046 12736
rect 29181 12733 29193 12736
rect 29227 12733 29239 12767
rect 29181 12727 29239 12733
rect 17770 12696 17776 12708
rect 17328 12668 17776 12696
rect 15160 12656 15166 12668
rect 17770 12656 17776 12668
rect 17828 12696 17834 12708
rect 19426 12696 19432 12708
rect 17828 12668 19432 12696
rect 17828 12656 17834 12668
rect 19426 12656 19432 12668
rect 19484 12696 19490 12708
rect 19484 12668 23612 12696
rect 19484 12656 19490 12668
rect 7653 12631 7711 12637
rect 7653 12597 7665 12631
rect 7699 12628 7711 12631
rect 7834 12628 7840 12640
rect 7699 12600 7840 12628
rect 7699 12597 7711 12600
rect 7653 12591 7711 12597
rect 7834 12588 7840 12600
rect 7892 12588 7898 12640
rect 8757 12631 8815 12637
rect 8757 12597 8769 12631
rect 8803 12628 8815 12631
rect 10410 12628 10416 12640
rect 8803 12600 10416 12628
rect 8803 12597 8815 12600
rect 8757 12591 8815 12597
rect 10410 12588 10416 12600
rect 10468 12588 10474 12640
rect 22462 12588 22468 12640
rect 22520 12628 22526 12640
rect 22833 12631 22891 12637
rect 22833 12628 22845 12631
rect 22520 12600 22845 12628
rect 22520 12588 22526 12600
rect 22833 12597 22845 12600
rect 22879 12597 22891 12631
rect 22833 12591 22891 12597
rect 23474 12588 23480 12640
rect 23532 12588 23538 12640
rect 23584 12628 23612 12668
rect 25038 12628 25044 12640
rect 23584 12600 25044 12628
rect 25038 12588 25044 12600
rect 25096 12588 25102 12640
rect 1104 12538 30820 12560
rect 1104 12486 4664 12538
rect 4716 12486 4728 12538
rect 4780 12486 4792 12538
rect 4844 12486 4856 12538
rect 4908 12486 4920 12538
rect 4972 12486 12092 12538
rect 12144 12486 12156 12538
rect 12208 12486 12220 12538
rect 12272 12486 12284 12538
rect 12336 12486 12348 12538
rect 12400 12486 19520 12538
rect 19572 12486 19584 12538
rect 19636 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 26948 12538
rect 27000 12486 27012 12538
rect 27064 12486 27076 12538
rect 27128 12486 27140 12538
rect 27192 12486 27204 12538
rect 27256 12486 30820 12538
rect 1104 12464 30820 12486
rect 17221 12427 17279 12433
rect 17221 12393 17233 12427
rect 17267 12424 17279 12427
rect 17310 12424 17316 12436
rect 17267 12396 17316 12424
rect 17267 12393 17279 12396
rect 17221 12387 17279 12393
rect 17310 12384 17316 12396
rect 17368 12384 17374 12436
rect 23474 12424 23480 12436
rect 22296 12396 23480 12424
rect 7009 12291 7067 12297
rect 7009 12257 7021 12291
rect 7055 12288 7067 12291
rect 22189 12291 22247 12297
rect 7055 12260 7696 12288
rect 7055 12257 7067 12260
rect 7009 12251 7067 12257
rect 4982 12180 4988 12232
rect 5040 12180 5046 12232
rect 5166 12180 5172 12232
rect 5224 12220 5230 12232
rect 5629 12223 5687 12229
rect 5629 12220 5641 12223
rect 5224 12192 5641 12220
rect 5224 12180 5230 12192
rect 5629 12189 5641 12192
rect 5675 12220 5687 12223
rect 6914 12220 6920 12232
rect 5675 12192 6920 12220
rect 5675 12189 5687 12192
rect 5629 12183 5687 12189
rect 6914 12180 6920 12192
rect 6972 12180 6978 12232
rect 7098 12180 7104 12232
rect 7156 12180 7162 12232
rect 7190 12180 7196 12232
rect 7248 12220 7254 12232
rect 7668 12229 7696 12260
rect 22189 12257 22201 12291
rect 22235 12288 22247 12291
rect 22296 12288 22324 12396
rect 23474 12384 23480 12396
rect 23532 12384 23538 12436
rect 23934 12384 23940 12436
rect 23992 12384 23998 12436
rect 27430 12356 27436 12368
rect 25332 12328 27436 12356
rect 22235 12260 22324 12288
rect 22235 12257 22247 12260
rect 22189 12251 22247 12257
rect 22462 12248 22468 12300
rect 22520 12248 22526 12300
rect 22922 12248 22928 12300
rect 22980 12288 22986 12300
rect 25332 12297 25360 12328
rect 27430 12316 27436 12328
rect 27488 12316 27494 12368
rect 25317 12291 25375 12297
rect 25317 12288 25329 12291
rect 22980 12260 25329 12288
rect 22980 12248 22986 12260
rect 25317 12257 25329 12260
rect 25363 12257 25375 12291
rect 25317 12251 25375 12257
rect 26142 12248 26148 12300
rect 26200 12248 26206 12300
rect 7561 12223 7619 12229
rect 7561 12220 7573 12223
rect 7248 12192 7573 12220
rect 7248 12180 7254 12192
rect 7561 12189 7573 12192
rect 7607 12189 7619 12223
rect 7561 12183 7619 12189
rect 7654 12223 7712 12229
rect 7654 12189 7666 12223
rect 7700 12189 7712 12223
rect 7654 12183 7712 12189
rect 7834 12180 7840 12232
rect 7892 12180 7898 12232
rect 8110 12229 8116 12232
rect 8067 12223 8116 12229
rect 8067 12189 8079 12223
rect 8113 12189 8116 12223
rect 8067 12183 8116 12189
rect 8110 12180 8116 12183
rect 8168 12180 8174 12232
rect 11790 12220 11796 12232
rect 8220 12192 11796 12220
rect 4154 12112 4160 12164
rect 4212 12152 4218 12164
rect 5537 12155 5595 12161
rect 5537 12152 5549 12155
rect 4212 12124 5549 12152
rect 4212 12112 4218 12124
rect 5537 12121 5549 12124
rect 5583 12121 5595 12155
rect 5537 12115 5595 12121
rect 7926 12112 7932 12164
rect 7984 12112 7990 12164
rect 4430 12044 4436 12096
rect 4488 12084 4494 12096
rect 8220 12093 8248 12192
rect 11790 12180 11796 12192
rect 11848 12220 11854 12232
rect 12345 12223 12403 12229
rect 12345 12220 12357 12223
rect 11848 12192 12357 12220
rect 11848 12180 11854 12192
rect 12345 12189 12357 12192
rect 12391 12189 12403 12223
rect 12345 12183 12403 12189
rect 12434 12180 12440 12232
rect 12492 12220 12498 12232
rect 12529 12223 12587 12229
rect 12529 12220 12541 12223
rect 12492 12192 12541 12220
rect 12492 12180 12498 12192
rect 12529 12189 12541 12192
rect 12575 12189 12587 12223
rect 12529 12183 12587 12189
rect 15841 12223 15899 12229
rect 15841 12189 15853 12223
rect 15887 12189 15899 12223
rect 15841 12183 15899 12189
rect 16108 12223 16166 12229
rect 16108 12189 16120 12223
rect 16154 12220 16166 12223
rect 16390 12220 16396 12232
rect 16154 12192 16396 12220
rect 16154 12189 16166 12192
rect 16108 12183 16166 12189
rect 15856 12152 15884 12183
rect 16390 12180 16396 12192
rect 16448 12180 16454 12232
rect 17865 12223 17923 12229
rect 17865 12189 17877 12223
rect 17911 12220 17923 12223
rect 18230 12220 18236 12232
rect 17911 12192 18236 12220
rect 17911 12189 17923 12192
rect 17865 12183 17923 12189
rect 18230 12180 18236 12192
rect 18288 12180 18294 12232
rect 26050 12220 26056 12232
rect 25806 12192 26056 12220
rect 26050 12180 26056 12192
rect 26108 12180 26114 12232
rect 16206 12152 16212 12164
rect 15856 12124 16212 12152
rect 16206 12112 16212 12124
rect 16264 12112 16270 12164
rect 23750 12152 23756 12164
rect 23690 12124 23756 12152
rect 23750 12112 23756 12124
rect 23808 12112 23814 12164
rect 4893 12087 4951 12093
rect 4893 12084 4905 12087
rect 4488 12056 4905 12084
rect 4488 12044 4494 12056
rect 4893 12053 4905 12056
rect 4939 12053 4951 12087
rect 4893 12047 4951 12053
rect 8205 12087 8263 12093
rect 8205 12053 8217 12087
rect 8251 12053 8263 12087
rect 8205 12047 8263 12053
rect 12437 12087 12495 12093
rect 12437 12053 12449 12087
rect 12483 12084 12495 12087
rect 12526 12084 12532 12096
rect 12483 12056 12532 12084
rect 12483 12053 12495 12056
rect 12437 12047 12495 12053
rect 12526 12044 12532 12056
rect 12584 12044 12590 12096
rect 17310 12044 17316 12096
rect 17368 12084 17374 12096
rect 17773 12087 17831 12093
rect 17773 12084 17785 12087
rect 17368 12056 17785 12084
rect 17368 12044 17374 12056
rect 17773 12053 17785 12056
rect 17819 12053 17831 12087
rect 17773 12047 17831 12053
rect 1104 11994 30976 12016
rect 1104 11942 8378 11994
rect 8430 11942 8442 11994
rect 8494 11942 8506 11994
rect 8558 11942 8570 11994
rect 8622 11942 8634 11994
rect 8686 11942 15806 11994
rect 15858 11942 15870 11994
rect 15922 11942 15934 11994
rect 15986 11942 15998 11994
rect 16050 11942 16062 11994
rect 16114 11942 23234 11994
rect 23286 11942 23298 11994
rect 23350 11942 23362 11994
rect 23414 11942 23426 11994
rect 23478 11942 23490 11994
rect 23542 11942 30662 11994
rect 30714 11942 30726 11994
rect 30778 11942 30790 11994
rect 30842 11942 30854 11994
rect 30906 11942 30918 11994
rect 30970 11942 30976 11994
rect 1104 11920 30976 11942
rect 7650 11880 7656 11892
rect 5920 11852 7656 11880
rect 4430 11772 4436 11824
rect 4488 11772 4494 11824
rect 5718 11812 5724 11824
rect 5658 11784 5724 11812
rect 5718 11772 5724 11784
rect 5776 11772 5782 11824
rect 4154 11704 4160 11756
rect 4212 11704 4218 11756
rect 4982 11636 4988 11688
rect 5040 11676 5046 11688
rect 5920 11685 5948 11852
rect 7650 11840 7656 11852
rect 7708 11840 7714 11892
rect 7926 11840 7932 11892
rect 7984 11880 7990 11892
rect 8665 11883 8723 11889
rect 8665 11880 8677 11883
rect 7984 11852 8677 11880
rect 7984 11840 7990 11852
rect 8665 11849 8677 11852
rect 8711 11849 8723 11883
rect 8665 11843 8723 11849
rect 12618 11840 12624 11892
rect 12676 11880 12682 11892
rect 12802 11880 12808 11892
rect 12676 11852 12808 11880
rect 12676 11840 12682 11852
rect 12802 11840 12808 11852
rect 12860 11880 12866 11892
rect 12989 11883 13047 11889
rect 12989 11880 13001 11883
rect 12860 11852 13001 11880
rect 12860 11840 12866 11852
rect 12989 11849 13001 11852
rect 13035 11849 13047 11883
rect 12989 11843 13047 11849
rect 7092 11747 7150 11753
rect 7092 11713 7104 11747
rect 7138 11744 7150 11747
rect 7558 11744 7564 11756
rect 7138 11716 7564 11744
rect 7138 11713 7150 11716
rect 7092 11707 7150 11713
rect 7558 11704 7564 11716
rect 7616 11704 7622 11756
rect 7834 11704 7840 11756
rect 7892 11744 7898 11756
rect 8665 11747 8723 11753
rect 8665 11744 8677 11747
rect 7892 11716 8677 11744
rect 7892 11704 7898 11716
rect 8665 11713 8677 11716
rect 8711 11713 8723 11747
rect 8665 11707 8723 11713
rect 8849 11747 8907 11753
rect 8849 11713 8861 11747
rect 8895 11713 8907 11747
rect 8849 11707 8907 11713
rect 5905 11679 5963 11685
rect 5905 11676 5917 11679
rect 5040 11648 5917 11676
rect 5040 11636 5046 11648
rect 5905 11645 5917 11648
rect 5951 11645 5963 11679
rect 5905 11639 5963 11645
rect 6822 11636 6828 11688
rect 6880 11636 6886 11688
rect 8018 11568 8024 11620
rect 8076 11608 8082 11620
rect 8205 11611 8263 11617
rect 8205 11608 8217 11611
rect 8076 11580 8217 11608
rect 8076 11568 8082 11580
rect 8205 11577 8217 11580
rect 8251 11608 8263 11611
rect 8864 11608 8892 11707
rect 8938 11704 8944 11756
rect 8996 11744 9002 11756
rect 9585 11747 9643 11753
rect 9585 11744 9597 11747
rect 8996 11716 9597 11744
rect 8996 11704 9002 11716
rect 9585 11713 9597 11716
rect 9631 11713 9643 11747
rect 9585 11707 9643 11713
rect 9674 11704 9680 11756
rect 9732 11744 9738 11756
rect 10413 11747 10471 11753
rect 10413 11744 10425 11747
rect 9732 11716 10425 11744
rect 9732 11704 9738 11716
rect 10413 11713 10425 11716
rect 10459 11713 10471 11747
rect 10413 11707 10471 11713
rect 10686 11704 10692 11756
rect 10744 11704 10750 11756
rect 13004 11744 13032 11843
rect 18230 11772 18236 11824
rect 18288 11812 18294 11824
rect 23661 11815 23719 11821
rect 18288 11784 19012 11812
rect 18288 11772 18294 11784
rect 17770 11744 17776 11756
rect 13004 11716 17776 11744
rect 17770 11704 17776 11716
rect 17828 11704 17834 11756
rect 18506 11704 18512 11756
rect 18564 11704 18570 11756
rect 18984 11753 19012 11784
rect 23661 11781 23673 11815
rect 23707 11812 23719 11815
rect 23750 11812 23756 11824
rect 23707 11784 23756 11812
rect 23707 11781 23719 11784
rect 23661 11775 23719 11781
rect 23750 11772 23756 11784
rect 23808 11772 23814 11824
rect 23020 11756 23072 11762
rect 18969 11747 19027 11753
rect 18969 11713 18981 11747
rect 19015 11713 19027 11747
rect 18969 11707 19027 11713
rect 19886 11704 19892 11756
rect 19944 11744 19950 11756
rect 20438 11744 20444 11756
rect 19944 11716 20444 11744
rect 19944 11704 19950 11716
rect 20438 11704 20444 11716
rect 20496 11744 20502 11756
rect 20717 11747 20775 11753
rect 20717 11744 20729 11747
rect 20496 11716 20729 11744
rect 20496 11704 20502 11716
rect 20717 11713 20729 11716
rect 20763 11713 20775 11747
rect 20717 11707 20775 11713
rect 22189 11747 22247 11753
rect 22189 11713 22201 11747
rect 22235 11713 22247 11747
rect 22189 11707 22247 11713
rect 9490 11636 9496 11688
rect 9548 11636 9554 11688
rect 9953 11679 10011 11685
rect 9953 11645 9965 11679
rect 9999 11676 10011 11679
rect 10505 11679 10563 11685
rect 10505 11676 10517 11679
rect 9999 11648 10517 11676
rect 9999 11645 10011 11648
rect 9953 11639 10011 11645
rect 10505 11645 10517 11648
rect 10551 11645 10563 11679
rect 10505 11639 10563 11645
rect 13078 11636 13084 11688
rect 13136 11636 13142 11688
rect 13262 11636 13268 11688
rect 13320 11636 13326 11688
rect 17862 11636 17868 11688
rect 17920 11636 17926 11688
rect 8251 11580 8892 11608
rect 22204 11608 22232 11707
rect 22922 11704 22928 11756
rect 22980 11704 22986 11756
rect 23020 11698 23072 11704
rect 23106 11608 23112 11620
rect 22204 11580 23112 11608
rect 8251 11577 8263 11580
rect 8205 11571 8263 11577
rect 23106 11568 23112 11580
rect 23164 11568 23170 11620
rect 10410 11500 10416 11552
rect 10468 11500 10474 11552
rect 10873 11543 10931 11549
rect 10873 11509 10885 11543
rect 10919 11540 10931 11543
rect 11974 11540 11980 11552
rect 10919 11512 11980 11540
rect 10919 11509 10931 11512
rect 10873 11503 10931 11509
rect 11974 11500 11980 11512
rect 12032 11500 12038 11552
rect 12618 11500 12624 11552
rect 12676 11500 12682 11552
rect 19061 11543 19119 11549
rect 19061 11509 19073 11543
rect 19107 11540 19119 11543
rect 19426 11540 19432 11552
rect 19107 11512 19432 11540
rect 19107 11509 19119 11512
rect 19061 11503 19119 11509
rect 19426 11500 19432 11512
rect 19484 11500 19490 11552
rect 19797 11543 19855 11549
rect 19797 11509 19809 11543
rect 19843 11540 19855 11543
rect 19886 11540 19892 11552
rect 19843 11512 19892 11540
rect 19843 11509 19855 11512
rect 19797 11503 19855 11509
rect 19886 11500 19892 11512
rect 19944 11500 19950 11552
rect 20809 11543 20867 11549
rect 20809 11509 20821 11543
rect 20855 11540 20867 11543
rect 21726 11540 21732 11552
rect 20855 11512 21732 11540
rect 20855 11509 20867 11512
rect 20809 11503 20867 11509
rect 21726 11500 21732 11512
rect 21784 11500 21790 11552
rect 22002 11500 22008 11552
rect 22060 11540 22066 11552
rect 22097 11543 22155 11549
rect 22097 11540 22109 11543
rect 22060 11512 22109 11540
rect 22060 11500 22066 11512
rect 22097 11509 22109 11512
rect 22143 11509 22155 11543
rect 22097 11503 22155 11509
rect 1104 11450 30820 11472
rect 1104 11398 4664 11450
rect 4716 11398 4728 11450
rect 4780 11398 4792 11450
rect 4844 11398 4856 11450
rect 4908 11398 4920 11450
rect 4972 11398 12092 11450
rect 12144 11398 12156 11450
rect 12208 11398 12220 11450
rect 12272 11398 12284 11450
rect 12336 11398 12348 11450
rect 12400 11398 19520 11450
rect 19572 11398 19584 11450
rect 19636 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 26948 11450
rect 27000 11398 27012 11450
rect 27064 11398 27076 11450
rect 27128 11398 27140 11450
rect 27192 11398 27204 11450
rect 27256 11398 30820 11450
rect 1104 11376 30820 11398
rect 7558 11296 7564 11348
rect 7616 11296 7622 11348
rect 12066 11296 12072 11348
rect 12124 11336 12130 11348
rect 13078 11336 13084 11348
rect 12124 11308 13084 11336
rect 12124 11296 12130 11308
rect 13078 11296 13084 11308
rect 13136 11336 13142 11348
rect 13449 11339 13507 11345
rect 13449 11336 13461 11339
rect 13136 11308 13461 11336
rect 13136 11296 13142 11308
rect 13449 11305 13461 11308
rect 13495 11305 13507 11339
rect 13449 11299 13507 11305
rect 18230 11296 18236 11348
rect 18288 11336 18294 11348
rect 18417 11339 18475 11345
rect 18417 11336 18429 11339
rect 18288 11308 18429 11336
rect 18288 11296 18294 11308
rect 18417 11305 18429 11308
rect 18463 11305 18475 11339
rect 18417 11299 18475 11305
rect 20438 11296 20444 11348
rect 20496 11336 20502 11348
rect 21177 11339 21235 11345
rect 21177 11336 21189 11339
rect 20496 11308 21189 11336
rect 20496 11296 20502 11308
rect 21177 11305 21189 11308
rect 21223 11305 21235 11339
rect 21177 11299 21235 11305
rect 23106 11296 23112 11348
rect 23164 11336 23170 11348
rect 23477 11339 23535 11345
rect 23477 11336 23489 11339
rect 23164 11308 23489 11336
rect 23164 11296 23170 11308
rect 23477 11305 23489 11308
rect 23523 11305 23535 11339
rect 23477 11299 23535 11305
rect 28994 11228 29000 11280
rect 29052 11228 29058 11280
rect 30282 11228 30288 11280
rect 30340 11228 30346 11280
rect 5166 11200 5172 11212
rect 4264 11172 5172 11200
rect 4264 11144 4292 11172
rect 5166 11160 5172 11172
rect 5224 11160 5230 11212
rect 5258 11160 5264 11212
rect 5316 11200 5322 11212
rect 5534 11200 5540 11212
rect 5316 11172 5540 11200
rect 5316 11160 5322 11172
rect 5534 11160 5540 11172
rect 5592 11160 5598 11212
rect 5718 11160 5724 11212
rect 5776 11160 5782 11212
rect 8018 11160 8024 11212
rect 8076 11160 8082 11212
rect 8202 11160 8208 11212
rect 8260 11200 8266 11212
rect 9122 11200 9128 11212
rect 8260 11172 9128 11200
rect 8260 11160 8266 11172
rect 9122 11160 9128 11172
rect 9180 11160 9186 11212
rect 11882 11160 11888 11212
rect 11940 11200 11946 11212
rect 12069 11203 12127 11209
rect 12069 11200 12081 11203
rect 11940 11172 12081 11200
rect 11940 11160 11946 11172
rect 12069 11169 12081 11172
rect 12115 11169 12127 11203
rect 12069 11163 12127 11169
rect 16117 11203 16175 11209
rect 16117 11169 16129 11203
rect 16163 11200 16175 11203
rect 16669 11203 16727 11209
rect 16669 11200 16681 11203
rect 16163 11172 16681 11200
rect 16163 11169 16175 11172
rect 16117 11163 16175 11169
rect 16669 11169 16681 11172
rect 16715 11169 16727 11203
rect 16669 11163 16727 11169
rect 16945 11203 17003 11209
rect 16945 11169 16957 11203
rect 16991 11200 17003 11203
rect 17310 11200 17316 11212
rect 16991 11172 17316 11200
rect 16991 11169 17003 11172
rect 16945 11163 17003 11169
rect 17310 11160 17316 11172
rect 17368 11160 17374 11212
rect 19426 11160 19432 11212
rect 19484 11160 19490 11212
rect 19705 11203 19763 11209
rect 19705 11169 19717 11203
rect 19751 11200 19763 11203
rect 19794 11200 19800 11212
rect 19751 11172 19800 11200
rect 19751 11169 19763 11172
rect 19705 11163 19763 11169
rect 19794 11160 19800 11172
rect 19852 11160 19858 11212
rect 21726 11160 21732 11212
rect 21784 11160 21790 11212
rect 22002 11160 22008 11212
rect 22060 11160 22066 11212
rect 23658 11160 23664 11212
rect 23716 11200 23722 11212
rect 24762 11200 24768 11212
rect 23716 11172 24768 11200
rect 23716 11160 23722 11172
rect 24762 11160 24768 11172
rect 24820 11200 24826 11212
rect 24820 11172 24900 11200
rect 24820 11160 24826 11172
rect 4246 11092 4252 11144
rect 4304 11092 4310 11144
rect 5077 11135 5135 11141
rect 5077 11101 5089 11135
rect 5123 11132 5135 11135
rect 5442 11132 5448 11144
rect 5123 11104 5448 11132
rect 5123 11101 5135 11104
rect 5077 11095 5135 11101
rect 5442 11092 5448 11104
rect 5500 11132 5506 11144
rect 5626 11132 5632 11144
rect 5500 11104 5632 11132
rect 5500 11092 5506 11104
rect 5626 11092 5632 11104
rect 5684 11092 5690 11144
rect 9858 11092 9864 11144
rect 9916 11092 9922 11144
rect 12336 11135 12394 11141
rect 12336 11101 12348 11135
rect 12382 11132 12394 11135
rect 12618 11132 12624 11144
rect 12382 11104 12624 11132
rect 12382 11101 12394 11104
rect 12336 11095 12394 11101
rect 12618 11092 12624 11104
rect 12676 11092 12682 11144
rect 16209 11135 16267 11141
rect 16209 11101 16221 11135
rect 16255 11101 16267 11135
rect 16209 11095 16267 11101
rect 4157 11067 4215 11073
rect 4157 11033 4169 11067
rect 4203 11064 4215 11067
rect 5718 11064 5724 11076
rect 4203 11036 5724 11064
rect 4203 11033 4215 11036
rect 4157 11027 4215 11033
rect 5718 11024 5724 11036
rect 5776 11024 5782 11076
rect 7929 11067 7987 11073
rect 7929 11033 7941 11067
rect 7975 11064 7987 11067
rect 14918 11064 14924 11076
rect 7975 11036 14924 11064
rect 7975 11033 7987 11036
rect 7929 11027 7987 11033
rect 14918 11024 14924 11036
rect 14976 11024 14982 11076
rect 9953 10999 10011 11005
rect 9953 10965 9965 10999
rect 9999 10996 10011 10999
rect 10042 10996 10048 11008
rect 9999 10968 10048 10996
rect 9999 10965 10011 10968
rect 9953 10959 10011 10965
rect 10042 10956 10048 10968
rect 10100 10956 10106 11008
rect 16224 10996 16252 11095
rect 23106 11092 23112 11144
rect 23164 11092 23170 11144
rect 24670 11092 24676 11144
rect 24728 11092 24734 11144
rect 24872 11141 24900 11172
rect 25406 11160 25412 11212
rect 25464 11200 25470 11212
rect 25869 11203 25927 11209
rect 25869 11200 25881 11203
rect 25464 11172 25881 11200
rect 25464 11160 25470 11172
rect 25869 11169 25881 11172
rect 25915 11169 25927 11203
rect 25869 11163 25927 11169
rect 29181 11203 29239 11209
rect 29181 11169 29193 11203
rect 29227 11169 29239 11203
rect 29181 11163 29239 11169
rect 24857 11135 24915 11141
rect 24857 11101 24869 11135
rect 24903 11101 24915 11135
rect 24857 11095 24915 11101
rect 25682 11092 25688 11144
rect 25740 11092 25746 11144
rect 29196 11132 29224 11163
rect 29822 11160 29828 11212
rect 29880 11160 29886 11212
rect 29917 11135 29975 11141
rect 29917 11132 29929 11135
rect 29196 11104 29929 11132
rect 29917 11101 29929 11104
rect 29963 11101 29975 11135
rect 29917 11095 29975 11101
rect 17954 11024 17960 11076
rect 18012 11024 18018 11076
rect 20714 11024 20720 11076
rect 20772 11024 20778 11076
rect 25777 11067 25835 11073
rect 25777 11033 25789 11067
rect 25823 11064 25835 11067
rect 26510 11064 26516 11076
rect 25823 11036 26516 11064
rect 25823 11033 25835 11036
rect 25777 11027 25835 11033
rect 26510 11024 26516 11036
rect 26568 11024 26574 11076
rect 28718 11024 28724 11076
rect 28776 11024 28782 11076
rect 16298 10996 16304 11008
rect 16224 10968 16304 10996
rect 16298 10956 16304 10968
rect 16356 10996 16362 11008
rect 18598 10996 18604 11008
rect 16356 10968 18604 10996
rect 16356 10956 16362 10968
rect 18598 10956 18604 10968
rect 18656 10956 18662 11008
rect 24854 10956 24860 11008
rect 24912 10956 24918 11008
rect 25314 10956 25320 11008
rect 25372 10956 25378 11008
rect 1104 10906 30976 10928
rect 1104 10854 8378 10906
rect 8430 10854 8442 10906
rect 8494 10854 8506 10906
rect 8558 10854 8570 10906
rect 8622 10854 8634 10906
rect 8686 10854 15806 10906
rect 15858 10854 15870 10906
rect 15922 10854 15934 10906
rect 15986 10854 15998 10906
rect 16050 10854 16062 10906
rect 16114 10854 23234 10906
rect 23286 10854 23298 10906
rect 23350 10854 23362 10906
rect 23414 10854 23426 10906
rect 23478 10854 23490 10906
rect 23542 10854 30662 10906
rect 30714 10854 30726 10906
rect 30778 10854 30790 10906
rect 30842 10854 30854 10906
rect 30906 10854 30918 10906
rect 30970 10854 30976 10906
rect 1104 10832 30976 10854
rect 4246 10752 4252 10804
rect 4304 10752 4310 10804
rect 7561 10795 7619 10801
rect 7561 10761 7573 10795
rect 7607 10792 7619 10795
rect 8110 10792 8116 10804
rect 7607 10764 8116 10792
rect 7607 10761 7619 10764
rect 7561 10755 7619 10761
rect 8110 10752 8116 10764
rect 8168 10752 8174 10804
rect 12434 10752 12440 10804
rect 12492 10792 12498 10804
rect 12621 10795 12679 10801
rect 12621 10792 12633 10795
rect 12492 10764 12633 10792
rect 12492 10752 12498 10764
rect 12621 10761 12633 10764
rect 12667 10761 12679 10795
rect 12621 10755 12679 10761
rect 18598 10752 18604 10804
rect 18656 10752 18662 10804
rect 24854 10752 24860 10804
rect 24912 10792 24918 10804
rect 28077 10795 28135 10801
rect 24912 10764 25452 10792
rect 24912 10752 24918 10764
rect 4982 10684 4988 10736
rect 5040 10684 5046 10736
rect 5718 10684 5724 10736
rect 5776 10684 5782 10736
rect 7745 10727 7803 10733
rect 7745 10693 7757 10727
rect 7791 10724 7803 10727
rect 7834 10724 7840 10736
rect 7791 10696 7840 10724
rect 7791 10693 7803 10696
rect 7745 10687 7803 10693
rect 7834 10684 7840 10696
rect 7892 10684 7898 10736
rect 7929 10727 7987 10733
rect 7929 10693 7941 10727
rect 7975 10724 7987 10727
rect 8018 10724 8024 10736
rect 7975 10696 8024 10724
rect 7975 10693 7987 10696
rect 7929 10687 7987 10693
rect 8018 10684 8024 10696
rect 8076 10684 8082 10736
rect 10505 10727 10563 10733
rect 10505 10693 10517 10727
rect 10551 10724 10563 10727
rect 11514 10724 11520 10736
rect 10551 10696 11520 10724
rect 10551 10693 10563 10696
rect 10505 10687 10563 10693
rect 11514 10684 11520 10696
rect 11572 10684 11578 10736
rect 11974 10684 11980 10736
rect 12032 10724 12038 10736
rect 12161 10727 12219 10733
rect 12161 10724 12173 10727
rect 12032 10696 12173 10724
rect 12032 10684 12038 10696
rect 12161 10693 12173 10696
rect 12207 10693 12219 10727
rect 12161 10687 12219 10693
rect 16209 10727 16267 10733
rect 16209 10693 16221 10727
rect 16255 10724 16267 10727
rect 17129 10727 17187 10733
rect 17129 10724 17141 10727
rect 16255 10696 17141 10724
rect 16255 10693 16267 10696
rect 16209 10687 16267 10693
rect 17129 10693 17141 10696
rect 17175 10693 17187 10727
rect 17129 10687 17187 10693
rect 18138 10684 18144 10736
rect 18196 10684 18202 10736
rect 20349 10727 20407 10733
rect 20349 10693 20361 10727
rect 20395 10724 20407 10727
rect 20714 10724 20720 10736
rect 20395 10696 20720 10724
rect 20395 10693 20407 10696
rect 20349 10687 20407 10693
rect 20714 10684 20720 10696
rect 20772 10684 20778 10736
rect 23106 10684 23112 10736
rect 23164 10684 23170 10736
rect 25041 10727 25099 10733
rect 25041 10693 25053 10727
rect 25087 10724 25099 10727
rect 25314 10724 25320 10736
rect 25087 10696 25320 10724
rect 25087 10693 25099 10696
rect 25041 10687 25099 10693
rect 25314 10684 25320 10696
rect 25372 10684 25378 10736
rect 25424 10724 25452 10764
rect 28077 10761 28089 10795
rect 28123 10761 28135 10795
rect 28077 10755 28135 10761
rect 29733 10795 29791 10801
rect 29733 10761 29745 10795
rect 29779 10792 29791 10795
rect 29822 10792 29828 10804
rect 29779 10764 29828 10792
rect 29779 10761 29791 10764
rect 29733 10755 29791 10761
rect 25424 10696 25530 10724
rect 27430 10684 27436 10736
rect 27488 10724 27494 10736
rect 27709 10727 27767 10733
rect 27709 10724 27721 10727
rect 27488 10696 27721 10724
rect 27488 10684 27494 10696
rect 27709 10693 27721 10696
rect 27755 10693 27767 10727
rect 27709 10687 27767 10693
rect 27801 10727 27859 10733
rect 27801 10693 27813 10727
rect 27847 10724 27859 10727
rect 27982 10724 27988 10736
rect 27847 10696 27988 10724
rect 27847 10693 27859 10696
rect 27801 10687 27859 10693
rect 27982 10684 27988 10696
rect 28040 10684 28046 10736
rect 28092 10724 28120 10755
rect 29822 10752 29828 10764
rect 29880 10752 29886 10804
rect 28994 10724 29000 10736
rect 28092 10696 29000 10724
rect 19984 10668 20036 10674
rect 6733 10659 6791 10665
rect 6733 10625 6745 10659
rect 6779 10656 6791 10659
rect 6779 10628 6914 10656
rect 6779 10625 6791 10628
rect 6733 10619 6791 10625
rect 5997 10591 6055 10597
rect 5997 10557 6009 10591
rect 6043 10588 6055 10591
rect 6641 10591 6699 10597
rect 6641 10588 6653 10591
rect 6043 10560 6653 10588
rect 6043 10557 6055 10560
rect 5997 10551 6055 10557
rect 6641 10557 6653 10560
rect 6687 10557 6699 10591
rect 6886 10588 6914 10628
rect 11146 10616 11152 10668
rect 11204 10616 11210 10668
rect 12437 10659 12495 10665
rect 12437 10625 12449 10659
rect 12483 10656 12495 10659
rect 12894 10656 12900 10668
rect 12483 10628 12900 10656
rect 12483 10625 12495 10628
rect 12437 10619 12495 10625
rect 12894 10616 12900 10628
rect 12952 10616 12958 10668
rect 13440 10659 13498 10665
rect 13440 10625 13452 10659
rect 13486 10656 13498 10659
rect 14274 10656 14280 10668
rect 13486 10628 14280 10656
rect 13486 10625 13498 10628
rect 13440 10619 13498 10625
rect 14274 10616 14280 10628
rect 14332 10616 14338 10668
rect 16298 10616 16304 10668
rect 16356 10616 16362 10668
rect 16758 10616 16764 10668
rect 16816 10656 16822 10668
rect 16853 10659 16911 10665
rect 16853 10656 16865 10659
rect 16816 10628 16865 10656
rect 16816 10616 16822 10628
rect 16853 10625 16865 10628
rect 16899 10625 16911 10659
rect 16853 10619 16911 10625
rect 23014 10656 23020 10668
rect 22770 10628 23020 10656
rect 23014 10616 23020 10628
rect 23072 10616 23078 10668
rect 24762 10616 24768 10668
rect 24820 10616 24826 10668
rect 27525 10659 27583 10665
rect 27525 10625 27537 10659
rect 27571 10656 27583 10659
rect 27893 10659 27951 10665
rect 27571 10628 27752 10656
rect 27571 10625 27583 10628
rect 27525 10619 27583 10625
rect 19984 10610 20036 10616
rect 27724 10600 27752 10628
rect 27893 10625 27905 10659
rect 27939 10656 27951 10659
rect 28166 10656 28172 10668
rect 27939 10628 28172 10656
rect 27939 10625 27951 10628
rect 27893 10619 27951 10625
rect 28166 10616 28172 10628
rect 28224 10616 28230 10668
rect 28644 10665 28672 10696
rect 28994 10684 29000 10696
rect 29052 10684 29058 10736
rect 29089 10727 29147 10733
rect 29089 10693 29101 10727
rect 29135 10724 29147 10727
rect 29914 10724 29920 10736
rect 29135 10696 29920 10724
rect 29135 10693 29147 10696
rect 29089 10687 29147 10693
rect 29914 10684 29920 10696
rect 29972 10684 29978 10736
rect 28629 10659 28687 10665
rect 28629 10625 28641 10659
rect 28675 10625 28687 10659
rect 28629 10619 28687 10625
rect 28718 10616 28724 10668
rect 28776 10616 28782 10668
rect 28813 10659 28871 10665
rect 28813 10625 28825 10659
rect 28859 10625 28871 10659
rect 28813 10619 28871 10625
rect 9858 10588 9864 10600
rect 6886 10560 9864 10588
rect 6641 10551 6699 10557
rect 9858 10548 9864 10560
rect 9916 10548 9922 10600
rect 12345 10591 12403 10597
rect 12345 10557 12357 10591
rect 12391 10588 12403 10591
rect 12526 10588 12532 10600
rect 12391 10560 12532 10588
rect 12391 10557 12403 10560
rect 12345 10551 12403 10557
rect 12526 10548 12532 10560
rect 12584 10548 12590 10600
rect 12710 10548 12716 10600
rect 12768 10588 12774 10600
rect 13173 10591 13231 10597
rect 13173 10588 13185 10591
rect 12768 10560 13185 10588
rect 12768 10548 12774 10560
rect 13173 10557 13185 10560
rect 13219 10557 13231 10591
rect 13173 10551 13231 10557
rect 17862 10548 17868 10600
rect 17920 10588 17926 10600
rect 19521 10591 19579 10597
rect 19521 10588 19533 10591
rect 17920 10560 19533 10588
rect 17920 10548 17926 10560
rect 19521 10557 19533 10560
rect 19567 10557 19579 10591
rect 19521 10551 19579 10557
rect 22281 10591 22339 10597
rect 22281 10557 22293 10591
rect 22327 10588 22339 10591
rect 22922 10588 22928 10600
rect 22327 10560 22928 10588
rect 22327 10557 22339 10560
rect 22281 10551 22339 10557
rect 19536 10520 19564 10551
rect 22296 10520 22324 10551
rect 22922 10548 22928 10560
rect 22980 10548 22986 10600
rect 26510 10548 26516 10600
rect 26568 10588 26574 10600
rect 27706 10588 27712 10600
rect 26568 10560 27712 10588
rect 26568 10548 26574 10560
rect 27706 10548 27712 10560
rect 27764 10548 27770 10600
rect 28828 10588 28856 10619
rect 28902 10616 28908 10668
rect 28960 10656 28966 10668
rect 29641 10659 29699 10665
rect 29641 10656 29653 10659
rect 28960 10628 29653 10656
rect 28960 10616 28966 10628
rect 29641 10625 29653 10628
rect 29687 10625 29699 10659
rect 29641 10619 29699 10625
rect 29825 10659 29883 10665
rect 29825 10625 29837 10659
rect 29871 10625 29883 10659
rect 29825 10619 29883 10625
rect 29730 10588 29736 10600
rect 28828 10560 29736 10588
rect 29730 10548 29736 10560
rect 29788 10588 29794 10600
rect 29840 10588 29868 10619
rect 29788 10560 29868 10588
rect 29788 10548 29794 10560
rect 19536 10492 22324 10520
rect 9214 10412 9220 10464
rect 9272 10412 9278 10464
rect 9766 10412 9772 10464
rect 9824 10452 9830 10464
rect 11057 10455 11115 10461
rect 11057 10452 11069 10455
rect 9824 10424 11069 10452
rect 9824 10412 9830 10424
rect 11057 10421 11069 10424
rect 11103 10421 11115 10455
rect 11057 10415 11115 10421
rect 12434 10412 12440 10464
rect 12492 10412 12498 10464
rect 14550 10412 14556 10464
rect 14608 10412 14614 10464
rect 1104 10362 30820 10384
rect 1104 10310 4664 10362
rect 4716 10310 4728 10362
rect 4780 10310 4792 10362
rect 4844 10310 4856 10362
rect 4908 10310 4920 10362
rect 4972 10310 12092 10362
rect 12144 10310 12156 10362
rect 12208 10310 12220 10362
rect 12272 10310 12284 10362
rect 12336 10310 12348 10362
rect 12400 10310 19520 10362
rect 19572 10310 19584 10362
rect 19636 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 26948 10362
rect 27000 10310 27012 10362
rect 27064 10310 27076 10362
rect 27128 10310 27140 10362
rect 27192 10310 27204 10362
rect 27256 10310 30820 10362
rect 1104 10288 30820 10310
rect 5534 10208 5540 10260
rect 5592 10208 5598 10260
rect 9858 10208 9864 10260
rect 9916 10248 9922 10260
rect 11517 10251 11575 10257
rect 11517 10248 11529 10251
rect 9916 10220 11529 10248
rect 9916 10208 9922 10220
rect 11517 10217 11529 10220
rect 11563 10248 11575 10251
rect 12066 10248 12072 10260
rect 11563 10220 12072 10248
rect 11563 10217 11575 10220
rect 11517 10211 11575 10217
rect 12066 10208 12072 10220
rect 12124 10208 12130 10260
rect 12526 10208 12532 10260
rect 12584 10208 12590 10260
rect 14274 10208 14280 10260
rect 14332 10208 14338 10260
rect 17862 10208 17868 10260
rect 17920 10208 17926 10260
rect 19978 10208 19984 10260
rect 20036 10248 20042 10260
rect 21269 10251 21327 10257
rect 21269 10248 21281 10251
rect 20036 10220 21281 10248
rect 20036 10208 20042 10220
rect 21269 10217 21281 10220
rect 21315 10248 21327 10251
rect 23014 10248 23020 10260
rect 21315 10220 23020 10248
rect 21315 10217 21327 10220
rect 21269 10211 21327 10217
rect 23014 10208 23020 10220
rect 23072 10208 23078 10260
rect 28445 10251 28503 10257
rect 28445 10217 28457 10251
rect 28491 10248 28503 10251
rect 28718 10248 28724 10260
rect 28491 10220 28724 10248
rect 28491 10217 28503 10220
rect 28445 10211 28503 10217
rect 28718 10208 28724 10220
rect 28776 10208 28782 10260
rect 29730 10208 29736 10260
rect 29788 10208 29794 10260
rect 17880 10180 17908 10208
rect 17144 10152 17908 10180
rect 8202 10072 8208 10124
rect 8260 10072 8266 10124
rect 9766 10072 9772 10124
rect 9824 10072 9830 10124
rect 10042 10072 10048 10124
rect 10100 10072 10106 10124
rect 12989 10115 13047 10121
rect 12989 10081 13001 10115
rect 13035 10112 13047 10115
rect 14550 10112 14556 10124
rect 13035 10084 14556 10112
rect 13035 10081 13047 10084
rect 12989 10075 13047 10081
rect 14550 10072 14556 10084
rect 14608 10112 14614 10124
rect 14737 10115 14795 10121
rect 14737 10112 14749 10115
rect 14608 10084 14749 10112
rect 14608 10072 14614 10084
rect 14737 10081 14749 10084
rect 14783 10081 14795 10115
rect 14737 10075 14795 10081
rect 14921 10115 14979 10121
rect 14921 10081 14933 10115
rect 14967 10112 14979 10115
rect 15102 10112 15108 10124
rect 14967 10084 15108 10112
rect 14967 10081 14979 10084
rect 14921 10075 14979 10081
rect 15102 10072 15108 10084
rect 15160 10072 15166 10124
rect 17144 10121 17172 10152
rect 17129 10115 17187 10121
rect 17129 10081 17141 10115
rect 17175 10081 17187 10115
rect 17129 10075 17187 10081
rect 17865 10115 17923 10121
rect 17865 10081 17877 10115
rect 17911 10112 17923 10115
rect 17954 10112 17960 10124
rect 17911 10084 17960 10112
rect 17911 10081 17923 10084
rect 17865 10075 17923 10081
rect 17954 10072 17960 10084
rect 18012 10072 18018 10124
rect 17592 10056 17644 10062
rect 8021 10047 8079 10053
rect 8021 10013 8033 10047
rect 8067 10044 8079 10047
rect 8067 10016 9812 10044
rect 8067 10013 8079 10016
rect 8021 10007 8079 10013
rect 7009 9979 7067 9985
rect 7009 9945 7021 9979
rect 7055 9976 7067 9979
rect 9214 9976 9220 9988
rect 7055 9948 9220 9976
rect 7055 9945 7067 9948
rect 7009 9939 7067 9945
rect 9214 9936 9220 9948
rect 9272 9936 9278 9988
rect 9784 9976 9812 10016
rect 11330 10004 11336 10056
rect 11388 10044 11394 10056
rect 12526 10044 12532 10056
rect 11388 10016 12532 10044
rect 11388 10004 11394 10016
rect 12526 10004 12532 10016
rect 12584 10044 12590 10056
rect 12897 10047 12955 10053
rect 12897 10044 12909 10047
rect 12584 10016 12909 10044
rect 12584 10004 12590 10016
rect 12897 10013 12909 10016
rect 12943 10013 12955 10047
rect 12897 10007 12955 10013
rect 14642 10004 14648 10056
rect 14700 10004 14706 10056
rect 19996 10044 20024 10208
rect 29917 10183 29975 10189
rect 29917 10149 29929 10183
rect 29963 10180 29975 10183
rect 30006 10180 30012 10192
rect 29963 10152 30012 10180
rect 29963 10149 29975 10152
rect 29917 10143 29975 10149
rect 30006 10140 30012 10152
rect 30064 10140 30070 10192
rect 25406 10072 25412 10124
rect 25464 10112 25470 10124
rect 25501 10115 25559 10121
rect 25501 10112 25513 10115
rect 25464 10084 25513 10112
rect 25464 10072 25470 10084
rect 25501 10081 25513 10084
rect 25547 10081 25559 10115
rect 25501 10075 25559 10081
rect 17644 10016 20024 10044
rect 22557 10047 22615 10053
rect 22557 10013 22569 10047
rect 22603 10044 22615 10047
rect 24578 10044 24584 10056
rect 22603 10016 24584 10044
rect 22603 10013 22615 10016
rect 22557 10007 22615 10013
rect 24578 10004 24584 10016
rect 24636 10004 24642 10056
rect 25038 10004 25044 10056
rect 25096 10044 25102 10056
rect 25317 10047 25375 10053
rect 25317 10044 25329 10047
rect 25096 10016 25329 10044
rect 25096 10004 25102 10016
rect 25317 10013 25329 10016
rect 25363 10013 25375 10047
rect 25317 10007 25375 10013
rect 27982 10004 27988 10056
rect 28040 10044 28046 10056
rect 28077 10047 28135 10053
rect 28077 10044 28089 10047
rect 28040 10016 28089 10044
rect 28040 10004 28046 10016
rect 28077 10013 28089 10016
rect 28123 10013 28135 10047
rect 28077 10007 28135 10013
rect 28166 10004 28172 10056
rect 28224 10044 28230 10056
rect 28905 10047 28963 10053
rect 28905 10044 28917 10047
rect 28224 10016 28917 10044
rect 28224 10004 28230 10016
rect 28905 10013 28917 10016
rect 28951 10013 28963 10047
rect 28905 10007 28963 10013
rect 17592 9998 17644 10004
rect 9784 9948 10456 9976
rect 7650 9868 7656 9920
rect 7708 9868 7714 9920
rect 8113 9911 8171 9917
rect 8113 9877 8125 9911
rect 8159 9908 8171 9911
rect 8294 9908 8300 9920
rect 8159 9880 8300 9908
rect 8159 9877 8171 9880
rect 8113 9871 8171 9877
rect 8294 9868 8300 9880
rect 8352 9868 8358 9920
rect 10428 9908 10456 9948
rect 11054 9936 11060 9988
rect 11112 9936 11118 9988
rect 27706 9936 27712 9988
rect 27764 9976 27770 9988
rect 27893 9979 27951 9985
rect 27893 9976 27905 9979
rect 27764 9948 27905 9976
rect 27764 9936 27770 9948
rect 27893 9945 27905 9948
rect 27939 9945 27951 9979
rect 28261 9979 28319 9985
rect 28261 9976 28273 9979
rect 27893 9939 27951 9945
rect 28000 9948 28273 9976
rect 12802 9908 12808 9920
rect 10428 9880 12808 9908
rect 12802 9868 12808 9880
rect 12860 9868 12866 9920
rect 24854 9868 24860 9920
rect 24912 9908 24918 9920
rect 24949 9911 25007 9917
rect 24949 9908 24961 9911
rect 24912 9880 24961 9908
rect 24912 9868 24918 9880
rect 24949 9877 24961 9880
rect 24995 9877 25007 9911
rect 24949 9871 25007 9877
rect 25409 9911 25467 9917
rect 25409 9877 25421 9911
rect 25455 9908 25467 9911
rect 26050 9908 26056 9920
rect 25455 9880 26056 9908
rect 25455 9877 25467 9880
rect 25409 9871 25467 9877
rect 26050 9868 26056 9880
rect 26108 9868 26114 9920
rect 27430 9868 27436 9920
rect 27488 9908 27494 9920
rect 28000 9908 28028 9948
rect 28261 9945 28273 9948
rect 28307 9945 28319 9979
rect 28261 9939 28319 9945
rect 30190 9936 30196 9988
rect 30248 9936 30254 9988
rect 27488 9880 28028 9908
rect 27488 9868 27494 9880
rect 28994 9868 29000 9920
rect 29052 9868 29058 9920
rect 1104 9818 30976 9840
rect 1104 9766 8378 9818
rect 8430 9766 8442 9818
rect 8494 9766 8506 9818
rect 8558 9766 8570 9818
rect 8622 9766 8634 9818
rect 8686 9766 15806 9818
rect 15858 9766 15870 9818
rect 15922 9766 15934 9818
rect 15986 9766 15998 9818
rect 16050 9766 16062 9818
rect 16114 9766 23234 9818
rect 23286 9766 23298 9818
rect 23350 9766 23362 9818
rect 23414 9766 23426 9818
rect 23478 9766 23490 9818
rect 23542 9766 30662 9818
rect 30714 9766 30726 9818
rect 30778 9766 30790 9818
rect 30842 9766 30854 9818
rect 30906 9766 30918 9818
rect 30970 9766 30976 9818
rect 1104 9744 30976 9766
rect 8294 9664 8300 9716
rect 8352 9704 8358 9716
rect 8386 9704 8392 9716
rect 8352 9676 8392 9704
rect 8352 9664 8358 9676
rect 8386 9664 8392 9676
rect 8444 9664 8450 9716
rect 14642 9664 14648 9716
rect 14700 9704 14706 9716
rect 24762 9704 24768 9716
rect 14700 9676 15240 9704
rect 14700 9664 14706 9676
rect 4801 9639 4859 9645
rect 4801 9605 4813 9639
rect 4847 9636 4859 9639
rect 4982 9636 4988 9648
rect 4847 9608 4988 9636
rect 4847 9605 4859 9608
rect 4801 9599 4859 9605
rect 4982 9596 4988 9608
rect 5040 9596 5046 9648
rect 7276 9639 7334 9645
rect 7276 9605 7288 9639
rect 7322 9636 7334 9639
rect 7650 9636 7656 9648
rect 7322 9608 7656 9636
rect 7322 9605 7334 9608
rect 7276 9599 7334 9605
rect 7650 9596 7656 9608
rect 7708 9596 7714 9648
rect 10965 9639 11023 9645
rect 10965 9605 10977 9639
rect 11011 9636 11023 9639
rect 11054 9636 11060 9648
rect 11011 9608 11060 9636
rect 11011 9605 11023 9608
rect 10965 9599 11023 9605
rect 11054 9596 11060 9608
rect 11112 9596 11118 9648
rect 15212 9645 15240 9676
rect 24412 9676 24768 9704
rect 15197 9639 15255 9645
rect 15197 9605 15209 9639
rect 15243 9605 15255 9639
rect 24412 9636 24440 9676
rect 24762 9664 24768 9676
rect 24820 9664 24826 9716
rect 26050 9664 26056 9716
rect 26108 9704 26114 9716
rect 27985 9707 28043 9713
rect 26108 9676 26234 9704
rect 26108 9664 26114 9676
rect 15197 9599 15255 9605
rect 24320 9608 24440 9636
rect 24581 9639 24639 9645
rect 17592 9580 17644 9586
rect 5626 9528 5632 9580
rect 5684 9528 5690 9580
rect 6822 9528 6828 9580
rect 6880 9568 6886 9580
rect 7009 9571 7067 9577
rect 7009 9568 7021 9571
rect 6880 9540 7021 9568
rect 6880 9528 6886 9540
rect 7009 9537 7021 9540
rect 7055 9537 7067 9571
rect 7009 9531 7067 9537
rect 8294 9528 8300 9580
rect 8352 9568 8358 9580
rect 9582 9568 9588 9580
rect 8352 9540 9588 9568
rect 8352 9528 8358 9540
rect 9582 9528 9588 9540
rect 9640 9568 9646 9580
rect 9953 9571 10011 9577
rect 9953 9568 9965 9571
rect 9640 9540 9965 9568
rect 9640 9528 9646 9540
rect 9953 9537 9965 9540
rect 9999 9537 10011 9571
rect 9953 9531 10011 9537
rect 10137 9571 10195 9577
rect 10137 9537 10149 9571
rect 10183 9537 10195 9571
rect 10137 9531 10195 9537
rect 5534 9460 5540 9512
rect 5592 9460 5598 9512
rect 9490 9460 9496 9512
rect 9548 9500 9554 9512
rect 10152 9500 10180 9531
rect 12066 9528 12072 9580
rect 12124 9528 12130 9580
rect 16390 9528 16396 9580
rect 16448 9568 16454 9580
rect 16574 9568 16580 9580
rect 16448 9540 16580 9568
rect 16448 9528 16454 9540
rect 16574 9528 16580 9540
rect 16632 9568 16638 9580
rect 16945 9571 17003 9577
rect 16945 9568 16957 9571
rect 16632 9540 16957 9568
rect 16632 9528 16638 9540
rect 16945 9537 16957 9540
rect 16991 9537 17003 9571
rect 16945 9531 17003 9537
rect 21910 9528 21916 9580
rect 21968 9568 21974 9580
rect 22005 9571 22063 9577
rect 22005 9568 22017 9571
rect 21968 9540 22017 9568
rect 21968 9528 21974 9540
rect 22005 9537 22017 9540
rect 22051 9537 22063 9571
rect 22005 9531 22063 9537
rect 22272 9571 22330 9577
rect 22272 9537 22284 9571
rect 22318 9568 22330 9571
rect 22830 9568 22836 9580
rect 22318 9540 22836 9568
rect 22318 9537 22330 9540
rect 22272 9531 22330 9537
rect 22830 9528 22836 9540
rect 22888 9528 22894 9580
rect 24320 9577 24348 9608
rect 24581 9605 24593 9639
rect 24627 9636 24639 9639
rect 24854 9636 24860 9648
rect 24627 9608 24860 9636
rect 24627 9605 24639 9608
rect 24581 9599 24639 9605
rect 24854 9596 24860 9608
rect 24912 9596 24918 9648
rect 25038 9596 25044 9648
rect 25096 9596 25102 9648
rect 26206 9636 26234 9676
rect 27985 9673 27997 9707
rect 28031 9704 28043 9707
rect 28166 9704 28172 9716
rect 28031 9676 28172 9704
rect 28031 9673 28043 9676
rect 27985 9667 28043 9673
rect 28166 9664 28172 9676
rect 28224 9664 28230 9716
rect 31018 9704 31024 9716
rect 30116 9676 31024 9704
rect 27890 9636 27896 9648
rect 26206 9608 27896 9636
rect 27890 9596 27896 9608
rect 27948 9596 27954 9648
rect 28994 9596 29000 9648
rect 29052 9636 29058 9648
rect 30116 9645 30144 9676
rect 31018 9664 31024 9676
rect 31076 9664 31082 9716
rect 29098 9639 29156 9645
rect 29098 9636 29110 9639
rect 29052 9608 29110 9636
rect 29052 9596 29058 9608
rect 29098 9605 29110 9608
rect 29144 9605 29156 9639
rect 29098 9599 29156 9605
rect 30101 9639 30159 9645
rect 30101 9605 30113 9639
rect 30147 9605 30159 9639
rect 30101 9599 30159 9605
rect 24305 9571 24363 9577
rect 24305 9537 24317 9571
rect 24351 9537 24363 9571
rect 24305 9531 24363 9537
rect 29822 9528 29828 9580
rect 29880 9528 29886 9580
rect 17592 9522 17644 9528
rect 9548 9472 10180 9500
rect 9548 9460 9554 9472
rect 11974 9460 11980 9512
rect 12032 9460 12038 9512
rect 12434 9460 12440 9512
rect 12492 9460 12498 9512
rect 14458 9460 14464 9512
rect 14516 9500 14522 9512
rect 15289 9503 15347 9509
rect 15289 9500 15301 9503
rect 14516 9472 15301 9500
rect 14516 9460 14522 9472
rect 15289 9469 15301 9472
rect 15335 9469 15347 9503
rect 15289 9463 15347 9469
rect 15378 9460 15384 9512
rect 15436 9460 15442 9512
rect 17865 9503 17923 9509
rect 17865 9469 17877 9503
rect 17911 9500 17923 9503
rect 18138 9500 18144 9512
rect 17911 9472 18144 9500
rect 17911 9469 17923 9472
rect 17865 9463 17923 9469
rect 18138 9460 18144 9472
rect 18196 9460 18202 9512
rect 29362 9460 29368 9512
rect 29420 9460 29426 9512
rect 14826 9324 14832 9376
rect 14884 9324 14890 9376
rect 23385 9367 23443 9373
rect 23385 9333 23397 9367
rect 23431 9364 23443 9367
rect 23842 9364 23848 9376
rect 23431 9336 23848 9364
rect 23431 9333 23443 9336
rect 23385 9327 23443 9333
rect 23842 9324 23848 9336
rect 23900 9324 23906 9376
rect 1104 9274 30820 9296
rect 1104 9222 4664 9274
rect 4716 9222 4728 9274
rect 4780 9222 4792 9274
rect 4844 9222 4856 9274
rect 4908 9222 4920 9274
rect 4972 9222 12092 9274
rect 12144 9222 12156 9274
rect 12208 9222 12220 9274
rect 12272 9222 12284 9274
rect 12336 9222 12348 9274
rect 12400 9222 19520 9274
rect 19572 9222 19584 9274
rect 19636 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 26948 9274
rect 27000 9222 27012 9274
rect 27064 9222 27076 9274
rect 27128 9222 27140 9274
rect 27192 9222 27204 9274
rect 27256 9222 30820 9274
rect 1104 9200 30820 9222
rect 9674 9120 9680 9172
rect 9732 9120 9738 9172
rect 14458 9120 14464 9172
rect 14516 9120 14522 9172
rect 22830 9120 22836 9172
rect 22888 9120 22894 9172
rect 24673 9163 24731 9169
rect 24673 9129 24685 9163
rect 24719 9160 24731 9163
rect 25038 9160 25044 9172
rect 24719 9132 25044 9160
rect 24719 9129 24731 9132
rect 24673 9123 24731 9129
rect 25038 9120 25044 9132
rect 25096 9120 25102 9172
rect 29822 9120 29828 9172
rect 29880 9120 29886 9172
rect 8386 8984 8392 9036
rect 8444 9024 8450 9036
rect 9217 9027 9275 9033
rect 9217 9024 9229 9027
rect 8444 8996 9229 9024
rect 8444 8984 8450 8996
rect 9217 8993 9229 8996
rect 9263 8993 9275 9027
rect 9217 8987 9275 8993
rect 30006 8984 30012 9036
rect 30064 8984 30070 9036
rect 5626 8916 5632 8968
rect 5684 8956 5690 8968
rect 7929 8959 7987 8965
rect 7929 8956 7941 8959
rect 5684 8928 7941 8956
rect 5684 8916 5690 8928
rect 7929 8925 7941 8928
rect 7975 8925 7987 8959
rect 7929 8919 7987 8925
rect 8205 8959 8263 8965
rect 8205 8925 8217 8959
rect 8251 8956 8263 8959
rect 8294 8956 8300 8968
rect 8251 8928 8300 8956
rect 8251 8925 8263 8928
rect 8205 8919 8263 8925
rect 7944 8888 7972 8919
rect 8294 8916 8300 8928
rect 8352 8916 8358 8968
rect 9306 8916 9312 8968
rect 9364 8916 9370 8968
rect 12250 8916 12256 8968
rect 12308 8956 12314 8968
rect 13173 8959 13231 8965
rect 13173 8956 13185 8959
rect 12308 8928 13185 8956
rect 12308 8916 12314 8928
rect 13173 8925 13185 8928
rect 13219 8925 13231 8959
rect 13173 8919 13231 8925
rect 14826 8916 14832 8968
rect 14884 8956 14890 8968
rect 15574 8959 15632 8965
rect 15574 8956 15586 8959
rect 14884 8928 15586 8956
rect 14884 8916 14890 8928
rect 15574 8925 15586 8928
rect 15620 8925 15632 8959
rect 15574 8919 15632 8925
rect 15841 8959 15899 8965
rect 15841 8925 15853 8959
rect 15887 8956 15899 8959
rect 16206 8956 16212 8968
rect 15887 8928 16212 8956
rect 15887 8925 15899 8928
rect 15841 8919 15899 8925
rect 16206 8916 16212 8928
rect 16264 8916 16270 8968
rect 19886 8916 19892 8968
rect 19944 8916 19950 8968
rect 20073 8959 20131 8965
rect 20073 8925 20085 8959
rect 20119 8956 20131 8959
rect 21450 8956 21456 8968
rect 20119 8928 21456 8956
rect 20119 8925 20131 8928
rect 20073 8919 20131 8925
rect 21450 8916 21456 8928
rect 21508 8916 21514 8968
rect 22925 8959 22983 8965
rect 22925 8925 22937 8959
rect 22971 8956 22983 8959
rect 23842 8956 23848 8968
rect 22971 8928 23848 8956
rect 22971 8925 22983 8928
rect 22925 8919 22983 8925
rect 23842 8916 23848 8928
rect 23900 8916 23906 8968
rect 24581 8959 24639 8965
rect 24581 8925 24593 8959
rect 24627 8956 24639 8959
rect 24670 8956 24676 8968
rect 24627 8928 24676 8956
rect 24627 8925 24639 8928
rect 24581 8919 24639 8925
rect 9490 8888 9496 8900
rect 7944 8860 9496 8888
rect 9490 8848 9496 8860
rect 9548 8848 9554 8900
rect 12986 8848 12992 8900
rect 13044 8848 13050 8900
rect 22278 8848 22284 8900
rect 22336 8888 22342 8900
rect 24596 8888 24624 8919
rect 24670 8916 24676 8928
rect 24728 8916 24734 8968
rect 24762 8916 24768 8968
rect 24820 8916 24826 8968
rect 27522 8916 27528 8968
rect 27580 8956 27586 8968
rect 28077 8959 28135 8965
rect 28077 8956 28089 8959
rect 27580 8928 28089 8956
rect 27580 8916 27586 8928
rect 28077 8925 28089 8928
rect 28123 8925 28135 8959
rect 28077 8919 28135 8925
rect 28261 8959 28319 8965
rect 28261 8925 28273 8959
rect 28307 8956 28319 8959
rect 28902 8956 28908 8968
rect 28307 8928 28908 8956
rect 28307 8925 28319 8928
rect 28261 8919 28319 8925
rect 28902 8916 28908 8928
rect 28960 8916 28966 8968
rect 29089 8959 29147 8965
rect 29089 8925 29101 8959
rect 29135 8956 29147 8959
rect 30101 8959 30159 8965
rect 30101 8956 30113 8959
rect 29135 8928 30113 8956
rect 29135 8925 29147 8928
rect 29089 8919 29147 8925
rect 30101 8925 30113 8928
rect 30147 8956 30159 8959
rect 30190 8956 30196 8968
rect 30147 8928 30196 8956
rect 30147 8925 30159 8928
rect 30101 8919 30159 8925
rect 30190 8916 30196 8928
rect 30248 8916 30254 8968
rect 22336 8860 24624 8888
rect 22336 8848 22342 8860
rect 27706 8848 27712 8900
rect 27764 8848 27770 8900
rect 27798 8848 27804 8900
rect 27856 8888 27862 8900
rect 28721 8891 28779 8897
rect 28721 8888 28733 8891
rect 27856 8860 28733 8888
rect 27856 8848 27862 8860
rect 28721 8857 28733 8860
rect 28767 8857 28779 8891
rect 28721 8851 28779 8857
rect 8573 8823 8631 8829
rect 8573 8789 8585 8823
rect 8619 8820 8631 8823
rect 8754 8820 8760 8832
rect 8619 8792 8760 8820
rect 8619 8789 8631 8792
rect 8573 8783 8631 8789
rect 8754 8780 8760 8792
rect 8812 8780 8818 8832
rect 13078 8780 13084 8832
rect 13136 8820 13142 8832
rect 13357 8823 13415 8829
rect 13357 8820 13369 8823
rect 13136 8792 13369 8820
rect 13136 8780 13142 8792
rect 13357 8789 13369 8792
rect 13403 8789 13415 8823
rect 13357 8783 13415 8789
rect 19978 8780 19984 8832
rect 20036 8780 20042 8832
rect 27890 8780 27896 8832
rect 27948 8780 27954 8832
rect 27982 8780 27988 8832
rect 28040 8780 28046 8832
rect 1104 8730 30976 8752
rect 1104 8678 8378 8730
rect 8430 8678 8442 8730
rect 8494 8678 8506 8730
rect 8558 8678 8570 8730
rect 8622 8678 8634 8730
rect 8686 8678 15806 8730
rect 15858 8678 15870 8730
rect 15922 8678 15934 8730
rect 15986 8678 15998 8730
rect 16050 8678 16062 8730
rect 16114 8678 23234 8730
rect 23286 8678 23298 8730
rect 23350 8678 23362 8730
rect 23414 8678 23426 8730
rect 23478 8678 23490 8730
rect 23542 8678 30662 8730
rect 30714 8678 30726 8730
rect 30778 8678 30790 8730
rect 30842 8678 30854 8730
rect 30906 8678 30918 8730
rect 30970 8678 30976 8730
rect 1104 8656 30976 8678
rect 8294 8576 8300 8628
rect 8352 8576 8358 8628
rect 12894 8576 12900 8628
rect 12952 8576 12958 8628
rect 18601 8619 18659 8625
rect 18601 8585 18613 8619
rect 18647 8616 18659 8619
rect 19058 8616 19064 8628
rect 18647 8588 19064 8616
rect 18647 8585 18659 8588
rect 18601 8579 18659 8585
rect 19058 8576 19064 8588
rect 19116 8576 19122 8628
rect 19426 8616 19432 8628
rect 19168 8588 19432 8616
rect 9214 8508 9220 8560
rect 9272 8548 9278 8560
rect 9585 8551 9643 8557
rect 9585 8548 9597 8551
rect 9272 8520 9597 8548
rect 9272 8508 9278 8520
rect 9585 8517 9597 8520
rect 9631 8517 9643 8551
rect 9585 8511 9643 8517
rect 12345 8551 12403 8557
rect 12345 8517 12357 8551
rect 12391 8548 12403 8551
rect 13173 8551 13231 8557
rect 13173 8548 13185 8551
rect 12391 8520 13185 8548
rect 12391 8517 12403 8520
rect 12345 8511 12403 8517
rect 13173 8517 13185 8520
rect 13219 8517 13231 8551
rect 13173 8511 13231 8517
rect 13265 8551 13323 8557
rect 13265 8517 13277 8551
rect 13311 8548 13323 8551
rect 14001 8551 14059 8557
rect 14001 8548 14013 8551
rect 13311 8520 14013 8548
rect 13311 8517 13323 8520
rect 13265 8511 13323 8517
rect 14001 8517 14013 8520
rect 14047 8517 14059 8551
rect 19168 8548 19196 8588
rect 19426 8576 19432 8588
rect 19484 8576 19490 8628
rect 25225 8619 25283 8625
rect 25225 8585 25237 8619
rect 25271 8616 25283 8619
rect 27430 8616 27436 8628
rect 25271 8588 27436 8616
rect 25271 8585 25283 8588
rect 25225 8579 25283 8585
rect 27430 8576 27436 8588
rect 27488 8576 27494 8628
rect 28629 8619 28687 8625
rect 28629 8585 28641 8619
rect 28675 8616 28687 8619
rect 29362 8616 29368 8628
rect 28675 8588 29368 8616
rect 28675 8585 28687 8588
rect 28629 8579 28687 8585
rect 29362 8576 29368 8588
rect 29420 8576 29426 8628
rect 18354 8520 19196 8548
rect 14001 8511 14059 8517
rect 19978 8508 19984 8560
rect 20036 8508 20042 8560
rect 24762 8548 24768 8560
rect 22020 8520 24768 8548
rect 5350 8440 5356 8492
rect 5408 8480 5414 8492
rect 5813 8483 5871 8489
rect 5813 8480 5825 8483
rect 5408 8452 5825 8480
rect 5408 8440 5414 8452
rect 5813 8449 5825 8452
rect 5859 8480 5871 8483
rect 6549 8483 6607 8489
rect 6549 8480 6561 8483
rect 5859 8452 6561 8480
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 6549 8449 6561 8452
rect 6595 8480 6607 8483
rect 9306 8480 9312 8492
rect 6595 8452 9312 8480
rect 6595 8449 6607 8452
rect 6549 8443 6607 8449
rect 9306 8440 9312 8452
rect 9364 8440 9370 8492
rect 11146 8440 11152 8492
rect 11204 8440 11210 8492
rect 11238 8440 11244 8492
rect 11296 8480 11302 8492
rect 12250 8480 12256 8492
rect 11296 8452 12256 8480
rect 11296 8440 11302 8452
rect 12250 8440 12256 8452
rect 12308 8440 12314 8492
rect 12437 8483 12495 8489
rect 12437 8449 12449 8483
rect 12483 8480 12495 8483
rect 12986 8480 12992 8492
rect 12483 8452 12992 8480
rect 12483 8449 12495 8452
rect 12437 8443 12495 8449
rect 12986 8440 12992 8452
rect 13044 8440 13050 8492
rect 13078 8440 13084 8492
rect 13136 8440 13142 8492
rect 13446 8440 13452 8492
rect 13504 8440 13510 8492
rect 13906 8440 13912 8492
rect 13964 8440 13970 8492
rect 14093 8483 14151 8489
rect 14093 8449 14105 8483
rect 14139 8480 14151 8483
rect 14458 8480 14464 8492
rect 14139 8452 14464 8480
rect 14139 8449 14151 8452
rect 14093 8443 14151 8449
rect 14458 8440 14464 8452
rect 14516 8440 14522 8492
rect 19061 8483 19119 8489
rect 19061 8480 19073 8483
rect 18984 8452 19073 8480
rect 18984 8424 19012 8452
rect 19061 8449 19073 8452
rect 19107 8449 19119 8483
rect 19061 8443 19119 8449
rect 19150 8440 19156 8492
rect 19208 8480 19214 8492
rect 19429 8483 19487 8489
rect 19429 8480 19441 8483
rect 19208 8452 19441 8480
rect 19208 8440 19214 8452
rect 19429 8449 19441 8452
rect 19475 8449 19487 8483
rect 19429 8443 19487 8449
rect 21450 8440 21456 8492
rect 21508 8480 21514 8492
rect 22020 8489 22048 8520
rect 24762 8508 24768 8520
rect 24820 8508 24826 8560
rect 27522 8508 27528 8560
rect 27580 8548 27586 8560
rect 27801 8551 27859 8557
rect 27801 8548 27813 8551
rect 27580 8520 27813 8548
rect 27580 8508 27586 8520
rect 27801 8517 27813 8520
rect 27847 8517 27859 8551
rect 27801 8511 27859 8517
rect 22005 8483 22063 8489
rect 22005 8480 22017 8483
rect 21508 8452 22017 8480
rect 21508 8440 21514 8452
rect 22005 8449 22017 8452
rect 22051 8449 22063 8483
rect 22005 8443 22063 8449
rect 22189 8483 22247 8489
rect 22189 8449 22201 8483
rect 22235 8480 22247 8483
rect 22278 8480 22284 8492
rect 22235 8452 22284 8480
rect 22235 8449 22247 8452
rect 22189 8443 22247 8449
rect 22278 8440 22284 8452
rect 22336 8440 22342 8492
rect 23842 8440 23848 8492
rect 23900 8440 23906 8492
rect 24101 8483 24159 8489
rect 24101 8480 24113 8483
rect 23952 8452 24113 8480
rect 5442 8372 5448 8424
rect 5500 8412 5506 8424
rect 8294 8412 8300 8424
rect 5500 8384 8300 8412
rect 5500 8372 5506 8384
rect 8294 8372 8300 8384
rect 8352 8372 8358 8424
rect 16853 8415 16911 8421
rect 16853 8381 16865 8415
rect 16899 8381 16911 8415
rect 16853 8375 16911 8381
rect 6641 8347 6699 8353
rect 6641 8313 6653 8347
rect 6687 8344 6699 8347
rect 6914 8344 6920 8356
rect 6687 8316 6920 8344
rect 6687 8313 6699 8316
rect 6641 8307 6699 8313
rect 6914 8304 6920 8316
rect 6972 8304 6978 8356
rect 5718 8236 5724 8288
rect 5776 8236 5782 8288
rect 11054 8236 11060 8288
rect 11112 8236 11118 8288
rect 16666 8236 16672 8288
rect 16724 8276 16730 8288
rect 16868 8276 16896 8375
rect 17126 8372 17132 8424
rect 17184 8412 17190 8424
rect 17184 8384 18552 8412
rect 17184 8372 17190 8384
rect 18524 8344 18552 8384
rect 18966 8372 18972 8424
rect 19024 8372 19030 8424
rect 23952 8412 23980 8452
rect 24101 8449 24113 8452
rect 24147 8449 24159 8483
rect 24101 8443 24159 8449
rect 27617 8483 27675 8489
rect 27617 8449 27629 8483
rect 27663 8480 27675 8483
rect 27706 8480 27712 8492
rect 27663 8452 27712 8480
rect 27663 8449 27675 8452
rect 27617 8443 27675 8449
rect 27706 8440 27712 8452
rect 27764 8440 27770 8492
rect 27890 8440 27896 8492
rect 27948 8440 27954 8492
rect 27982 8440 27988 8492
rect 28040 8489 28046 8492
rect 28040 8483 28079 8489
rect 28067 8480 28079 8483
rect 28534 8480 28540 8492
rect 28067 8452 28540 8480
rect 28067 8449 28079 8452
rect 28040 8443 28079 8449
rect 28040 8440 28046 8443
rect 28534 8440 28540 8452
rect 28592 8440 28598 8492
rect 19076 8384 23980 8412
rect 19076 8344 19104 8384
rect 27798 8372 27804 8424
rect 27856 8372 27862 8424
rect 18524 8316 19104 8344
rect 18598 8276 18604 8288
rect 16724 8248 18604 8276
rect 16724 8236 16730 8248
rect 18598 8236 18604 8248
rect 18656 8236 18662 8288
rect 20806 8236 20812 8288
rect 20864 8285 20870 8288
rect 20864 8279 20913 8285
rect 20864 8245 20867 8279
rect 20901 8245 20913 8279
rect 20864 8239 20913 8245
rect 20864 8236 20870 8239
rect 22094 8236 22100 8288
rect 22152 8236 22158 8288
rect 1104 8186 30820 8208
rect 1104 8134 4664 8186
rect 4716 8134 4728 8186
rect 4780 8134 4792 8186
rect 4844 8134 4856 8186
rect 4908 8134 4920 8186
rect 4972 8134 12092 8186
rect 12144 8134 12156 8186
rect 12208 8134 12220 8186
rect 12272 8134 12284 8186
rect 12336 8134 12348 8186
rect 12400 8134 19520 8186
rect 19572 8134 19584 8186
rect 19636 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 26948 8186
rect 27000 8134 27012 8186
rect 27064 8134 27076 8186
rect 27128 8134 27140 8186
rect 27192 8134 27204 8186
rect 27256 8134 30820 8186
rect 1104 8112 30820 8134
rect 12526 8032 12532 8084
rect 12584 8032 12590 8084
rect 13081 8075 13139 8081
rect 13081 8041 13093 8075
rect 13127 8072 13139 8075
rect 13446 8072 13452 8084
rect 13127 8044 13452 8072
rect 13127 8041 13139 8044
rect 13081 8035 13139 8041
rect 13446 8032 13452 8044
rect 13504 8032 13510 8084
rect 16209 8075 16267 8081
rect 16209 8041 16221 8075
rect 16255 8072 16267 8075
rect 16666 8072 16672 8084
rect 16255 8044 16672 8072
rect 16255 8041 16267 8044
rect 16209 8035 16267 8041
rect 16666 8032 16672 8044
rect 16724 8032 16730 8084
rect 16807 8075 16865 8081
rect 16807 8041 16819 8075
rect 16853 8072 16865 8075
rect 17126 8072 17132 8084
rect 16853 8044 17132 8072
rect 16853 8041 16865 8044
rect 16807 8035 16865 8041
rect 17126 8032 17132 8044
rect 17184 8032 17190 8084
rect 19426 8032 19432 8084
rect 19484 8072 19490 8084
rect 19521 8075 19579 8081
rect 19521 8072 19533 8075
rect 19484 8044 19533 8072
rect 19484 8032 19490 8044
rect 19521 8041 19533 8044
rect 19567 8041 19579 8075
rect 19521 8035 19579 8041
rect 25961 8075 26019 8081
rect 25961 8041 25973 8075
rect 26007 8072 26019 8075
rect 27522 8072 27528 8084
rect 26007 8044 27528 8072
rect 26007 8041 26019 8044
rect 25961 8035 26019 8041
rect 27522 8032 27528 8044
rect 27580 8032 27586 8084
rect 5353 7939 5411 7945
rect 5353 7905 5365 7939
rect 5399 7936 5411 7939
rect 5718 7936 5724 7948
rect 5399 7908 5724 7936
rect 5399 7905 5411 7908
rect 5353 7899 5411 7905
rect 5718 7896 5724 7908
rect 5776 7896 5782 7948
rect 11054 7896 11060 7948
rect 11112 7896 11118 7948
rect 18598 7896 18604 7948
rect 18656 7936 18662 7948
rect 18966 7936 18972 7948
rect 18656 7908 18972 7936
rect 18656 7896 18662 7908
rect 18966 7896 18972 7908
rect 19024 7936 19030 7948
rect 19024 7908 20484 7936
rect 19024 7896 19030 7908
rect 20456 7880 20484 7908
rect 20806 7896 20812 7948
rect 20864 7896 20870 7948
rect 7653 7871 7711 7877
rect 7653 7837 7665 7871
rect 7699 7868 7711 7871
rect 7834 7868 7840 7880
rect 7699 7840 7840 7868
rect 7699 7837 7711 7840
rect 7653 7831 7711 7837
rect 5629 7803 5687 7809
rect 5629 7769 5641 7803
rect 5675 7769 5687 7803
rect 5629 7763 5687 7769
rect 5644 7732 5672 7763
rect 6086 7760 6092 7812
rect 6144 7760 6150 7812
rect 6638 7732 6644 7744
rect 5644 7704 6644 7732
rect 6638 7692 6644 7704
rect 6696 7692 6702 7744
rect 7098 7692 7104 7744
rect 7156 7732 7162 7744
rect 7668 7732 7696 7831
rect 7834 7828 7840 7840
rect 7892 7828 7898 7880
rect 9306 7828 9312 7880
rect 9364 7828 9370 7880
rect 10778 7828 10784 7880
rect 10836 7828 10842 7880
rect 13449 7871 13507 7877
rect 13449 7837 13461 7871
rect 13495 7868 13507 7871
rect 14458 7868 14464 7880
rect 13495 7840 14464 7868
rect 13495 7837 13507 7840
rect 13449 7831 13507 7837
rect 14458 7828 14464 7840
rect 14516 7828 14522 7880
rect 15194 7828 15200 7880
rect 15252 7868 15258 7880
rect 15933 7871 15991 7877
rect 15933 7868 15945 7871
rect 15252 7840 15945 7868
rect 15252 7828 15258 7840
rect 15933 7837 15945 7840
rect 15979 7837 15991 7871
rect 15933 7831 15991 7837
rect 18233 7871 18291 7877
rect 18233 7837 18245 7871
rect 18279 7868 18291 7871
rect 18506 7868 18512 7880
rect 18279 7840 18512 7868
rect 18279 7837 18291 7840
rect 18233 7831 18291 7837
rect 18506 7828 18512 7840
rect 18564 7828 18570 7880
rect 19429 7871 19487 7877
rect 19429 7837 19441 7871
rect 19475 7837 19487 7871
rect 19429 7831 19487 7837
rect 11698 7760 11704 7812
rect 11756 7760 11762 7812
rect 13265 7803 13323 7809
rect 13265 7769 13277 7803
rect 13311 7800 13323 7803
rect 13906 7800 13912 7812
rect 13311 7772 13912 7800
rect 13311 7769 13323 7772
rect 13265 7763 13323 7769
rect 7156 7704 7696 7732
rect 7156 7692 7162 7704
rect 7742 7692 7748 7744
rect 7800 7692 7806 7744
rect 8018 7692 8024 7744
rect 8076 7732 8082 7744
rect 9217 7735 9275 7741
rect 9217 7732 9229 7735
rect 8076 7704 9229 7732
rect 8076 7692 8082 7704
rect 9217 7701 9229 7704
rect 9263 7701 9275 7735
rect 9217 7695 9275 7701
rect 11054 7692 11060 7744
rect 11112 7732 11118 7744
rect 13280 7732 13308 7763
rect 13906 7760 13912 7772
rect 13964 7760 13970 7812
rect 17402 7760 17408 7812
rect 17460 7760 17466 7812
rect 11112 7704 13308 7732
rect 11112 7692 11118 7704
rect 17678 7692 17684 7744
rect 17736 7732 17742 7744
rect 19444 7732 19472 7831
rect 19610 7828 19616 7880
rect 19668 7868 19674 7880
rect 19886 7868 19892 7880
rect 19668 7840 19892 7868
rect 19668 7828 19674 7840
rect 19886 7828 19892 7840
rect 19944 7828 19950 7880
rect 20438 7828 20444 7880
rect 20496 7868 20502 7880
rect 20533 7871 20591 7877
rect 20533 7868 20545 7871
rect 20496 7840 20545 7868
rect 20496 7828 20502 7840
rect 20533 7837 20545 7840
rect 20579 7837 20591 7871
rect 20533 7831 20591 7837
rect 23842 7828 23848 7880
rect 23900 7868 23906 7880
rect 24302 7868 24308 7880
rect 23900 7840 24308 7868
rect 23900 7828 23906 7840
rect 24302 7828 24308 7840
rect 24360 7868 24366 7880
rect 24581 7871 24639 7877
rect 24581 7868 24593 7871
rect 24360 7840 24593 7868
rect 24360 7828 24366 7840
rect 24581 7837 24593 7840
rect 24627 7837 24639 7871
rect 24581 7831 24639 7837
rect 28534 7828 28540 7880
rect 28592 7828 28598 7880
rect 22094 7800 22100 7812
rect 22034 7772 22100 7800
rect 22094 7760 22100 7772
rect 22152 7760 22158 7812
rect 24826 7803 24884 7809
rect 24826 7800 24838 7803
rect 22296 7772 24838 7800
rect 17736 7704 19472 7732
rect 17736 7692 17742 7704
rect 22186 7692 22192 7744
rect 22244 7732 22250 7744
rect 22296 7741 22324 7772
rect 24826 7769 24838 7772
rect 24872 7769 24884 7803
rect 24826 7763 24884 7769
rect 22281 7735 22339 7741
rect 22281 7732 22293 7735
rect 22244 7704 22293 7732
rect 22244 7692 22250 7704
rect 22281 7701 22293 7704
rect 22327 7701 22339 7735
rect 22281 7695 22339 7701
rect 28442 7692 28448 7744
rect 28500 7692 28506 7744
rect 1104 7642 30976 7664
rect 1104 7590 8378 7642
rect 8430 7590 8442 7642
rect 8494 7590 8506 7642
rect 8558 7590 8570 7642
rect 8622 7590 8634 7642
rect 8686 7590 15806 7642
rect 15858 7590 15870 7642
rect 15922 7590 15934 7642
rect 15986 7590 15998 7642
rect 16050 7590 16062 7642
rect 16114 7590 23234 7642
rect 23286 7590 23298 7642
rect 23350 7590 23362 7642
rect 23414 7590 23426 7642
rect 23478 7590 23490 7642
rect 23542 7590 30662 7642
rect 30714 7590 30726 7642
rect 30778 7590 30790 7642
rect 30842 7590 30854 7642
rect 30906 7590 30918 7642
rect 30970 7590 30976 7642
rect 1104 7568 30976 7590
rect 5997 7531 6055 7537
rect 5997 7497 6009 7531
rect 6043 7528 6055 7531
rect 6086 7528 6092 7540
rect 6043 7500 6092 7528
rect 6043 7497 6055 7500
rect 5997 7491 6055 7497
rect 6086 7488 6092 7500
rect 6144 7488 6150 7540
rect 6638 7488 6644 7540
rect 6696 7488 6702 7540
rect 10778 7488 10784 7540
rect 10836 7488 10842 7540
rect 11698 7488 11704 7540
rect 11756 7488 11762 7540
rect 13354 7528 13360 7540
rect 12636 7500 13360 7528
rect 5626 7460 5632 7472
rect 5368 7432 5632 7460
rect 5258 7352 5264 7404
rect 5316 7392 5322 7404
rect 5368 7401 5396 7432
rect 5626 7420 5632 7432
rect 5684 7420 5690 7472
rect 8018 7420 8024 7472
rect 8076 7420 8082 7472
rect 8754 7420 8760 7472
rect 8812 7420 8818 7472
rect 5353 7395 5411 7401
rect 5353 7392 5365 7395
rect 5316 7364 5365 7392
rect 5316 7352 5322 7364
rect 5353 7361 5365 7364
rect 5399 7361 5411 7395
rect 5353 7355 5411 7361
rect 5442 7352 5448 7404
rect 5500 7352 5506 7404
rect 6733 7395 6791 7401
rect 6733 7361 6745 7395
rect 6779 7392 6791 7395
rect 7098 7392 7104 7404
rect 6779 7364 7104 7392
rect 6779 7361 6791 7364
rect 6733 7355 6791 7361
rect 7098 7352 7104 7364
rect 7156 7352 7162 7404
rect 7742 7352 7748 7404
rect 7800 7352 7806 7404
rect 10689 7395 10747 7401
rect 10689 7361 10701 7395
rect 10735 7392 10747 7395
rect 11238 7392 11244 7404
rect 10735 7364 11244 7392
rect 10735 7361 10747 7364
rect 10689 7355 10747 7361
rect 9306 7284 9312 7336
rect 9364 7324 9370 7336
rect 9493 7327 9551 7333
rect 9493 7324 9505 7327
rect 9364 7296 9505 7324
rect 9364 7284 9370 7296
rect 9493 7293 9505 7296
rect 9539 7324 9551 7327
rect 10704 7324 10732 7355
rect 11238 7352 11244 7364
rect 11296 7352 11302 7404
rect 12529 7395 12587 7401
rect 12529 7361 12541 7395
rect 12575 7392 12587 7395
rect 12636 7392 12664 7500
rect 13354 7488 13360 7500
rect 13412 7528 13418 7540
rect 16390 7528 16396 7540
rect 13412 7500 16396 7528
rect 13412 7488 13418 7500
rect 16390 7488 16396 7500
rect 16448 7488 16454 7540
rect 18506 7488 18512 7540
rect 18564 7528 18570 7540
rect 18601 7531 18659 7537
rect 18601 7528 18613 7531
rect 18564 7500 18613 7528
rect 18564 7488 18570 7500
rect 18601 7497 18613 7500
rect 18647 7497 18659 7531
rect 18601 7491 18659 7497
rect 28534 7488 28540 7540
rect 28592 7528 28598 7540
rect 29457 7531 29515 7537
rect 29457 7528 29469 7531
rect 28592 7500 29469 7528
rect 28592 7488 28598 7500
rect 29457 7497 29469 7500
rect 29503 7497 29515 7531
rect 29457 7491 29515 7497
rect 16209 7463 16267 7469
rect 16209 7429 16221 7463
rect 16255 7460 16267 7463
rect 22278 7460 22284 7472
rect 16255 7432 17618 7460
rect 21284 7432 22284 7460
rect 16255 7429 16267 7432
rect 16209 7423 16267 7429
rect 12575 7364 12664 7392
rect 16117 7395 16175 7401
rect 12575 7361 12587 7364
rect 12529 7355 12587 7361
rect 16117 7361 16129 7395
rect 16163 7361 16175 7395
rect 16117 7355 16175 7361
rect 16301 7395 16359 7401
rect 16301 7361 16313 7395
rect 16347 7392 16359 7395
rect 16666 7392 16672 7404
rect 16347 7364 16672 7392
rect 16347 7361 16359 7364
rect 16301 7355 16359 7361
rect 9539 7296 10732 7324
rect 9539 7293 9551 7296
rect 9493 7287 9551 7293
rect 12434 7284 12440 7336
rect 12492 7284 12498 7336
rect 16132 7324 16160 7355
rect 16666 7352 16672 7364
rect 16724 7352 16730 7404
rect 16758 7352 16764 7404
rect 16816 7392 16822 7404
rect 21284 7401 21312 7432
rect 16853 7395 16911 7401
rect 16853 7392 16865 7395
rect 16816 7364 16865 7392
rect 16816 7352 16822 7364
rect 16853 7361 16865 7364
rect 16899 7361 16911 7395
rect 21269 7395 21327 7401
rect 21269 7392 21281 7395
rect 16853 7355 16911 7361
rect 19628 7364 21281 7392
rect 19628 7336 19656 7364
rect 21269 7361 21281 7364
rect 21315 7361 21327 7395
rect 21269 7355 21327 7361
rect 21450 7352 21456 7404
rect 21508 7352 21514 7404
rect 21928 7390 21956 7432
rect 22278 7420 22284 7432
rect 22336 7460 22342 7472
rect 28344 7463 28402 7469
rect 22336 7432 22876 7460
rect 22336 7420 22342 7432
rect 22848 7401 22876 7432
rect 28344 7429 28356 7463
rect 28390 7460 28402 7463
rect 28442 7460 28448 7472
rect 28390 7432 28448 7460
rect 28390 7429 28402 7432
rect 28344 7423 28402 7429
rect 28442 7420 28448 7432
rect 28500 7420 28506 7472
rect 22005 7395 22063 7401
rect 22005 7390 22017 7395
rect 21928 7362 22017 7390
rect 22005 7361 22017 7362
rect 22051 7361 22063 7395
rect 22005 7355 22063 7361
rect 22189 7395 22247 7401
rect 22189 7361 22201 7395
rect 22235 7392 22247 7395
rect 22649 7395 22707 7401
rect 22649 7392 22661 7395
rect 22235 7364 22661 7392
rect 22235 7361 22247 7364
rect 22189 7355 22247 7361
rect 22649 7361 22661 7364
rect 22695 7361 22707 7395
rect 22649 7355 22707 7361
rect 22833 7395 22891 7401
rect 22833 7361 22845 7395
rect 22879 7361 22891 7395
rect 22833 7355 22891 7361
rect 25409 7395 25467 7401
rect 25409 7361 25421 7395
rect 25455 7392 25467 7395
rect 25958 7392 25964 7404
rect 25455 7364 25964 7392
rect 25455 7361 25467 7364
rect 25409 7355 25467 7361
rect 16206 7324 16212 7336
rect 16132 7296 16212 7324
rect 16206 7284 16212 7296
rect 16264 7324 16270 7336
rect 16264 7296 16574 7324
rect 16264 7284 16270 7296
rect 16546 7188 16574 7296
rect 17126 7284 17132 7336
rect 17184 7284 17190 7336
rect 17494 7284 17500 7336
rect 17552 7324 17558 7336
rect 19610 7324 19616 7336
rect 17552 7296 19616 7324
rect 17552 7284 17558 7296
rect 19610 7284 19616 7296
rect 19668 7284 19674 7336
rect 21468 7256 21496 7352
rect 22204 7256 22232 7355
rect 25958 7352 25964 7364
rect 26016 7352 26022 7404
rect 27614 7352 27620 7404
rect 27672 7352 27678 7404
rect 27525 7327 27583 7333
rect 27525 7293 27537 7327
rect 27571 7324 27583 7327
rect 28077 7327 28135 7333
rect 28077 7324 28089 7327
rect 27571 7296 28089 7324
rect 27571 7293 27583 7296
rect 27525 7287 27583 7293
rect 28077 7293 28089 7296
rect 28123 7293 28135 7327
rect 28077 7287 28135 7293
rect 21468 7228 22232 7256
rect 17678 7188 17684 7200
rect 16546 7160 17684 7188
rect 17678 7148 17684 7160
rect 17736 7148 17742 7200
rect 21358 7148 21364 7200
rect 21416 7148 21422 7200
rect 22097 7191 22155 7197
rect 22097 7157 22109 7191
rect 22143 7188 22155 7191
rect 22646 7188 22652 7200
rect 22143 7160 22652 7188
rect 22143 7157 22155 7160
rect 22097 7151 22155 7157
rect 22646 7148 22652 7160
rect 22704 7148 22710 7200
rect 22741 7191 22799 7197
rect 22741 7157 22753 7191
rect 22787 7188 22799 7191
rect 22830 7188 22836 7200
rect 22787 7160 22836 7188
rect 22787 7157 22799 7160
rect 22741 7151 22799 7157
rect 22830 7148 22836 7160
rect 22888 7148 22894 7200
rect 25314 7148 25320 7200
rect 25372 7148 25378 7200
rect 1104 7098 30820 7120
rect 1104 7046 4664 7098
rect 4716 7046 4728 7098
rect 4780 7046 4792 7098
rect 4844 7046 4856 7098
rect 4908 7046 4920 7098
rect 4972 7046 12092 7098
rect 12144 7046 12156 7098
rect 12208 7046 12220 7098
rect 12272 7046 12284 7098
rect 12336 7046 12348 7098
rect 12400 7046 19520 7098
rect 19572 7046 19584 7098
rect 19636 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 26948 7098
rect 27000 7046 27012 7098
rect 27064 7046 27076 7098
rect 27128 7046 27140 7098
rect 27192 7046 27204 7098
rect 27256 7046 30820 7098
rect 1104 7024 30820 7046
rect 6914 6944 6920 6996
rect 6972 6993 6978 6996
rect 6972 6987 6987 6993
rect 6975 6953 6987 6987
rect 6972 6947 6987 6953
rect 6972 6944 6978 6947
rect 25958 6944 25964 6996
rect 26016 6944 26022 6996
rect 5350 6808 5356 6860
rect 5408 6848 5414 6860
rect 5445 6851 5503 6857
rect 5445 6848 5457 6851
rect 5408 6820 5457 6848
rect 5408 6808 5414 6820
rect 5445 6817 5457 6820
rect 5491 6817 5503 6851
rect 5445 6811 5503 6817
rect 8481 6851 8539 6857
rect 8481 6817 8493 6851
rect 8527 6848 8539 6851
rect 9125 6851 9183 6857
rect 9125 6848 9137 6851
rect 8527 6820 9137 6848
rect 8527 6817 8539 6820
rect 8481 6811 8539 6817
rect 9125 6817 9137 6820
rect 9171 6817 9183 6851
rect 9125 6811 9183 6817
rect 9950 6808 9956 6860
rect 10008 6848 10014 6860
rect 16071 6851 16129 6857
rect 10008 6820 15424 6848
rect 10008 6808 10014 6820
rect 7190 6740 7196 6792
rect 7248 6740 7254 6792
rect 8573 6783 8631 6789
rect 8573 6749 8585 6783
rect 8619 6780 8631 6783
rect 8754 6780 8760 6792
rect 8619 6752 8760 6780
rect 8619 6749 8631 6752
rect 8573 6743 8631 6749
rect 8754 6740 8760 6752
rect 8812 6740 8818 6792
rect 14277 6783 14335 6789
rect 14277 6749 14289 6783
rect 14323 6749 14335 6783
rect 14277 6743 14335 6749
rect 5902 6672 5908 6724
rect 5960 6672 5966 6724
rect 9398 6672 9404 6724
rect 9456 6672 9462 6724
rect 10042 6672 10048 6724
rect 10100 6672 10106 6724
rect 8294 6604 8300 6656
rect 8352 6644 8358 6656
rect 10873 6647 10931 6653
rect 10873 6644 10885 6647
rect 8352 6616 10885 6644
rect 8352 6604 8358 6616
rect 10873 6613 10885 6616
rect 10919 6644 10931 6647
rect 11054 6644 11060 6656
rect 10919 6616 11060 6644
rect 10919 6613 10931 6616
rect 10873 6607 10931 6613
rect 11054 6604 11060 6616
rect 11112 6604 11118 6656
rect 13538 6604 13544 6656
rect 13596 6644 13602 6656
rect 14292 6644 14320 6743
rect 14642 6740 14648 6792
rect 14700 6740 14706 6792
rect 15396 6780 15424 6820
rect 16071 6817 16083 6851
rect 16117 6848 16129 6851
rect 17126 6848 17132 6860
rect 16117 6820 17132 6848
rect 16117 6817 16129 6820
rect 16071 6811 16129 6817
rect 17126 6808 17132 6820
rect 17184 6808 17190 6860
rect 17402 6808 17408 6860
rect 17460 6848 17466 6860
rect 17589 6851 17647 6857
rect 17589 6848 17601 6851
rect 17460 6820 17601 6848
rect 17460 6808 17466 6820
rect 17589 6817 17601 6820
rect 17635 6817 17647 6851
rect 17589 6811 17647 6817
rect 20438 6808 20444 6860
rect 20496 6808 20502 6860
rect 20809 6851 20867 6857
rect 20809 6817 20821 6851
rect 20855 6848 20867 6851
rect 22186 6848 22192 6860
rect 20855 6820 22192 6848
rect 20855 6817 20867 6820
rect 20809 6811 20867 6817
rect 22186 6808 22192 6820
rect 22244 6808 22250 6860
rect 26881 6851 26939 6857
rect 26881 6817 26893 6851
rect 26927 6848 26939 6851
rect 27706 6848 27712 6860
rect 26927 6820 27712 6848
rect 26927 6817 26939 6820
rect 26881 6811 26939 6817
rect 27706 6808 27712 6820
rect 27764 6808 27770 6860
rect 29089 6851 29147 6857
rect 29089 6817 29101 6851
rect 29135 6848 29147 6851
rect 30006 6848 30012 6860
rect 29135 6820 30012 6848
rect 29135 6817 29147 6820
rect 29089 6811 29147 6817
rect 30006 6808 30012 6820
rect 30064 6808 30070 6860
rect 16577 6783 16635 6789
rect 16577 6780 16589 6783
rect 15396 6752 16589 6780
rect 16577 6749 16589 6752
rect 16623 6749 16635 6783
rect 16577 6743 16635 6749
rect 16666 6740 16672 6792
rect 16724 6780 16730 6792
rect 16853 6783 16911 6789
rect 16853 6780 16865 6783
rect 16724 6752 16865 6780
rect 16724 6740 16730 6752
rect 16853 6749 16865 6752
rect 16899 6780 16911 6783
rect 17494 6780 17500 6792
rect 16899 6752 17500 6780
rect 16899 6749 16911 6752
rect 16853 6743 16911 6749
rect 17494 6740 17500 6752
rect 17552 6740 17558 6792
rect 17678 6740 17684 6792
rect 17736 6740 17742 6792
rect 24578 6740 24584 6792
rect 24636 6740 24642 6792
rect 24848 6783 24906 6789
rect 24848 6749 24860 6783
rect 24894 6780 24906 6783
rect 25314 6780 25320 6792
rect 24894 6752 25320 6780
rect 24894 6749 24906 6752
rect 24848 6743 24906 6749
rect 25314 6740 25320 6752
rect 25372 6740 25378 6792
rect 25958 6740 25964 6792
rect 26016 6780 26022 6792
rect 27157 6783 27215 6789
rect 27157 6780 27169 6783
rect 26016 6752 27169 6780
rect 26016 6740 26022 6752
rect 27157 6749 27169 6752
rect 27203 6749 27215 6783
rect 27157 6743 27215 6749
rect 27433 6783 27491 6789
rect 27433 6749 27445 6783
rect 27479 6780 27491 6783
rect 28810 6780 28816 6792
rect 27479 6752 28816 6780
rect 27479 6749 27491 6752
rect 27433 6743 27491 6749
rect 28810 6740 28816 6752
rect 28868 6740 28874 6792
rect 28902 6740 28908 6792
rect 28960 6740 28966 6792
rect 16482 6712 16488 6724
rect 15686 6684 16488 6712
rect 16482 6672 16488 6684
rect 16540 6672 16546 6724
rect 21358 6672 21364 6724
rect 21416 6672 21422 6724
rect 27065 6715 27123 6721
rect 27065 6681 27077 6715
rect 27111 6712 27123 6715
rect 27890 6712 27896 6724
rect 27111 6684 27896 6712
rect 27111 6681 27123 6684
rect 27065 6675 27123 6681
rect 27890 6672 27896 6684
rect 27948 6672 27954 6724
rect 14366 6644 14372 6656
rect 13596 6616 14372 6644
rect 13596 6604 13602 6616
rect 14366 6604 14372 6616
rect 14424 6644 14430 6656
rect 16850 6644 16856 6656
rect 14424 6616 16856 6644
rect 14424 6604 14430 6616
rect 16850 6604 16856 6616
rect 16908 6604 16914 6656
rect 22235 6647 22293 6653
rect 22235 6613 22247 6647
rect 22281 6644 22293 6647
rect 22370 6644 22376 6656
rect 22281 6616 22376 6644
rect 22281 6613 22293 6616
rect 22235 6607 22293 6613
rect 22370 6604 22376 6616
rect 22428 6604 22434 6656
rect 27249 6647 27307 6653
rect 27249 6613 27261 6647
rect 27295 6644 27307 6647
rect 27338 6644 27344 6656
rect 27295 6616 27344 6644
rect 27295 6613 27307 6616
rect 27249 6607 27307 6613
rect 27338 6604 27344 6616
rect 27396 6604 27402 6656
rect 28442 6604 28448 6656
rect 28500 6604 28506 6656
rect 1104 6554 30976 6576
rect 1104 6502 8378 6554
rect 8430 6502 8442 6554
rect 8494 6502 8506 6554
rect 8558 6502 8570 6554
rect 8622 6502 8634 6554
rect 8686 6502 15806 6554
rect 15858 6502 15870 6554
rect 15922 6502 15934 6554
rect 15986 6502 15998 6554
rect 16050 6502 16062 6554
rect 16114 6502 23234 6554
rect 23286 6502 23298 6554
rect 23350 6502 23362 6554
rect 23414 6502 23426 6554
rect 23478 6502 23490 6554
rect 23542 6502 30662 6554
rect 30714 6502 30726 6554
rect 30778 6502 30790 6554
rect 30842 6502 30854 6554
rect 30906 6502 30918 6554
rect 30970 6502 30976 6554
rect 1104 6480 30976 6502
rect 5902 6400 5908 6452
rect 5960 6440 5966 6452
rect 5997 6443 6055 6449
rect 5997 6440 6009 6443
rect 5960 6412 6009 6440
rect 5960 6400 5966 6412
rect 5997 6409 6009 6412
rect 6043 6409 6055 6443
rect 5997 6403 6055 6409
rect 6641 6443 6699 6449
rect 6641 6409 6653 6443
rect 6687 6440 6699 6443
rect 7190 6440 7196 6452
rect 6687 6412 7196 6440
rect 6687 6409 6699 6412
rect 6641 6403 6699 6409
rect 7190 6400 7196 6412
rect 7248 6400 7254 6452
rect 8389 6443 8447 6449
rect 8389 6409 8401 6443
rect 8435 6440 8447 6443
rect 9398 6440 9404 6452
rect 8435 6412 9404 6440
rect 8435 6409 8447 6412
rect 8389 6403 8447 6409
rect 9398 6400 9404 6412
rect 9456 6400 9462 6452
rect 9950 6440 9956 6452
rect 9508 6412 9956 6440
rect 5074 6332 5080 6384
rect 5132 6372 5138 6384
rect 9508 6372 9536 6412
rect 9950 6400 9956 6412
rect 10008 6400 10014 6452
rect 10042 6400 10048 6452
rect 10100 6400 10106 6452
rect 12618 6400 12624 6452
rect 12676 6440 12682 6452
rect 24578 6440 24584 6452
rect 12676 6412 24584 6440
rect 12676 6400 12682 6412
rect 24578 6400 24584 6412
rect 24636 6400 24642 6452
rect 27614 6400 27620 6452
rect 27672 6440 27678 6452
rect 28350 6440 28356 6452
rect 27672 6412 28356 6440
rect 27672 6400 27678 6412
rect 28350 6400 28356 6412
rect 28408 6440 28414 6452
rect 28537 6443 28595 6449
rect 28537 6440 28549 6443
rect 28408 6412 28549 6440
rect 28408 6400 28414 6412
rect 28537 6409 28549 6412
rect 28583 6409 28595 6443
rect 28537 6403 28595 6409
rect 5132 6344 9536 6372
rect 5132 6332 5138 6344
rect 11974 6332 11980 6384
rect 12032 6372 12038 6384
rect 12032 6344 12098 6372
rect 12032 6332 12038 6344
rect 22738 6332 22744 6384
rect 22796 6332 22802 6384
rect 28902 6332 28908 6384
rect 28960 6372 28966 6384
rect 28960 6344 30144 6372
rect 28960 6332 28966 6344
rect 5258 6264 5264 6316
rect 5316 6264 5322 6316
rect 5442 6264 5448 6316
rect 5500 6264 5506 6316
rect 6733 6307 6791 6313
rect 6733 6273 6745 6307
rect 6779 6304 6791 6307
rect 8294 6304 8300 6316
rect 6779 6276 8300 6304
rect 6779 6273 6791 6276
rect 6733 6267 6791 6273
rect 8294 6264 8300 6276
rect 8352 6264 8358 6316
rect 9398 6264 9404 6316
rect 9456 6264 9462 6316
rect 9493 6307 9551 6313
rect 9493 6273 9505 6307
rect 9539 6304 9551 6307
rect 9582 6304 9588 6316
rect 9539 6276 9588 6304
rect 9539 6273 9551 6276
rect 9493 6267 9551 6273
rect 9582 6264 9588 6276
rect 9640 6264 9646 6316
rect 10965 6307 11023 6313
rect 10965 6273 10977 6307
rect 11011 6273 11023 6307
rect 10965 6267 11023 6273
rect 8754 6196 8760 6248
rect 8812 6236 8818 6248
rect 10980 6236 11008 6267
rect 13538 6264 13544 6316
rect 13596 6264 13602 6316
rect 22370 6264 22376 6316
rect 22428 6264 22434 6316
rect 24302 6264 24308 6316
rect 24360 6264 24366 6316
rect 24561 6307 24619 6313
rect 24561 6304 24573 6307
rect 24412 6276 24573 6304
rect 8812 6208 11008 6236
rect 8812 6196 8818 6208
rect 10980 6168 11008 6208
rect 11057 6239 11115 6245
rect 11057 6205 11069 6239
rect 11103 6236 11115 6239
rect 13265 6239 13323 6245
rect 13265 6236 13277 6239
rect 11103 6208 13277 6236
rect 11103 6205 11115 6208
rect 11057 6199 11115 6205
rect 13265 6205 13277 6208
rect 13311 6205 13323 6239
rect 13265 6199 13323 6205
rect 21450 6196 21456 6248
rect 21508 6236 21514 6248
rect 22005 6239 22063 6245
rect 22005 6236 22017 6239
rect 21508 6208 22017 6236
rect 21508 6196 21514 6208
rect 22005 6205 22017 6208
rect 22051 6205 22063 6239
rect 24412 6236 24440 6276
rect 24561 6273 24573 6276
rect 24607 6273 24619 6307
rect 24561 6267 24619 6273
rect 25958 6264 25964 6316
rect 26016 6304 26022 6316
rect 26421 6307 26479 6313
rect 26421 6304 26433 6307
rect 26016 6276 26433 6304
rect 26016 6264 26022 6276
rect 26421 6273 26433 6276
rect 26467 6273 26479 6307
rect 26421 6267 26479 6273
rect 27424 6307 27482 6313
rect 27424 6273 27436 6307
rect 27470 6304 27482 6307
rect 29086 6304 29092 6316
rect 27470 6276 29092 6304
rect 27470 6273 27482 6276
rect 27424 6267 27482 6273
rect 29086 6264 29092 6276
rect 29144 6264 29150 6316
rect 30116 6313 30144 6344
rect 29273 6307 29331 6313
rect 29273 6273 29285 6307
rect 29319 6273 29331 6307
rect 29273 6267 29331 6273
rect 30101 6307 30159 6313
rect 30101 6273 30113 6307
rect 30147 6273 30159 6307
rect 30101 6267 30159 6273
rect 30285 6307 30343 6313
rect 30285 6273 30297 6307
rect 30331 6273 30343 6307
rect 30285 6267 30343 6273
rect 22005 6199 22063 6205
rect 24320 6208 24440 6236
rect 26513 6239 26571 6245
rect 11793 6171 11851 6177
rect 11793 6168 11805 6171
rect 10980 6140 11805 6168
rect 11793 6137 11805 6140
rect 11839 6137 11851 6171
rect 11793 6131 11851 6137
rect 21726 6060 21732 6112
rect 21784 6100 21790 6112
rect 23799 6103 23857 6109
rect 23799 6100 23811 6103
rect 21784 6072 23811 6100
rect 21784 6060 21790 6072
rect 23799 6069 23811 6072
rect 23845 6100 23857 6103
rect 24320 6100 24348 6208
rect 26513 6205 26525 6239
rect 26559 6236 26571 6239
rect 27157 6239 27215 6245
rect 27157 6236 27169 6239
rect 26559 6208 27169 6236
rect 26559 6205 26571 6208
rect 26513 6199 26571 6205
rect 27157 6205 27169 6208
rect 27203 6205 27215 6239
rect 27157 6199 27215 6205
rect 28810 6196 28816 6248
rect 28868 6236 28874 6248
rect 29288 6236 29316 6267
rect 28868 6208 29316 6236
rect 29365 6239 29423 6245
rect 28868 6196 28874 6208
rect 29365 6205 29377 6239
rect 29411 6236 29423 6239
rect 30193 6239 30251 6245
rect 30193 6236 30205 6239
rect 29411 6208 30205 6236
rect 29411 6205 29423 6208
rect 29365 6199 29423 6205
rect 30193 6205 30205 6208
rect 30239 6205 30251 6239
rect 30193 6199 30251 6205
rect 28442 6128 28448 6180
rect 28500 6168 28506 6180
rect 30300 6168 30328 6267
rect 28500 6140 30328 6168
rect 28500 6128 28506 6140
rect 23845 6072 24348 6100
rect 25685 6103 25743 6109
rect 23845 6069 23857 6072
rect 23799 6063 23857 6069
rect 25685 6069 25697 6103
rect 25731 6100 25743 6103
rect 27430 6100 27436 6112
rect 25731 6072 27436 6100
rect 25731 6069 25743 6072
rect 25685 6063 25743 6069
rect 27430 6060 27436 6072
rect 27488 6060 27494 6112
rect 29549 6103 29607 6109
rect 29549 6069 29561 6103
rect 29595 6100 29607 6103
rect 29822 6100 29828 6112
rect 29595 6072 29828 6100
rect 29595 6069 29607 6072
rect 29549 6063 29607 6069
rect 29822 6060 29828 6072
rect 29880 6060 29886 6112
rect 1104 6010 30820 6032
rect 1104 5958 4664 6010
rect 4716 5958 4728 6010
rect 4780 5958 4792 6010
rect 4844 5958 4856 6010
rect 4908 5958 4920 6010
rect 4972 5958 12092 6010
rect 12144 5958 12156 6010
rect 12208 5958 12220 6010
rect 12272 5958 12284 6010
rect 12336 5958 12348 6010
rect 12400 5958 19520 6010
rect 19572 5958 19584 6010
rect 19636 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 26948 6010
rect 27000 5958 27012 6010
rect 27064 5958 27076 6010
rect 27128 5958 27140 6010
rect 27192 5958 27204 6010
rect 27256 5958 30820 6010
rect 1104 5936 30820 5958
rect 14277 5899 14335 5905
rect 14277 5865 14289 5899
rect 14323 5896 14335 5899
rect 14642 5896 14648 5908
rect 14323 5868 14648 5896
rect 14323 5865 14335 5868
rect 14277 5859 14335 5865
rect 14642 5856 14648 5868
rect 14700 5856 14706 5908
rect 28537 5899 28595 5905
rect 28537 5865 28549 5899
rect 28583 5896 28595 5899
rect 28902 5896 28908 5908
rect 28583 5868 28908 5896
rect 28583 5865 28595 5868
rect 28537 5859 28595 5865
rect 28902 5856 28908 5868
rect 28960 5856 28966 5908
rect 29086 5856 29092 5908
rect 29144 5856 29150 5908
rect 27890 5828 27896 5840
rect 27172 5800 27896 5828
rect 9582 5720 9588 5772
rect 9640 5760 9646 5772
rect 9640 5732 11836 5760
rect 9640 5720 9646 5732
rect 9398 5652 9404 5704
rect 9456 5692 9462 5704
rect 11808 5701 11836 5732
rect 11974 5720 11980 5772
rect 12032 5760 12038 5772
rect 12069 5763 12127 5769
rect 12069 5760 12081 5763
rect 12032 5732 12081 5760
rect 12032 5720 12038 5732
rect 12069 5729 12081 5732
rect 12115 5729 12127 5763
rect 12069 5723 12127 5729
rect 15657 5763 15715 5769
rect 15657 5729 15669 5763
rect 15703 5760 15715 5763
rect 16850 5760 16856 5772
rect 15703 5732 16856 5760
rect 15703 5729 15715 5732
rect 15657 5723 15715 5729
rect 16850 5720 16856 5732
rect 16908 5720 16914 5772
rect 19702 5720 19708 5772
rect 19760 5720 19766 5772
rect 19978 5720 19984 5772
rect 20036 5720 20042 5772
rect 20438 5720 20444 5772
rect 20496 5760 20502 5772
rect 20806 5760 20812 5772
rect 20496 5732 20812 5760
rect 20496 5720 20502 5732
rect 20806 5720 20812 5732
rect 20864 5760 20870 5772
rect 21450 5760 21456 5772
rect 20864 5732 21456 5760
rect 20864 5720 20870 5732
rect 21450 5720 21456 5732
rect 21508 5720 21514 5772
rect 21726 5720 21732 5772
rect 21784 5720 21790 5772
rect 24302 5720 24308 5772
rect 24360 5760 24366 5772
rect 24581 5763 24639 5769
rect 24581 5760 24593 5763
rect 24360 5732 24593 5760
rect 24360 5720 24366 5732
rect 24581 5729 24593 5732
rect 24627 5729 24639 5763
rect 24581 5723 24639 5729
rect 11333 5695 11391 5701
rect 11333 5692 11345 5695
rect 9456 5664 11345 5692
rect 9456 5652 9462 5664
rect 11333 5661 11345 5664
rect 11379 5661 11391 5695
rect 11333 5655 11391 5661
rect 11793 5695 11851 5701
rect 11793 5661 11805 5695
rect 11839 5692 11851 5695
rect 12434 5692 12440 5704
rect 11839 5664 12440 5692
rect 11839 5661 11851 5664
rect 11793 5655 11851 5661
rect 12434 5652 12440 5664
rect 12492 5652 12498 5704
rect 19613 5695 19671 5701
rect 19613 5661 19625 5695
rect 19659 5661 19671 5695
rect 19613 5655 19671 5661
rect 15412 5627 15470 5633
rect 15412 5593 15424 5627
rect 15458 5624 15470 5627
rect 19426 5624 19432 5636
rect 15458 5596 19432 5624
rect 15458 5593 15470 5596
rect 15412 5587 15470 5593
rect 19426 5584 19432 5596
rect 19484 5584 19490 5636
rect 17954 5516 17960 5568
rect 18012 5556 18018 5568
rect 19628 5556 19656 5655
rect 22830 5652 22836 5704
rect 22888 5652 22894 5704
rect 25958 5652 25964 5704
rect 26016 5692 26022 5704
rect 26697 5695 26755 5701
rect 26697 5692 26709 5695
rect 26016 5664 26709 5692
rect 26016 5652 26022 5664
rect 26697 5661 26709 5664
rect 26743 5661 26755 5695
rect 26697 5655 26755 5661
rect 27065 5695 27123 5701
rect 27065 5661 27077 5695
rect 27111 5692 27123 5695
rect 27172 5692 27200 5800
rect 27890 5788 27896 5800
rect 27948 5788 27954 5840
rect 27525 5763 27583 5769
rect 27525 5729 27537 5763
rect 27571 5760 27583 5763
rect 28718 5760 28724 5772
rect 27571 5732 28724 5760
rect 27571 5729 27583 5732
rect 27525 5723 27583 5729
rect 28718 5720 28724 5732
rect 28776 5720 28782 5772
rect 30101 5763 30159 5769
rect 30101 5729 30113 5763
rect 30147 5760 30159 5763
rect 31018 5760 31024 5772
rect 30147 5732 31024 5760
rect 30147 5729 30159 5732
rect 30101 5723 30159 5729
rect 31018 5720 31024 5732
rect 31076 5720 31082 5772
rect 27111 5664 27200 5692
rect 27249 5695 27307 5701
rect 27111 5661 27123 5664
rect 27065 5655 27123 5661
rect 27249 5661 27261 5695
rect 27295 5692 27307 5695
rect 27338 5692 27344 5704
rect 27295 5664 27344 5692
rect 27295 5661 27307 5664
rect 27249 5655 27307 5661
rect 24826 5627 24884 5633
rect 24826 5624 24838 5627
rect 23216 5596 24838 5624
rect 23216 5565 23244 5596
rect 24826 5593 24838 5596
rect 24872 5593 24884 5627
rect 27264 5624 27292 5655
rect 27338 5652 27344 5664
rect 27396 5652 27402 5704
rect 27433 5695 27491 5701
rect 27433 5661 27445 5695
rect 27479 5692 27491 5695
rect 27706 5692 27712 5704
rect 27479 5664 27712 5692
rect 27479 5661 27491 5664
rect 27433 5655 27491 5661
rect 27706 5652 27712 5664
rect 27764 5692 27770 5704
rect 27985 5695 28043 5701
rect 27985 5692 27997 5695
rect 27764 5664 27997 5692
rect 27764 5652 27770 5664
rect 27985 5661 27997 5664
rect 28031 5661 28043 5695
rect 28261 5695 28319 5701
rect 28261 5692 28273 5695
rect 27985 5655 28043 5661
rect 28092 5664 28273 5692
rect 24826 5587 24884 5593
rect 26206 5596 27292 5624
rect 23201 5559 23259 5565
rect 23201 5556 23213 5559
rect 18012 5528 23213 5556
rect 18012 5516 18018 5528
rect 23201 5525 23213 5528
rect 23247 5525 23259 5559
rect 23201 5519 23259 5525
rect 25961 5559 26019 5565
rect 25961 5525 25973 5559
rect 26007 5556 26019 5559
rect 26206 5556 26234 5596
rect 27890 5584 27896 5636
rect 27948 5624 27954 5636
rect 28092 5624 28120 5664
rect 28261 5661 28273 5664
rect 28307 5661 28319 5695
rect 28261 5655 28319 5661
rect 28350 5652 28356 5704
rect 28408 5692 28414 5704
rect 28997 5695 29055 5701
rect 28997 5692 29009 5695
rect 28408 5664 29009 5692
rect 28408 5652 28414 5664
rect 28997 5661 29009 5664
rect 29043 5661 29055 5695
rect 28997 5655 29055 5661
rect 29822 5652 29828 5704
rect 29880 5652 29886 5704
rect 27948 5596 28120 5624
rect 28169 5627 28227 5633
rect 27948 5584 27954 5596
rect 28169 5593 28181 5627
rect 28215 5593 28227 5627
rect 28169 5587 28227 5593
rect 26007 5528 26234 5556
rect 26007 5525 26019 5528
rect 25961 5519 26019 5525
rect 27430 5516 27436 5568
rect 27488 5556 27494 5568
rect 28184 5556 28212 5587
rect 27488 5528 28212 5556
rect 27488 5516 27494 5528
rect 1104 5466 30976 5488
rect 1104 5414 8378 5466
rect 8430 5414 8442 5466
rect 8494 5414 8506 5466
rect 8558 5414 8570 5466
rect 8622 5414 8634 5466
rect 8686 5414 15806 5466
rect 15858 5414 15870 5466
rect 15922 5414 15934 5466
rect 15986 5414 15998 5466
rect 16050 5414 16062 5466
rect 16114 5414 23234 5466
rect 23286 5414 23298 5466
rect 23350 5414 23362 5466
rect 23414 5414 23426 5466
rect 23478 5414 23490 5466
rect 23542 5414 30662 5466
rect 30714 5414 30726 5466
rect 30778 5414 30790 5466
rect 30842 5414 30854 5466
rect 30906 5414 30918 5466
rect 30970 5414 30976 5466
rect 1104 5392 30976 5414
rect 18325 5355 18383 5361
rect 18325 5321 18337 5355
rect 18371 5321 18383 5355
rect 18325 5315 18383 5321
rect 18340 5284 18368 5315
rect 19702 5312 19708 5364
rect 19760 5352 19766 5364
rect 20165 5355 20223 5361
rect 20165 5352 20177 5355
rect 19760 5324 20177 5352
rect 19760 5312 19766 5324
rect 20165 5321 20177 5324
rect 20211 5321 20223 5355
rect 20165 5315 20223 5321
rect 27617 5355 27675 5361
rect 27617 5321 27629 5355
rect 27663 5352 27675 5355
rect 27890 5352 27896 5364
rect 27663 5324 27896 5352
rect 27663 5321 27675 5324
rect 27617 5315 27675 5321
rect 27890 5312 27896 5324
rect 27948 5312 27954 5364
rect 19030 5287 19088 5293
rect 19030 5284 19042 5287
rect 16960 5256 17356 5284
rect 18340 5256 19042 5284
rect 14113 5219 14171 5225
rect 14113 5185 14125 5219
rect 14159 5216 14171 5219
rect 14550 5216 14556 5228
rect 14159 5188 14556 5216
rect 14159 5185 14171 5188
rect 14113 5179 14171 5185
rect 14550 5176 14556 5188
rect 14608 5176 14614 5228
rect 16960 5225 16988 5256
rect 17218 5225 17224 5228
rect 16945 5219 17003 5225
rect 16945 5185 16957 5219
rect 16991 5185 17003 5219
rect 16945 5179 17003 5185
rect 17212 5179 17224 5225
rect 17218 5176 17224 5179
rect 17276 5176 17282 5228
rect 17328 5216 17356 5256
rect 19030 5253 19042 5256
rect 19076 5253 19088 5287
rect 19030 5247 19088 5253
rect 27525 5287 27583 5293
rect 27525 5253 27537 5287
rect 27571 5284 27583 5287
rect 28350 5284 28356 5296
rect 27571 5256 28356 5284
rect 27571 5253 27583 5256
rect 27525 5247 27583 5253
rect 28350 5244 28356 5256
rect 28408 5244 28414 5296
rect 18598 5216 18604 5228
rect 17328 5188 18604 5216
rect 18598 5176 18604 5188
rect 18656 5216 18662 5228
rect 18785 5219 18843 5225
rect 18785 5216 18797 5219
rect 18656 5188 18797 5216
rect 18656 5176 18662 5188
rect 18785 5185 18797 5188
rect 18831 5185 18843 5219
rect 18785 5179 18843 5185
rect 27430 5176 27436 5228
rect 27488 5176 27494 5228
rect 27706 5176 27712 5228
rect 27764 5216 27770 5228
rect 27801 5219 27859 5225
rect 27801 5216 27813 5219
rect 27764 5188 27813 5216
rect 27764 5176 27770 5188
rect 27801 5185 27813 5188
rect 27847 5185 27859 5219
rect 27801 5179 27859 5185
rect 28718 5176 28724 5228
rect 28776 5176 28782 5228
rect 28810 5176 28816 5228
rect 28868 5216 28874 5228
rect 28905 5219 28963 5225
rect 28905 5216 28917 5219
rect 28868 5188 28917 5216
rect 28868 5176 28874 5188
rect 28905 5185 28917 5188
rect 28951 5185 28963 5219
rect 28905 5179 28963 5185
rect 14366 5108 14372 5160
rect 14424 5108 14430 5160
rect 27709 5083 27767 5089
rect 27709 5049 27721 5083
rect 27755 5080 27767 5083
rect 28442 5080 28448 5092
rect 27755 5052 28448 5080
rect 27755 5049 27767 5052
rect 27709 5043 27767 5049
rect 28442 5040 28448 5052
rect 28500 5040 28506 5092
rect 12989 5015 13047 5021
rect 12989 4981 13001 5015
rect 13035 5012 13047 5015
rect 13998 5012 14004 5024
rect 13035 4984 14004 5012
rect 13035 4981 13047 4984
rect 12989 4975 13047 4981
rect 13998 4972 14004 4984
rect 14056 4972 14062 5024
rect 28718 4972 28724 5024
rect 28776 4972 28782 5024
rect 1104 4922 30820 4944
rect 1104 4870 4664 4922
rect 4716 4870 4728 4922
rect 4780 4870 4792 4922
rect 4844 4870 4856 4922
rect 4908 4870 4920 4922
rect 4972 4870 12092 4922
rect 12144 4870 12156 4922
rect 12208 4870 12220 4922
rect 12272 4870 12284 4922
rect 12336 4870 12348 4922
rect 12400 4870 19520 4922
rect 19572 4870 19584 4922
rect 19636 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 26948 4922
rect 27000 4870 27012 4922
rect 27064 4870 27076 4922
rect 27128 4870 27140 4922
rect 27192 4870 27204 4922
rect 27256 4870 30820 4922
rect 1104 4848 30820 4870
rect 17218 4768 17224 4820
rect 17276 4768 17282 4820
rect 19426 4768 19432 4820
rect 19484 4768 19490 4820
rect 14366 4700 14372 4752
rect 14424 4740 14430 4752
rect 16761 4743 16819 4749
rect 14424 4712 14780 4740
rect 14424 4700 14430 4712
rect 14642 4632 14648 4684
rect 14700 4632 14706 4684
rect 14550 4564 14556 4616
rect 14608 4564 14614 4616
rect 14752 4604 14780 4712
rect 16761 4709 16773 4743
rect 16807 4709 16819 4743
rect 16761 4703 16819 4709
rect 14921 4675 14979 4681
rect 14921 4641 14933 4675
rect 14967 4672 14979 4675
rect 16776 4672 16804 4703
rect 17497 4675 17555 4681
rect 17497 4672 17509 4675
rect 14967 4644 15516 4672
rect 16776 4644 17509 4672
rect 14967 4641 14979 4644
rect 14921 4635 14979 4641
rect 15381 4607 15439 4613
rect 15381 4604 15393 4607
rect 14752 4576 15393 4604
rect 15381 4573 15393 4576
rect 15427 4573 15439 4607
rect 15488 4604 15516 4644
rect 17497 4641 17509 4644
rect 17543 4641 17555 4675
rect 17497 4635 17555 4641
rect 20806 4632 20812 4684
rect 20864 4632 20870 4684
rect 15637 4607 15695 4613
rect 15637 4604 15649 4607
rect 15488 4576 15649 4604
rect 15381 4567 15439 4573
rect 15637 4573 15649 4576
rect 15683 4573 15695 4607
rect 17589 4607 17647 4613
rect 17589 4604 17601 4607
rect 15637 4567 15695 4573
rect 16546 4576 17601 4604
rect 14568 4536 14596 4564
rect 16546 4536 16574 4576
rect 17589 4573 17601 4576
rect 17635 4604 17647 4607
rect 17954 4604 17960 4616
rect 17635 4576 17960 4604
rect 17635 4573 17647 4576
rect 17589 4567 17647 4573
rect 17954 4564 17960 4576
rect 18012 4564 18018 4616
rect 19978 4564 19984 4616
rect 20036 4604 20042 4616
rect 20542 4607 20600 4613
rect 20542 4604 20554 4607
rect 20036 4576 20554 4604
rect 20036 4564 20042 4576
rect 20542 4573 20554 4576
rect 20588 4573 20600 4607
rect 20542 4567 20600 4573
rect 14568 4508 16574 4536
rect 1104 4378 30976 4400
rect 1104 4326 8378 4378
rect 8430 4326 8442 4378
rect 8494 4326 8506 4378
rect 8558 4326 8570 4378
rect 8622 4326 8634 4378
rect 8686 4326 15806 4378
rect 15858 4326 15870 4378
rect 15922 4326 15934 4378
rect 15986 4326 15998 4378
rect 16050 4326 16062 4378
rect 16114 4326 23234 4378
rect 23286 4326 23298 4378
rect 23350 4326 23362 4378
rect 23414 4326 23426 4378
rect 23478 4326 23490 4378
rect 23542 4326 30662 4378
rect 30714 4326 30726 4378
rect 30778 4326 30790 4378
rect 30842 4326 30854 4378
rect 30906 4326 30918 4378
rect 30970 4326 30976 4378
rect 1104 4304 30976 4326
rect 14642 4224 14648 4276
rect 14700 4264 14706 4276
rect 15105 4267 15163 4273
rect 15105 4264 15117 4267
rect 14700 4236 15117 4264
rect 14700 4224 14706 4236
rect 15105 4233 15117 4236
rect 15151 4233 15163 4267
rect 15105 4227 15163 4233
rect 14366 4196 14372 4208
rect 13832 4168 14372 4196
rect 13725 4131 13783 4137
rect 13725 4097 13737 4131
rect 13771 4128 13783 4131
rect 13832 4128 13860 4168
rect 14366 4156 14372 4168
rect 14424 4156 14430 4208
rect 13998 4137 14004 4140
rect 13992 4128 14004 4137
rect 13771 4100 13860 4128
rect 13959 4100 14004 4128
rect 13771 4097 13783 4100
rect 13725 4091 13783 4097
rect 13992 4091 14004 4100
rect 13998 4088 14004 4091
rect 14056 4088 14062 4140
rect 1104 3834 30820 3856
rect 1104 3782 4664 3834
rect 4716 3782 4728 3834
rect 4780 3782 4792 3834
rect 4844 3782 4856 3834
rect 4908 3782 4920 3834
rect 4972 3782 12092 3834
rect 12144 3782 12156 3834
rect 12208 3782 12220 3834
rect 12272 3782 12284 3834
rect 12336 3782 12348 3834
rect 12400 3782 19520 3834
rect 19572 3782 19584 3834
rect 19636 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 26948 3834
rect 27000 3782 27012 3834
rect 27064 3782 27076 3834
rect 27128 3782 27140 3834
rect 27192 3782 27204 3834
rect 27256 3782 30820 3834
rect 1104 3760 30820 3782
rect 1104 3290 30976 3312
rect 1104 3238 8378 3290
rect 8430 3238 8442 3290
rect 8494 3238 8506 3290
rect 8558 3238 8570 3290
rect 8622 3238 8634 3290
rect 8686 3238 15806 3290
rect 15858 3238 15870 3290
rect 15922 3238 15934 3290
rect 15986 3238 15998 3290
rect 16050 3238 16062 3290
rect 16114 3238 23234 3290
rect 23286 3238 23298 3290
rect 23350 3238 23362 3290
rect 23414 3238 23426 3290
rect 23478 3238 23490 3290
rect 23542 3238 30662 3290
rect 30714 3238 30726 3290
rect 30778 3238 30790 3290
rect 30842 3238 30854 3290
rect 30906 3238 30918 3290
rect 30970 3238 30976 3290
rect 1104 3216 30976 3238
rect 1104 2746 30820 2768
rect 1104 2694 4664 2746
rect 4716 2694 4728 2746
rect 4780 2694 4792 2746
rect 4844 2694 4856 2746
rect 4908 2694 4920 2746
rect 4972 2694 12092 2746
rect 12144 2694 12156 2746
rect 12208 2694 12220 2746
rect 12272 2694 12284 2746
rect 12336 2694 12348 2746
rect 12400 2694 19520 2746
rect 19572 2694 19584 2746
rect 19636 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 26948 2746
rect 27000 2694 27012 2746
rect 27064 2694 27076 2746
rect 27128 2694 27140 2746
rect 27192 2694 27204 2746
rect 27256 2694 30820 2746
rect 1104 2672 30820 2694
rect 28718 2388 28724 2440
rect 28776 2428 28782 2440
rect 29825 2431 29883 2437
rect 29825 2428 29837 2431
rect 28776 2400 29837 2428
rect 28776 2388 28782 2400
rect 29825 2397 29837 2400
rect 29871 2397 29883 2431
rect 29825 2391 29883 2397
rect 30101 2363 30159 2369
rect 30101 2329 30113 2363
rect 30147 2360 30159 2363
rect 31018 2360 31024 2372
rect 30147 2332 31024 2360
rect 30147 2329 30159 2332
rect 30101 2323 30159 2329
rect 31018 2320 31024 2332
rect 31076 2320 31082 2372
rect 1104 2202 30976 2224
rect 1104 2150 8378 2202
rect 8430 2150 8442 2202
rect 8494 2150 8506 2202
rect 8558 2150 8570 2202
rect 8622 2150 8634 2202
rect 8686 2150 15806 2202
rect 15858 2150 15870 2202
rect 15922 2150 15934 2202
rect 15986 2150 15998 2202
rect 16050 2150 16062 2202
rect 16114 2150 23234 2202
rect 23286 2150 23298 2202
rect 23350 2150 23362 2202
rect 23414 2150 23426 2202
rect 23478 2150 23490 2202
rect 23542 2150 30662 2202
rect 30714 2150 30726 2202
rect 30778 2150 30790 2202
rect 30842 2150 30854 2202
rect 30906 2150 30918 2202
rect 30970 2150 30976 2202
rect 1104 2128 30976 2150
<< via1 >>
rect 8378 29350 8430 29402
rect 8442 29350 8494 29402
rect 8506 29350 8558 29402
rect 8570 29350 8622 29402
rect 8634 29350 8686 29402
rect 15806 29350 15858 29402
rect 15870 29350 15922 29402
rect 15934 29350 15986 29402
rect 15998 29350 16050 29402
rect 16062 29350 16114 29402
rect 23234 29350 23286 29402
rect 23298 29350 23350 29402
rect 23362 29350 23414 29402
rect 23426 29350 23478 29402
rect 23490 29350 23542 29402
rect 30662 29350 30714 29402
rect 30726 29350 30778 29402
rect 30790 29350 30842 29402
rect 30854 29350 30906 29402
rect 30918 29350 30970 29402
rect 6092 29180 6144 29232
rect 15384 29180 15436 29232
rect 18144 29223 18196 29232
rect 18144 29189 18153 29223
rect 18153 29189 18187 29223
rect 18187 29189 18196 29223
rect 18144 29180 18196 29189
rect 31024 29180 31076 29232
rect 3240 29112 3292 29164
rect 3056 29044 3108 29096
rect 10232 29155 10284 29164
rect 10232 29121 10241 29155
rect 10241 29121 10275 29155
rect 10275 29121 10284 29155
rect 10232 29112 10284 29121
rect 14004 29112 14056 29164
rect 22008 29155 22060 29164
rect 22008 29121 22017 29155
rect 22017 29121 22051 29155
rect 22051 29121 22060 29155
rect 22008 29112 22060 29121
rect 25964 29155 26016 29164
rect 25964 29121 25973 29155
rect 25973 29121 26007 29155
rect 26007 29121 26016 29155
rect 25964 29112 26016 29121
rect 29736 29112 29788 29164
rect 14464 29044 14516 29096
rect 28540 29087 28592 29096
rect 28540 29053 28549 29087
rect 28549 29053 28583 29087
rect 28583 29053 28592 29087
rect 28540 29044 28592 29053
rect 29000 29044 29052 29096
rect 4528 28976 4580 29028
rect 7196 28976 7248 29028
rect 22192 29019 22244 29028
rect 22192 28985 22201 29019
rect 22201 28985 22235 29019
rect 22235 28985 22244 29019
rect 22192 28976 22244 28985
rect 25688 28976 25740 29028
rect 18144 28908 18196 28960
rect 4664 28806 4716 28858
rect 4728 28806 4780 28858
rect 4792 28806 4844 28858
rect 4856 28806 4908 28858
rect 4920 28806 4972 28858
rect 12092 28806 12144 28858
rect 12156 28806 12208 28858
rect 12220 28806 12272 28858
rect 12284 28806 12336 28858
rect 12348 28806 12400 28858
rect 19520 28806 19572 28858
rect 19584 28806 19636 28858
rect 19648 28806 19700 28858
rect 19712 28806 19764 28858
rect 19776 28806 19828 28858
rect 26948 28806 27000 28858
rect 27012 28806 27064 28858
rect 27076 28806 27128 28858
rect 27140 28806 27192 28858
rect 27204 28806 27256 28858
rect 2136 28704 2188 28756
rect 3516 28704 3568 28756
rect 3148 28679 3200 28688
rect 3148 28645 3157 28679
rect 3157 28645 3191 28679
rect 3191 28645 3200 28679
rect 3148 28636 3200 28645
rect 3240 28500 3292 28552
rect 3884 28500 3936 28552
rect 7196 28500 7248 28552
rect 8760 28500 8812 28552
rect 10324 28543 10376 28552
rect 10324 28509 10333 28543
rect 10333 28509 10367 28543
rect 10367 28509 10376 28543
rect 10324 28500 10376 28509
rect 11060 28543 11112 28552
rect 11060 28509 11069 28543
rect 11069 28509 11103 28543
rect 11103 28509 11112 28543
rect 11060 28500 11112 28509
rect 11704 28500 11756 28552
rect 12716 28500 12768 28552
rect 13728 28500 13780 28552
rect 14924 28500 14976 28552
rect 18144 28500 18196 28552
rect 20720 28500 20772 28552
rect 3056 28432 3108 28484
rect 11796 28475 11848 28484
rect 11796 28441 11805 28475
rect 11805 28441 11839 28475
rect 11839 28441 11848 28475
rect 11796 28432 11848 28441
rect 21824 28500 21876 28552
rect 22836 28500 22888 28552
rect 26424 28500 26476 28552
rect 27896 28500 27948 28552
rect 23572 28432 23624 28484
rect 27620 28432 27672 28484
rect 7012 28364 7064 28416
rect 8300 28407 8352 28416
rect 8300 28373 8309 28407
rect 8309 28373 8343 28407
rect 8343 28373 8352 28407
rect 8300 28364 8352 28373
rect 8852 28364 8904 28416
rect 10876 28364 10928 28416
rect 12072 28364 12124 28416
rect 15292 28364 15344 28416
rect 16212 28364 16264 28416
rect 18604 28364 18656 28416
rect 20904 28407 20956 28416
rect 20904 28373 20913 28407
rect 20913 28373 20947 28407
rect 20947 28373 20956 28407
rect 20904 28364 20956 28373
rect 22376 28364 22428 28416
rect 23756 28407 23808 28416
rect 23756 28373 23765 28407
rect 23765 28373 23799 28407
rect 23799 28373 23808 28407
rect 23756 28364 23808 28373
rect 27436 28364 27488 28416
rect 29184 28407 29236 28416
rect 29184 28373 29193 28407
rect 29193 28373 29227 28407
rect 29227 28373 29236 28407
rect 29184 28364 29236 28373
rect 8378 28262 8430 28314
rect 8442 28262 8494 28314
rect 8506 28262 8558 28314
rect 8570 28262 8622 28314
rect 8634 28262 8686 28314
rect 15806 28262 15858 28314
rect 15870 28262 15922 28314
rect 15934 28262 15986 28314
rect 15998 28262 16050 28314
rect 16062 28262 16114 28314
rect 23234 28262 23286 28314
rect 23298 28262 23350 28314
rect 23362 28262 23414 28314
rect 23426 28262 23478 28314
rect 23490 28262 23542 28314
rect 30662 28262 30714 28314
rect 30726 28262 30778 28314
rect 30790 28262 30842 28314
rect 30854 28262 30906 28314
rect 30918 28262 30970 28314
rect 12716 28160 12768 28212
rect 13820 28203 13872 28212
rect 13820 28169 13829 28203
rect 13829 28169 13863 28203
rect 13863 28169 13872 28203
rect 13820 28160 13872 28169
rect 14924 28160 14976 28212
rect 15292 28160 15344 28212
rect 2872 28092 2924 28144
rect 2964 28067 3016 28076
rect 2964 28033 2998 28067
rect 2998 28033 3016 28067
rect 2964 28024 3016 28033
rect 4528 28092 4580 28144
rect 8852 28092 8904 28144
rect 6920 28024 6972 28076
rect 8300 28067 8352 28076
rect 8300 28033 8309 28067
rect 8309 28033 8343 28067
rect 8343 28033 8352 28067
rect 8300 28024 8352 28033
rect 9680 28024 9732 28076
rect 13360 28092 13412 28144
rect 15476 28092 15528 28144
rect 12072 28067 12124 28076
rect 12072 28033 12081 28067
rect 12081 28033 12115 28067
rect 12115 28033 12124 28067
rect 12072 28024 12124 28033
rect 16212 28067 16264 28076
rect 16212 28033 16221 28067
rect 16221 28033 16255 28067
rect 16255 28033 16264 28067
rect 16212 28024 16264 28033
rect 18788 28160 18840 28212
rect 23572 28160 23624 28212
rect 18880 28092 18932 28144
rect 23756 28092 23808 28144
rect 27436 28135 27488 28144
rect 27436 28101 27445 28135
rect 27445 28101 27479 28135
rect 27479 28101 27488 28135
rect 27436 28092 27488 28101
rect 28172 28092 28224 28144
rect 20812 28067 20864 28076
rect 20812 28033 20821 28067
rect 20821 28033 20855 28067
rect 20855 28033 20864 28067
rect 20812 28024 20864 28033
rect 21088 28067 21140 28076
rect 21088 28033 21097 28067
rect 21097 28033 21131 28067
rect 21131 28033 21140 28067
rect 21088 28024 21140 28033
rect 21824 28024 21876 28076
rect 29460 28067 29512 28076
rect 29460 28033 29469 28067
rect 29469 28033 29503 28067
rect 29503 28033 29512 28067
rect 29460 28024 29512 28033
rect 3976 27956 4028 28008
rect 7380 27956 7432 28008
rect 7656 27956 7708 28008
rect 13636 27956 13688 28008
rect 19892 27999 19944 28008
rect 19892 27965 19901 27999
rect 19901 27965 19935 27999
rect 19935 27965 19944 27999
rect 19892 27956 19944 27965
rect 21364 27999 21416 28008
rect 21364 27965 21373 27999
rect 21373 27965 21407 27999
rect 21407 27965 21416 27999
rect 21364 27956 21416 27965
rect 10324 27888 10376 27940
rect 11888 27888 11940 27940
rect 13728 27888 13780 27940
rect 3884 27820 3936 27872
rect 5908 27863 5960 27872
rect 5908 27829 5917 27863
rect 5917 27829 5951 27863
rect 5951 27829 5960 27863
rect 5908 27820 5960 27829
rect 11152 27820 11204 27872
rect 22744 27999 22796 28008
rect 22744 27965 22753 27999
rect 22753 27965 22787 27999
rect 22787 27965 22796 27999
rect 22744 27956 22796 27965
rect 26608 27956 26660 28008
rect 23480 27820 23532 27872
rect 28908 27863 28960 27872
rect 28908 27829 28917 27863
rect 28917 27829 28951 27863
rect 28951 27829 28960 27863
rect 28908 27820 28960 27829
rect 29920 27820 29972 27872
rect 4664 27718 4716 27770
rect 4728 27718 4780 27770
rect 4792 27718 4844 27770
rect 4856 27718 4908 27770
rect 4920 27718 4972 27770
rect 12092 27718 12144 27770
rect 12156 27718 12208 27770
rect 12220 27718 12272 27770
rect 12284 27718 12336 27770
rect 12348 27718 12400 27770
rect 19520 27718 19572 27770
rect 19584 27718 19636 27770
rect 19648 27718 19700 27770
rect 19712 27718 19764 27770
rect 19776 27718 19828 27770
rect 26948 27718 27000 27770
rect 27012 27718 27064 27770
rect 27076 27718 27128 27770
rect 27140 27718 27192 27770
rect 27204 27718 27256 27770
rect 2964 27659 3016 27668
rect 2964 27625 2973 27659
rect 2973 27625 3007 27659
rect 3007 27625 3016 27659
rect 2964 27616 3016 27625
rect 3884 27616 3936 27668
rect 7012 27616 7064 27668
rect 10968 27616 11020 27668
rect 11152 27659 11204 27668
rect 11152 27625 11182 27659
rect 11182 27625 11204 27659
rect 11152 27616 11204 27625
rect 19892 27616 19944 27668
rect 20904 27616 20956 27668
rect 22744 27616 22796 27668
rect 26608 27659 26660 27668
rect 26608 27625 26617 27659
rect 26617 27625 26651 27659
rect 26651 27625 26660 27659
rect 26608 27616 26660 27625
rect 3240 27480 3292 27532
rect 3884 27480 3936 27532
rect 3976 27523 4028 27532
rect 3976 27489 3985 27523
rect 3985 27489 4019 27523
rect 4019 27489 4028 27523
rect 3976 27480 4028 27489
rect 5816 27591 5868 27600
rect 5816 27557 5825 27591
rect 5825 27557 5859 27591
rect 5859 27557 5868 27591
rect 5816 27548 5868 27557
rect 3148 27455 3200 27464
rect 3148 27421 3157 27455
rect 3157 27421 3191 27455
rect 3191 27421 3200 27455
rect 3148 27412 3200 27421
rect 5908 27412 5960 27464
rect 7380 27480 7432 27532
rect 9680 27548 9732 27600
rect 13636 27591 13688 27600
rect 13636 27557 13645 27591
rect 13645 27557 13679 27591
rect 13679 27557 13688 27591
rect 13636 27548 13688 27557
rect 6644 27455 6696 27464
rect 6644 27421 6653 27455
rect 6653 27421 6687 27455
rect 6687 27421 6696 27455
rect 6644 27412 6696 27421
rect 11704 27480 11756 27532
rect 15476 27523 15528 27532
rect 15476 27489 15485 27523
rect 15485 27489 15519 27523
rect 15519 27489 15528 27523
rect 15476 27480 15528 27489
rect 10876 27455 10928 27464
rect 10876 27421 10885 27455
rect 10885 27421 10919 27455
rect 10919 27421 10928 27455
rect 10876 27412 10928 27421
rect 13820 27412 13872 27464
rect 14096 27412 14148 27464
rect 14648 27412 14700 27464
rect 20812 27548 20864 27600
rect 23480 27548 23532 27600
rect 23664 27548 23716 27600
rect 29000 27548 29052 27600
rect 18880 27523 18932 27532
rect 18880 27489 18889 27523
rect 18889 27489 18923 27523
rect 18923 27489 18932 27523
rect 18880 27480 18932 27489
rect 21088 27480 21140 27532
rect 22376 27523 22428 27532
rect 22376 27489 22385 27523
rect 22385 27489 22419 27523
rect 22419 27489 22428 27523
rect 22376 27480 22428 27489
rect 25872 27480 25924 27532
rect 26056 27523 26108 27532
rect 26056 27489 26065 27523
rect 26065 27489 26099 27523
rect 26099 27489 26108 27523
rect 26056 27480 26108 27489
rect 28172 27523 28224 27532
rect 28172 27489 28181 27523
rect 28181 27489 28215 27523
rect 28215 27489 28224 27523
rect 28172 27480 28224 27489
rect 2320 27319 2372 27328
rect 2320 27285 2345 27319
rect 2345 27285 2372 27319
rect 2320 27276 2372 27285
rect 3424 27276 3476 27328
rect 3608 27344 3660 27396
rect 7656 27344 7708 27396
rect 11796 27344 11848 27396
rect 8760 27276 8812 27328
rect 9312 27276 9364 27328
rect 11060 27276 11112 27328
rect 12716 27276 12768 27328
rect 23572 27412 23624 27464
rect 21364 27344 21416 27396
rect 22928 27344 22980 27396
rect 26424 27412 26476 27464
rect 26608 27412 26660 27464
rect 27620 27455 27672 27464
rect 27620 27421 27629 27455
rect 27629 27421 27663 27455
rect 27663 27421 27672 27455
rect 27620 27412 27672 27421
rect 27896 27455 27948 27464
rect 27896 27421 27905 27455
rect 27905 27421 27939 27455
rect 27939 27421 27948 27455
rect 27896 27412 27948 27421
rect 26148 27344 26200 27396
rect 28908 27412 28960 27464
rect 20720 27276 20772 27328
rect 20812 27276 20864 27328
rect 27620 27276 27672 27328
rect 30196 27276 30248 27328
rect 8378 27174 8430 27226
rect 8442 27174 8494 27226
rect 8506 27174 8558 27226
rect 8570 27174 8622 27226
rect 8634 27174 8686 27226
rect 15806 27174 15858 27226
rect 15870 27174 15922 27226
rect 15934 27174 15986 27226
rect 15998 27174 16050 27226
rect 16062 27174 16114 27226
rect 23234 27174 23286 27226
rect 23298 27174 23350 27226
rect 23362 27174 23414 27226
rect 23426 27174 23478 27226
rect 23490 27174 23542 27226
rect 30662 27174 30714 27226
rect 30726 27174 30778 27226
rect 30790 27174 30842 27226
rect 30854 27174 30906 27226
rect 30918 27174 30970 27226
rect 3332 27072 3384 27124
rect 5816 27072 5868 27124
rect 6644 27072 6696 27124
rect 23664 27072 23716 27124
rect 11704 27004 11756 27056
rect 2872 26979 2924 26988
rect 2872 26945 2881 26979
rect 2881 26945 2915 26979
rect 2915 26945 2924 26979
rect 2872 26936 2924 26945
rect 3424 26936 3476 26988
rect 4988 26979 5040 26988
rect 4988 26945 4997 26979
rect 4997 26945 5031 26979
rect 5031 26945 5040 26979
rect 4988 26936 5040 26945
rect 8300 26936 8352 26988
rect 11888 26979 11940 26988
rect 11888 26945 11897 26979
rect 11897 26945 11931 26979
rect 11931 26945 11940 26979
rect 11888 26936 11940 26945
rect 13360 27047 13412 27056
rect 13360 27013 13369 27047
rect 13369 27013 13403 27047
rect 13403 27013 13412 27047
rect 13360 27004 13412 27013
rect 14648 27004 14700 27056
rect 23572 27004 23624 27056
rect 14096 26979 14148 26988
rect 14096 26945 14105 26979
rect 14105 26945 14139 26979
rect 14139 26945 14148 26979
rect 14096 26936 14148 26945
rect 16212 26936 16264 26988
rect 18604 26936 18656 26988
rect 20076 26936 20128 26988
rect 29184 27004 29236 27056
rect 29920 27047 29972 27056
rect 29920 27013 29929 27047
rect 29929 27013 29963 27047
rect 29963 27013 29972 27047
rect 29920 27004 29972 27013
rect 24952 26979 25004 26988
rect 24952 26945 24986 26979
rect 24986 26945 25004 26979
rect 24952 26936 25004 26945
rect 30196 26979 30248 26988
rect 30196 26945 30205 26979
rect 30205 26945 30239 26979
rect 30239 26945 30248 26979
rect 30196 26936 30248 26945
rect 11796 26911 11848 26920
rect 11796 26877 11805 26911
rect 11805 26877 11839 26911
rect 11839 26877 11848 26911
rect 11796 26868 11848 26877
rect 16580 26868 16632 26920
rect 18052 26911 18104 26920
rect 18052 26877 18061 26911
rect 18061 26877 18095 26911
rect 18095 26877 18104 26911
rect 18052 26868 18104 26877
rect 23112 26868 23164 26920
rect 24584 26868 24636 26920
rect 4252 26843 4304 26852
rect 4252 26809 4261 26843
rect 4261 26809 4295 26843
rect 4295 26809 4304 26843
rect 4252 26800 4304 26809
rect 25872 26800 25924 26852
rect 6736 26775 6788 26784
rect 6736 26741 6745 26775
rect 6745 26741 6779 26775
rect 6779 26741 6788 26775
rect 6736 26732 6788 26741
rect 12900 26732 12952 26784
rect 15016 26732 15068 26784
rect 25964 26732 26016 26784
rect 26148 26732 26200 26784
rect 29460 26732 29512 26784
rect 4664 26630 4716 26682
rect 4728 26630 4780 26682
rect 4792 26630 4844 26682
rect 4856 26630 4908 26682
rect 4920 26630 4972 26682
rect 12092 26630 12144 26682
rect 12156 26630 12208 26682
rect 12220 26630 12272 26682
rect 12284 26630 12336 26682
rect 12348 26630 12400 26682
rect 19520 26630 19572 26682
rect 19584 26630 19636 26682
rect 19648 26630 19700 26682
rect 19712 26630 19764 26682
rect 19776 26630 19828 26682
rect 26948 26630 27000 26682
rect 27012 26630 27064 26682
rect 27076 26630 27128 26682
rect 27140 26630 27192 26682
rect 27204 26630 27256 26682
rect 3608 26528 3660 26580
rect 3884 26528 3936 26580
rect 3332 26503 3384 26512
rect 3332 26469 3341 26503
rect 3341 26469 3375 26503
rect 3375 26469 3384 26503
rect 3332 26460 3384 26469
rect 2320 26392 2372 26444
rect 11796 26528 11848 26580
rect 12164 26528 12216 26580
rect 16212 26528 16264 26580
rect 24952 26528 25004 26580
rect 26056 26571 26108 26580
rect 26056 26537 26065 26571
rect 26065 26537 26099 26571
rect 26099 26537 26108 26571
rect 26056 26528 26108 26537
rect 26148 26528 26200 26580
rect 7380 26460 7432 26512
rect 3424 26367 3476 26376
rect 3424 26333 3433 26367
rect 3433 26333 3467 26367
rect 3467 26333 3476 26367
rect 3424 26324 3476 26333
rect 3792 26324 3844 26376
rect 3056 26256 3108 26308
rect 3976 26256 4028 26308
rect 4252 26367 4304 26376
rect 4252 26333 4261 26367
rect 4261 26333 4295 26367
rect 4295 26333 4304 26367
rect 4252 26324 4304 26333
rect 8024 26435 8076 26444
rect 8024 26401 8033 26435
rect 8033 26401 8067 26435
rect 8067 26401 8076 26435
rect 8024 26392 8076 26401
rect 6920 26324 6972 26376
rect 8300 26324 8352 26376
rect 9312 26367 9364 26376
rect 9312 26333 9321 26367
rect 9321 26333 9355 26367
rect 9355 26333 9364 26367
rect 9312 26324 9364 26333
rect 9680 26435 9732 26444
rect 9680 26401 9689 26435
rect 9689 26401 9723 26435
rect 9723 26401 9732 26435
rect 9680 26392 9732 26401
rect 10232 26324 10284 26376
rect 11152 26367 11204 26376
rect 11152 26333 11161 26367
rect 11161 26333 11195 26367
rect 11195 26333 11204 26367
rect 11152 26324 11204 26333
rect 14556 26435 14608 26444
rect 14556 26401 14565 26435
rect 14565 26401 14599 26435
rect 14599 26401 14608 26435
rect 14556 26392 14608 26401
rect 15016 26435 15068 26444
rect 15016 26401 15025 26435
rect 15025 26401 15059 26435
rect 15059 26401 15068 26435
rect 15016 26392 15068 26401
rect 15200 26392 15252 26444
rect 23112 26460 23164 26512
rect 12992 26324 13044 26376
rect 14924 26367 14976 26376
rect 14924 26333 14933 26367
rect 14933 26333 14967 26367
rect 14967 26333 14976 26367
rect 14924 26324 14976 26333
rect 7288 26299 7340 26308
rect 7288 26265 7297 26299
rect 7297 26265 7331 26299
rect 7331 26265 7340 26299
rect 7288 26256 7340 26265
rect 11704 26256 11756 26308
rect 15660 26256 15712 26308
rect 18788 26367 18840 26376
rect 18788 26333 18797 26367
rect 18797 26333 18831 26367
rect 18831 26333 18840 26367
rect 18788 26324 18840 26333
rect 20812 26392 20864 26444
rect 25872 26460 25924 26512
rect 25412 26435 25464 26444
rect 25412 26401 25421 26435
rect 25421 26401 25455 26435
rect 25455 26401 25464 26435
rect 25412 26392 25464 26401
rect 25964 26392 26016 26444
rect 27620 26392 27672 26444
rect 21088 26324 21140 26376
rect 21824 26367 21876 26376
rect 21824 26333 21833 26367
rect 21833 26333 21867 26367
rect 21867 26333 21876 26367
rect 21824 26324 21876 26333
rect 26332 26367 26384 26376
rect 26332 26333 26341 26367
rect 26341 26333 26375 26367
rect 26375 26333 26384 26367
rect 26332 26324 26384 26333
rect 27896 26324 27948 26376
rect 29920 26367 29972 26376
rect 29920 26333 29929 26367
rect 29929 26333 29963 26367
rect 29963 26333 29972 26367
rect 29920 26324 29972 26333
rect 4160 26188 4212 26240
rect 18420 26188 18472 26240
rect 19432 26231 19484 26240
rect 19432 26197 19441 26231
rect 19441 26197 19475 26231
rect 19475 26197 19484 26231
rect 19432 26188 19484 26197
rect 22284 26256 22336 26308
rect 22008 26188 22060 26240
rect 22192 26188 22244 26240
rect 25504 26256 25556 26308
rect 26056 26299 26108 26308
rect 26056 26265 26065 26299
rect 26065 26265 26099 26299
rect 26099 26265 26108 26299
rect 26056 26256 26108 26265
rect 26608 26256 26660 26308
rect 29184 26231 29236 26240
rect 29184 26197 29193 26231
rect 29193 26197 29227 26231
rect 29227 26197 29236 26231
rect 29184 26188 29236 26197
rect 29828 26231 29880 26240
rect 29828 26197 29837 26231
rect 29837 26197 29871 26231
rect 29871 26197 29880 26231
rect 29828 26188 29880 26197
rect 8378 26086 8430 26138
rect 8442 26086 8494 26138
rect 8506 26086 8558 26138
rect 8570 26086 8622 26138
rect 8634 26086 8686 26138
rect 15806 26086 15858 26138
rect 15870 26086 15922 26138
rect 15934 26086 15986 26138
rect 15998 26086 16050 26138
rect 16062 26086 16114 26138
rect 23234 26086 23286 26138
rect 23298 26086 23350 26138
rect 23362 26086 23414 26138
rect 23426 26086 23478 26138
rect 23490 26086 23542 26138
rect 30662 26086 30714 26138
rect 30726 26086 30778 26138
rect 30790 26086 30842 26138
rect 30854 26086 30906 26138
rect 30918 26086 30970 26138
rect 2872 26027 2924 26036
rect 2872 25993 2881 26027
rect 2881 25993 2915 26027
rect 2915 25993 2924 26027
rect 2872 25984 2924 25993
rect 8300 26027 8352 26036
rect 8300 25993 8309 26027
rect 8309 25993 8343 26027
rect 8343 25993 8352 26027
rect 8300 25984 8352 25993
rect 10232 26027 10284 26036
rect 10232 25993 10241 26027
rect 10241 25993 10275 26027
rect 10275 25993 10284 26027
rect 10232 25984 10284 25993
rect 11704 26027 11756 26036
rect 11704 25993 11713 26027
rect 11713 25993 11747 26027
rect 11747 25993 11756 26027
rect 11704 25984 11756 25993
rect 12164 26027 12216 26036
rect 12164 25993 12173 26027
rect 12173 25993 12207 26027
rect 12207 25993 12216 26027
rect 12164 25984 12216 25993
rect 6736 25916 6788 25968
rect 7288 25916 7340 25968
rect 12900 25959 12952 25968
rect 12900 25925 12909 25959
rect 12909 25925 12943 25959
rect 12943 25925 12952 25959
rect 12900 25916 12952 25925
rect 22284 26027 22336 26036
rect 22284 25993 22293 26027
rect 22293 25993 22327 26027
rect 22327 25993 22336 26027
rect 22284 25984 22336 25993
rect 23112 25984 23164 26036
rect 29920 26027 29972 26036
rect 29920 25993 29929 26027
rect 29929 25993 29963 26027
rect 29963 25993 29972 26027
rect 29920 25984 29972 25993
rect 19432 25916 19484 25968
rect 29184 25916 29236 25968
rect 4344 25891 4396 25900
rect 4344 25857 4353 25891
rect 4353 25857 4387 25891
rect 4387 25857 4396 25891
rect 4344 25848 4396 25857
rect 9496 25848 9548 25900
rect 11704 25848 11756 25900
rect 14556 25848 14608 25900
rect 18420 25891 18472 25900
rect 18420 25857 18429 25891
rect 18429 25857 18463 25891
rect 18463 25857 18472 25891
rect 18420 25848 18472 25857
rect 22008 25848 22060 25900
rect 24676 25848 24728 25900
rect 24860 25891 24912 25900
rect 24860 25857 24894 25891
rect 24894 25857 24912 25891
rect 24860 25848 24912 25857
rect 6552 25823 6604 25832
rect 6552 25789 6561 25823
rect 6561 25789 6595 25823
rect 6595 25789 6604 25823
rect 6552 25780 6604 25789
rect 11980 25780 12032 25832
rect 12992 25823 13044 25832
rect 12992 25789 13001 25823
rect 13001 25789 13035 25823
rect 13035 25789 13044 25823
rect 12992 25780 13044 25789
rect 20444 25823 20496 25832
rect 20444 25789 20453 25823
rect 20453 25789 20487 25823
rect 20487 25789 20496 25823
rect 20444 25780 20496 25789
rect 9128 25644 9180 25696
rect 15108 25712 15160 25764
rect 22652 25712 22704 25764
rect 24584 25823 24636 25832
rect 24584 25789 24593 25823
rect 24593 25789 24627 25823
rect 24627 25789 24636 25823
rect 24584 25780 24636 25789
rect 27988 25780 28040 25832
rect 29828 25780 29880 25832
rect 13176 25644 13228 25696
rect 25964 25687 26016 25696
rect 25964 25653 25973 25687
rect 25973 25653 26007 25687
rect 26007 25653 26016 25687
rect 25964 25644 26016 25653
rect 4664 25542 4716 25594
rect 4728 25542 4780 25594
rect 4792 25542 4844 25594
rect 4856 25542 4908 25594
rect 4920 25542 4972 25594
rect 12092 25542 12144 25594
rect 12156 25542 12208 25594
rect 12220 25542 12272 25594
rect 12284 25542 12336 25594
rect 12348 25542 12400 25594
rect 19520 25542 19572 25594
rect 19584 25542 19636 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 26948 25542 27000 25594
rect 27012 25542 27064 25594
rect 27076 25542 27128 25594
rect 27140 25542 27192 25594
rect 27204 25542 27256 25594
rect 4988 25440 5040 25492
rect 8024 25440 8076 25492
rect 9496 25483 9548 25492
rect 9496 25449 9505 25483
rect 9505 25449 9539 25483
rect 9539 25449 9548 25483
rect 9496 25440 9548 25449
rect 24860 25440 24912 25492
rect 27988 25483 28040 25492
rect 27988 25449 27997 25483
rect 27997 25449 28031 25483
rect 28031 25449 28040 25483
rect 27988 25440 28040 25449
rect 3148 25279 3200 25288
rect 3148 25245 3157 25279
rect 3157 25245 3191 25279
rect 3191 25245 3200 25279
rect 3148 25236 3200 25245
rect 3240 25279 3292 25288
rect 3240 25245 3249 25279
rect 3249 25245 3283 25279
rect 3283 25245 3292 25279
rect 3240 25236 3292 25245
rect 4068 25236 4120 25288
rect 4160 25279 4212 25288
rect 4160 25245 4169 25279
rect 4169 25245 4203 25279
rect 4203 25245 4212 25279
rect 4160 25236 4212 25245
rect 6828 25236 6880 25288
rect 11152 25372 11204 25424
rect 26332 25372 26384 25424
rect 11796 25304 11848 25356
rect 11980 25304 12032 25356
rect 19524 25347 19576 25356
rect 19524 25313 19533 25347
rect 19533 25313 19567 25347
rect 19567 25313 19576 25347
rect 19524 25304 19576 25313
rect 22652 25304 22704 25356
rect 25412 25304 25464 25356
rect 25964 25304 26016 25356
rect 26424 25304 26476 25356
rect 31024 25304 31076 25356
rect 10232 25236 10284 25288
rect 18788 25236 18840 25288
rect 22744 25279 22796 25288
rect 22744 25245 22753 25279
rect 22753 25245 22787 25279
rect 22787 25245 22796 25279
rect 22744 25236 22796 25245
rect 22928 25279 22980 25288
rect 22928 25245 22937 25279
rect 22937 25245 22971 25279
rect 22971 25245 22980 25279
rect 22928 25236 22980 25245
rect 26608 25236 26660 25288
rect 27804 25236 27856 25288
rect 28908 25236 28960 25288
rect 29828 25279 29880 25288
rect 29828 25245 29837 25279
rect 29837 25245 29871 25279
rect 29871 25245 29880 25279
rect 29828 25236 29880 25245
rect 5264 25168 5316 25220
rect 7012 25211 7064 25220
rect 7012 25177 7046 25211
rect 7046 25177 7064 25211
rect 7012 25168 7064 25177
rect 10784 25211 10836 25220
rect 10784 25177 10793 25211
rect 10793 25177 10827 25211
rect 10827 25177 10836 25211
rect 10784 25168 10836 25177
rect 14556 25168 14608 25220
rect 2872 25100 2924 25152
rect 9864 25143 9916 25152
rect 9864 25109 9873 25143
rect 9873 25109 9907 25143
rect 9907 25109 9916 25143
rect 9864 25100 9916 25109
rect 23664 25100 23716 25152
rect 25044 25100 25096 25152
rect 28448 25100 28500 25152
rect 8378 24998 8430 25050
rect 8442 24998 8494 25050
rect 8506 24998 8558 25050
rect 8570 24998 8622 25050
rect 8634 24998 8686 25050
rect 15806 24998 15858 25050
rect 15870 24998 15922 25050
rect 15934 24998 15986 25050
rect 15998 24998 16050 25050
rect 16062 24998 16114 25050
rect 23234 24998 23286 25050
rect 23298 24998 23350 25050
rect 23362 24998 23414 25050
rect 23426 24998 23478 25050
rect 23490 24998 23542 25050
rect 30662 24998 30714 25050
rect 30726 24998 30778 25050
rect 30790 24998 30842 25050
rect 30854 24998 30906 25050
rect 30918 24998 30970 25050
rect 6552 24896 6604 24948
rect 7012 24896 7064 24948
rect 8024 24896 8076 24948
rect 11152 24896 11204 24948
rect 11704 24896 11756 24948
rect 18236 24896 18288 24948
rect 22192 24896 22244 24948
rect 15660 24828 15712 24880
rect 28448 24871 28500 24880
rect 28448 24837 28457 24871
rect 28457 24837 28491 24871
rect 28491 24837 28500 24871
rect 28448 24828 28500 24837
rect 2964 24760 3016 24812
rect 3056 24803 3108 24812
rect 3056 24769 3065 24803
rect 3065 24769 3099 24803
rect 3099 24769 3108 24803
rect 3056 24760 3108 24769
rect 3516 24803 3568 24812
rect 3516 24769 3525 24803
rect 3525 24769 3559 24803
rect 3559 24769 3568 24803
rect 3516 24760 3568 24769
rect 6736 24760 6788 24812
rect 8760 24760 8812 24812
rect 9956 24692 10008 24744
rect 14004 24760 14056 24812
rect 14096 24803 14148 24812
rect 14096 24769 14105 24803
rect 14105 24769 14139 24803
rect 14139 24769 14148 24803
rect 14096 24760 14148 24769
rect 14648 24760 14700 24812
rect 15936 24803 15988 24812
rect 13360 24692 13412 24744
rect 15936 24769 15945 24803
rect 15945 24769 15979 24803
rect 15979 24769 15988 24803
rect 15936 24760 15988 24769
rect 17868 24760 17920 24812
rect 20444 24760 20496 24812
rect 15016 24735 15068 24744
rect 15016 24701 15025 24735
rect 15025 24701 15059 24735
rect 15059 24701 15068 24735
rect 15016 24692 15068 24701
rect 15108 24692 15160 24744
rect 16304 24692 16356 24744
rect 16580 24692 16632 24744
rect 11336 24624 11388 24676
rect 3424 24556 3476 24608
rect 4344 24556 4396 24608
rect 8116 24599 8168 24608
rect 8116 24565 8125 24599
rect 8125 24565 8159 24599
rect 8159 24565 8168 24599
rect 8116 24556 8168 24565
rect 11612 24556 11664 24608
rect 19892 24735 19944 24744
rect 19892 24701 19901 24735
rect 19901 24701 19935 24735
rect 19935 24701 19944 24735
rect 19892 24692 19944 24701
rect 19340 24624 19392 24676
rect 19524 24624 19576 24676
rect 22192 24760 22244 24812
rect 27804 24760 27856 24812
rect 29552 24760 29604 24812
rect 21364 24692 21416 24744
rect 21824 24692 21876 24744
rect 24584 24692 24636 24744
rect 25780 24735 25832 24744
rect 25780 24701 25789 24735
rect 25789 24701 25823 24735
rect 25823 24701 25832 24735
rect 25780 24692 25832 24701
rect 26056 24735 26108 24744
rect 26056 24701 26065 24735
rect 26065 24701 26099 24735
rect 26099 24701 26108 24735
rect 26056 24692 26108 24701
rect 18512 24556 18564 24608
rect 20352 24599 20404 24608
rect 20352 24565 20361 24599
rect 20361 24565 20395 24599
rect 20395 24565 20404 24599
rect 20352 24556 20404 24565
rect 23112 24556 23164 24608
rect 28908 24692 28960 24744
rect 28264 24556 28316 24608
rect 4664 24454 4716 24506
rect 4728 24454 4780 24506
rect 4792 24454 4844 24506
rect 4856 24454 4908 24506
rect 4920 24454 4972 24506
rect 12092 24454 12144 24506
rect 12156 24454 12208 24506
rect 12220 24454 12272 24506
rect 12284 24454 12336 24506
rect 12348 24454 12400 24506
rect 19520 24454 19572 24506
rect 19584 24454 19636 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 26948 24454 27000 24506
rect 27012 24454 27064 24506
rect 27076 24454 27128 24506
rect 27140 24454 27192 24506
rect 27204 24454 27256 24506
rect 2964 24395 3016 24404
rect 2964 24361 2973 24395
rect 2973 24361 3007 24395
rect 3007 24361 3016 24395
rect 2964 24352 3016 24361
rect 3240 24352 3292 24404
rect 3976 24352 4028 24404
rect 15936 24352 15988 24404
rect 17868 24395 17920 24404
rect 17868 24361 17877 24395
rect 17877 24361 17911 24395
rect 17911 24361 17920 24395
rect 17868 24352 17920 24361
rect 22744 24395 22796 24404
rect 22744 24361 22753 24395
rect 22753 24361 22787 24395
rect 22787 24361 22796 24395
rect 22744 24352 22796 24361
rect 3148 24284 3200 24336
rect 2320 24191 2372 24200
rect 2320 24157 2329 24191
rect 2329 24157 2363 24191
rect 2363 24157 2372 24191
rect 2320 24148 2372 24157
rect 3424 24259 3476 24268
rect 3424 24225 3433 24259
rect 3433 24225 3467 24259
rect 3467 24225 3476 24259
rect 3424 24216 3476 24225
rect 5172 24284 5224 24336
rect 7380 24259 7432 24268
rect 7380 24225 7389 24259
rect 7389 24225 7423 24259
rect 7423 24225 7432 24259
rect 7380 24216 7432 24225
rect 11336 24259 11388 24268
rect 11336 24225 11345 24259
rect 11345 24225 11379 24259
rect 11379 24225 11388 24259
rect 11336 24216 11388 24225
rect 11612 24259 11664 24268
rect 11612 24225 11621 24259
rect 11621 24225 11655 24259
rect 11655 24225 11664 24259
rect 11612 24216 11664 24225
rect 13360 24259 13412 24268
rect 13360 24225 13369 24259
rect 13369 24225 13403 24259
rect 13403 24225 13412 24259
rect 13360 24216 13412 24225
rect 18420 24259 18472 24268
rect 18420 24225 18429 24259
rect 18429 24225 18463 24259
rect 18463 24225 18472 24259
rect 18420 24216 18472 24225
rect 19892 24259 19944 24268
rect 19892 24225 19901 24259
rect 19901 24225 19935 24259
rect 19935 24225 19944 24259
rect 19892 24216 19944 24225
rect 19984 24259 20036 24268
rect 19984 24225 19993 24259
rect 19993 24225 20027 24259
rect 20027 24225 20036 24259
rect 19984 24216 20036 24225
rect 21364 24259 21416 24268
rect 21364 24225 21373 24259
rect 21373 24225 21407 24259
rect 21407 24225 21416 24259
rect 21364 24216 21416 24225
rect 25136 24259 25188 24268
rect 25136 24225 25145 24259
rect 25145 24225 25179 24259
rect 25179 24225 25188 24259
rect 25136 24216 25188 24225
rect 26148 24216 26200 24268
rect 27620 24216 27672 24268
rect 4160 24148 4212 24200
rect 6920 24148 6972 24200
rect 13452 24148 13504 24200
rect 18236 24191 18288 24200
rect 18236 24157 18245 24191
rect 18245 24157 18279 24191
rect 18279 24157 18288 24191
rect 18236 24148 18288 24157
rect 19340 24148 19392 24200
rect 22928 24148 22980 24200
rect 24952 24148 25004 24200
rect 26332 24191 26384 24200
rect 26332 24157 26341 24191
rect 26341 24157 26375 24191
rect 26375 24157 26384 24191
rect 26332 24148 26384 24157
rect 27896 24148 27948 24200
rect 28172 24191 28224 24200
rect 28172 24157 28181 24191
rect 28181 24157 28215 24191
rect 28215 24157 28224 24191
rect 28172 24148 28224 24157
rect 29552 24216 29604 24268
rect 28448 24148 28500 24200
rect 4160 24055 4212 24064
rect 4160 24021 4185 24055
rect 4185 24021 4212 24055
rect 12624 24080 12676 24132
rect 14096 24080 14148 24132
rect 15016 24080 15068 24132
rect 22008 24080 22060 24132
rect 22744 24080 22796 24132
rect 24676 24080 24728 24132
rect 4160 24012 4212 24021
rect 7104 24012 7156 24064
rect 19432 24055 19484 24064
rect 19432 24021 19441 24055
rect 19441 24021 19475 24055
rect 19475 24021 19484 24055
rect 19432 24012 19484 24021
rect 20168 24012 20220 24064
rect 22376 24012 22428 24064
rect 23572 24055 23624 24064
rect 23572 24021 23581 24055
rect 23581 24021 23615 24055
rect 23615 24021 23624 24055
rect 23572 24012 23624 24021
rect 24860 24012 24912 24064
rect 28540 24080 28592 24132
rect 25780 24012 25832 24064
rect 26148 24055 26200 24064
rect 26148 24021 26157 24055
rect 26157 24021 26191 24055
rect 26191 24021 26200 24055
rect 26148 24012 26200 24021
rect 8378 23910 8430 23962
rect 8442 23910 8494 23962
rect 8506 23910 8558 23962
rect 8570 23910 8622 23962
rect 8634 23910 8686 23962
rect 15806 23910 15858 23962
rect 15870 23910 15922 23962
rect 15934 23910 15986 23962
rect 15998 23910 16050 23962
rect 16062 23910 16114 23962
rect 23234 23910 23286 23962
rect 23298 23910 23350 23962
rect 23362 23910 23414 23962
rect 23426 23910 23478 23962
rect 23490 23910 23542 23962
rect 30662 23910 30714 23962
rect 30726 23910 30778 23962
rect 30790 23910 30842 23962
rect 30854 23910 30906 23962
rect 30918 23910 30970 23962
rect 2320 23740 2372 23792
rect 2872 23783 2924 23792
rect 2872 23749 2906 23783
rect 2906 23749 2924 23783
rect 2872 23740 2924 23749
rect 3976 23851 4028 23860
rect 3976 23817 3985 23851
rect 3985 23817 4019 23851
rect 4019 23817 4028 23851
rect 3976 23808 4028 23817
rect 5264 23851 5316 23860
rect 5264 23817 5273 23851
rect 5273 23817 5307 23851
rect 5307 23817 5316 23851
rect 5264 23808 5316 23817
rect 13452 23851 13504 23860
rect 13452 23817 13461 23851
rect 13461 23817 13495 23851
rect 13495 23817 13504 23851
rect 13452 23808 13504 23817
rect 14096 23851 14148 23860
rect 14096 23817 14105 23851
rect 14105 23817 14139 23851
rect 14139 23817 14148 23851
rect 14096 23808 14148 23817
rect 16304 23851 16356 23860
rect 16304 23817 16313 23851
rect 16313 23817 16347 23851
rect 16347 23817 16356 23851
rect 16304 23808 16356 23817
rect 19892 23851 19944 23860
rect 19892 23817 19901 23851
rect 19901 23817 19935 23851
rect 19935 23817 19944 23851
rect 19892 23808 19944 23817
rect 22008 23851 22060 23860
rect 22008 23817 22017 23851
rect 22017 23817 22051 23851
rect 22051 23817 22060 23851
rect 22008 23808 22060 23817
rect 22744 23808 22796 23860
rect 26332 23808 26384 23860
rect 28264 23808 28316 23860
rect 4068 23740 4120 23792
rect 2688 23672 2740 23724
rect 4988 23672 5040 23724
rect 6920 23740 6972 23792
rect 10784 23740 10836 23792
rect 11980 23740 12032 23792
rect 5172 23715 5224 23724
rect 5172 23681 5181 23715
rect 5181 23681 5215 23715
rect 5215 23681 5224 23715
rect 5172 23672 5224 23681
rect 5080 23604 5132 23656
rect 9680 23604 9732 23656
rect 10416 23715 10468 23724
rect 10416 23681 10425 23715
rect 10425 23681 10459 23715
rect 10459 23681 10468 23715
rect 10416 23672 10468 23681
rect 11060 23672 11112 23724
rect 12624 23740 12676 23792
rect 14648 23740 14700 23792
rect 19432 23740 19484 23792
rect 23112 23740 23164 23792
rect 28172 23740 28224 23792
rect 11244 23604 11296 23656
rect 12992 23604 13044 23656
rect 13728 23672 13780 23724
rect 14004 23715 14056 23724
rect 14004 23681 14013 23715
rect 14013 23681 14047 23715
rect 14047 23681 14056 23715
rect 14004 23672 14056 23681
rect 15476 23672 15528 23724
rect 18512 23715 18564 23724
rect 18512 23681 18521 23715
rect 18521 23681 18555 23715
rect 18555 23681 18564 23715
rect 18512 23672 18564 23681
rect 20720 23672 20772 23724
rect 22376 23715 22428 23724
rect 22376 23681 22385 23715
rect 22385 23681 22419 23715
rect 22419 23681 22428 23715
rect 22376 23672 22428 23681
rect 25688 23672 25740 23724
rect 25964 23672 26016 23724
rect 26516 23715 26568 23724
rect 26516 23681 26525 23715
rect 26525 23681 26559 23715
rect 26559 23681 26568 23715
rect 26516 23672 26568 23681
rect 28908 23672 28960 23724
rect 14924 23647 14976 23656
rect 14924 23613 14933 23647
rect 14933 23613 14967 23647
rect 14967 23613 14976 23647
rect 14924 23604 14976 23613
rect 20904 23647 20956 23656
rect 20904 23613 20913 23647
rect 20913 23613 20947 23647
rect 20947 23613 20956 23647
rect 20904 23604 20956 23613
rect 22652 23647 22704 23656
rect 22652 23613 22661 23647
rect 22661 23613 22695 23647
rect 22695 23613 22704 23647
rect 22652 23604 22704 23613
rect 26424 23647 26476 23656
rect 26424 23613 26433 23647
rect 26433 23613 26467 23647
rect 26467 23613 26476 23647
rect 26424 23604 26476 23613
rect 20352 23536 20404 23588
rect 4528 23511 4580 23520
rect 4528 23477 4537 23511
rect 4537 23477 4571 23511
rect 4571 23477 4580 23511
rect 4528 23468 4580 23477
rect 10140 23511 10192 23520
rect 10140 23477 10149 23511
rect 10149 23477 10183 23511
rect 10183 23477 10192 23511
rect 10140 23468 10192 23477
rect 11520 23468 11572 23520
rect 18420 23468 18472 23520
rect 19984 23468 20036 23520
rect 23020 23468 23072 23520
rect 4664 23366 4716 23418
rect 4728 23366 4780 23418
rect 4792 23366 4844 23418
rect 4856 23366 4908 23418
rect 4920 23366 4972 23418
rect 12092 23366 12144 23418
rect 12156 23366 12208 23418
rect 12220 23366 12272 23418
rect 12284 23366 12336 23418
rect 12348 23366 12400 23418
rect 19520 23366 19572 23418
rect 19584 23366 19636 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 26948 23366 27000 23418
rect 27012 23366 27064 23418
rect 27076 23366 27128 23418
rect 27140 23366 27192 23418
rect 27204 23366 27256 23418
rect 4252 23307 4304 23316
rect 4252 23273 4261 23307
rect 4261 23273 4295 23307
rect 4295 23273 4304 23307
rect 4252 23264 4304 23273
rect 4988 23307 5040 23316
rect 4988 23273 4997 23307
rect 4997 23273 5031 23307
rect 5031 23273 5040 23307
rect 4988 23264 5040 23273
rect 6736 23264 6788 23316
rect 5172 23196 5224 23248
rect 2320 23128 2372 23180
rect 1860 23103 1912 23112
rect 1860 23069 1869 23103
rect 1869 23069 1903 23103
rect 1903 23069 1912 23103
rect 1860 23060 1912 23069
rect 3700 23060 3752 23112
rect 4528 23060 4580 23112
rect 2320 22924 2372 22976
rect 4160 22924 4212 22976
rect 5816 23103 5868 23112
rect 5816 23069 5825 23103
rect 5825 23069 5859 23103
rect 5859 23069 5868 23103
rect 5816 23060 5868 23069
rect 10140 23264 10192 23316
rect 11980 23264 12032 23316
rect 15476 23307 15528 23316
rect 15476 23273 15485 23307
rect 15485 23273 15519 23307
rect 15519 23273 15528 23307
rect 15476 23264 15528 23273
rect 21088 23307 21140 23316
rect 21088 23273 21097 23307
rect 21097 23273 21131 23307
rect 21131 23273 21140 23307
rect 21088 23264 21140 23273
rect 24952 23264 25004 23316
rect 25780 23264 25832 23316
rect 26516 23264 26568 23316
rect 11244 23196 11296 23248
rect 23112 23196 23164 23248
rect 23572 23196 23624 23248
rect 8760 23128 8812 23180
rect 15660 23128 15712 23180
rect 16580 23128 16632 23180
rect 19984 23171 20036 23180
rect 19984 23137 19993 23171
rect 19993 23137 20027 23171
rect 20027 23137 20036 23171
rect 19984 23128 20036 23137
rect 10784 23060 10836 23112
rect 13360 23060 13412 23112
rect 16304 23060 16356 23112
rect 20904 23060 20956 23112
rect 23020 23103 23072 23112
rect 23020 23069 23029 23103
rect 23029 23069 23063 23103
rect 23063 23069 23072 23103
rect 23020 23060 23072 23069
rect 23112 23103 23164 23112
rect 23112 23069 23122 23103
rect 23122 23069 23156 23103
rect 23156 23069 23164 23103
rect 23112 23060 23164 23069
rect 24584 23171 24636 23180
rect 24584 23137 24593 23171
rect 24593 23137 24627 23171
rect 24627 23137 24636 23171
rect 24584 23128 24636 23137
rect 25872 23128 25924 23180
rect 23664 23060 23716 23112
rect 24860 23103 24912 23112
rect 24860 23069 24894 23103
rect 24894 23069 24912 23103
rect 24860 23060 24912 23069
rect 6092 23035 6144 23044
rect 6092 23001 6101 23035
rect 6101 23001 6135 23035
rect 6135 23001 6144 23035
rect 6092 22992 6144 23001
rect 7104 22992 7156 23044
rect 21456 22992 21508 23044
rect 28540 23103 28592 23112
rect 28540 23069 28549 23103
rect 28549 23069 28583 23103
rect 28583 23069 28592 23103
rect 28540 23060 28592 23069
rect 28908 23060 28960 23112
rect 14740 22924 14792 22976
rect 15476 22924 15528 22976
rect 19432 22967 19484 22976
rect 19432 22933 19441 22967
rect 19441 22933 19475 22967
rect 19475 22933 19484 22967
rect 19432 22924 19484 22933
rect 20076 22924 20128 22976
rect 21272 22924 21324 22976
rect 22376 22924 22428 22976
rect 25044 22924 25096 22976
rect 28356 22924 28408 22976
rect 28632 22924 28684 22976
rect 8378 22822 8430 22874
rect 8442 22822 8494 22874
rect 8506 22822 8558 22874
rect 8570 22822 8622 22874
rect 8634 22822 8686 22874
rect 15806 22822 15858 22874
rect 15870 22822 15922 22874
rect 15934 22822 15986 22874
rect 15998 22822 16050 22874
rect 16062 22822 16114 22874
rect 23234 22822 23286 22874
rect 23298 22822 23350 22874
rect 23362 22822 23414 22874
rect 23426 22822 23478 22874
rect 23490 22822 23542 22874
rect 30662 22822 30714 22874
rect 30726 22822 30778 22874
rect 30790 22822 30842 22874
rect 30854 22822 30906 22874
rect 30918 22822 30970 22874
rect 4068 22720 4120 22772
rect 6092 22720 6144 22772
rect 8760 22763 8812 22772
rect 8760 22729 8769 22763
rect 8769 22729 8803 22763
rect 8803 22729 8812 22763
rect 8760 22720 8812 22729
rect 15660 22720 15712 22772
rect 1860 22652 1912 22704
rect 3332 22652 3384 22704
rect 8116 22652 8168 22704
rect 2228 22627 2280 22636
rect 2228 22593 2237 22627
rect 2237 22593 2271 22627
rect 2271 22593 2280 22627
rect 2228 22584 2280 22593
rect 2964 22627 3016 22636
rect 2964 22593 2998 22627
rect 2998 22593 3016 22627
rect 2964 22584 3016 22593
rect 4252 22584 4304 22636
rect 2688 22559 2740 22568
rect 2688 22525 2697 22559
rect 2697 22525 2731 22559
rect 2731 22525 2740 22559
rect 2688 22516 2740 22525
rect 4988 22516 5040 22568
rect 5172 22584 5224 22636
rect 6736 22627 6788 22636
rect 6736 22593 6745 22627
rect 6745 22593 6779 22627
rect 6779 22593 6788 22627
rect 6736 22584 6788 22593
rect 6828 22584 6880 22636
rect 9772 22652 9824 22704
rect 11520 22652 11572 22704
rect 14740 22695 14792 22704
rect 14740 22661 14749 22695
rect 14749 22661 14783 22695
rect 14783 22661 14792 22695
rect 14740 22652 14792 22661
rect 20168 22720 20220 22772
rect 20904 22720 20956 22772
rect 21456 22763 21508 22772
rect 21456 22729 21465 22763
rect 21465 22729 21499 22763
rect 21499 22729 21508 22763
rect 21456 22720 21508 22729
rect 22376 22763 22428 22772
rect 22376 22729 22385 22763
rect 22385 22729 22419 22763
rect 22419 22729 22428 22763
rect 22376 22720 22428 22729
rect 23112 22720 23164 22772
rect 25872 22763 25924 22772
rect 25872 22729 25881 22763
rect 25881 22729 25915 22763
rect 25915 22729 25924 22763
rect 25872 22720 25924 22729
rect 28908 22720 28960 22772
rect 19432 22652 19484 22704
rect 22284 22652 22336 22704
rect 23020 22652 23072 22704
rect 28632 22695 28684 22704
rect 28632 22661 28641 22695
rect 28641 22661 28675 22695
rect 28675 22661 28684 22695
rect 28632 22652 28684 22661
rect 29184 22652 29236 22704
rect 8760 22584 8812 22636
rect 11428 22584 11480 22636
rect 12716 22584 12768 22636
rect 13176 22627 13228 22636
rect 13176 22593 13185 22627
rect 13185 22593 13219 22627
rect 13219 22593 13228 22627
rect 13176 22584 13228 22593
rect 5264 22516 5316 22568
rect 3700 22448 3752 22500
rect 9680 22516 9732 22568
rect 10416 22516 10468 22568
rect 11152 22516 11204 22568
rect 18512 22584 18564 22636
rect 23112 22584 23164 22636
rect 24584 22584 24636 22636
rect 24768 22627 24820 22636
rect 24768 22593 24802 22627
rect 24802 22593 24820 22627
rect 24768 22584 24820 22593
rect 28356 22627 28408 22636
rect 28356 22593 28365 22627
rect 28365 22593 28399 22627
rect 28399 22593 28408 22627
rect 28356 22584 28408 22593
rect 13084 22491 13136 22500
rect 13084 22457 13093 22491
rect 13093 22457 13127 22491
rect 13127 22457 13136 22491
rect 13084 22448 13136 22457
rect 22284 22516 22336 22568
rect 16580 22448 16632 22500
rect 17408 22448 17460 22500
rect 20352 22448 20404 22500
rect 3056 22380 3108 22432
rect 4160 22380 4212 22432
rect 4988 22380 5040 22432
rect 6828 22380 6880 22432
rect 12532 22380 12584 22432
rect 14740 22380 14792 22432
rect 15016 22423 15068 22432
rect 15016 22389 15025 22423
rect 15025 22389 15059 22423
rect 15059 22389 15068 22423
rect 15016 22380 15068 22389
rect 16672 22380 16724 22432
rect 22100 22380 22152 22432
rect 25136 22380 25188 22432
rect 4664 22278 4716 22330
rect 4728 22278 4780 22330
rect 4792 22278 4844 22330
rect 4856 22278 4908 22330
rect 4920 22278 4972 22330
rect 12092 22278 12144 22330
rect 12156 22278 12208 22330
rect 12220 22278 12272 22330
rect 12284 22278 12336 22330
rect 12348 22278 12400 22330
rect 19520 22278 19572 22330
rect 19584 22278 19636 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 26948 22278 27000 22330
rect 27012 22278 27064 22330
rect 27076 22278 27128 22330
rect 27140 22278 27192 22330
rect 27204 22278 27256 22330
rect 3700 22176 3752 22228
rect 5816 22176 5868 22228
rect 15660 22176 15712 22228
rect 24768 22219 24820 22228
rect 24768 22185 24777 22219
rect 24777 22185 24811 22219
rect 24811 22185 24820 22219
rect 24768 22176 24820 22185
rect 5264 22108 5316 22160
rect 9128 22108 9180 22160
rect 6828 22040 6880 22092
rect 10140 22083 10192 22092
rect 10140 22049 10149 22083
rect 10149 22049 10183 22083
rect 10183 22049 10192 22083
rect 10140 22040 10192 22049
rect 10416 22083 10468 22092
rect 10416 22049 10425 22083
rect 10425 22049 10459 22083
rect 10459 22049 10468 22083
rect 10416 22040 10468 22049
rect 11428 22083 11480 22092
rect 11428 22049 11437 22083
rect 11437 22049 11471 22083
rect 11471 22049 11480 22083
rect 11428 22040 11480 22049
rect 11796 22108 11848 22160
rect 15200 22108 15252 22160
rect 2688 21972 2740 22024
rect 4988 22015 5040 22024
rect 4988 21981 4997 22015
rect 4997 21981 5031 22015
rect 5031 21981 5040 22015
rect 4988 21972 5040 21981
rect 5724 22015 5776 22024
rect 5724 21981 5733 22015
rect 5733 21981 5767 22015
rect 5767 21981 5776 22015
rect 5724 21972 5776 21981
rect 6092 21972 6144 22024
rect 6460 21972 6512 22024
rect 10048 22015 10100 22024
rect 10048 21981 10057 22015
rect 10057 21981 10091 22015
rect 10091 21981 10100 22015
rect 10048 21972 10100 21981
rect 12992 22015 13044 22024
rect 12992 21981 13001 22015
rect 13001 21981 13035 22015
rect 13035 21981 13044 22015
rect 12992 21972 13044 21981
rect 14924 22040 14976 22092
rect 2320 21947 2372 21956
rect 2320 21913 2354 21947
rect 2354 21913 2372 21947
rect 2320 21904 2372 21913
rect 4160 21947 4212 21956
rect 4160 21913 4169 21947
rect 4169 21913 4203 21947
rect 4203 21913 4212 21947
rect 4160 21904 4212 21913
rect 7012 21947 7064 21956
rect 7012 21913 7021 21947
rect 7021 21913 7055 21947
rect 7055 21913 7064 21947
rect 7012 21904 7064 21913
rect 13176 21947 13228 21956
rect 13176 21913 13185 21947
rect 13185 21913 13219 21947
rect 13219 21913 13228 21947
rect 13176 21904 13228 21913
rect 15016 21947 15068 21956
rect 15016 21913 15025 21947
rect 15025 21913 15059 21947
rect 15059 21913 15068 21947
rect 15016 21904 15068 21913
rect 16672 22015 16724 22024
rect 16672 21981 16690 22015
rect 16690 21981 16724 22015
rect 16672 21972 16724 21981
rect 18512 22040 18564 22092
rect 20812 22040 20864 22092
rect 25136 22040 25188 22092
rect 25964 22083 26016 22092
rect 25964 22049 25973 22083
rect 25973 22049 26007 22083
rect 26007 22049 26016 22083
rect 25964 22040 26016 22049
rect 26240 22083 26292 22092
rect 26240 22049 26249 22083
rect 26249 22049 26283 22083
rect 26283 22049 26292 22083
rect 26240 22040 26292 22049
rect 29184 22083 29236 22092
rect 29184 22049 29193 22083
rect 29193 22049 29227 22083
rect 29227 22049 29236 22083
rect 29184 22040 29236 22049
rect 18144 21972 18196 22024
rect 21180 22015 21232 22024
rect 21180 21981 21189 22015
rect 21189 21981 21223 22015
rect 21223 21981 21232 22015
rect 21180 21972 21232 21981
rect 22836 21972 22888 22024
rect 25872 21972 25924 22024
rect 27620 21972 27672 22024
rect 28172 22015 28224 22024
rect 28172 21981 28181 22015
rect 28181 21981 28215 22015
rect 28215 21981 28224 22015
rect 28172 21972 28224 21981
rect 28448 22015 28500 22024
rect 28448 21981 28457 22015
rect 28457 21981 28491 22015
rect 28491 21981 28500 22015
rect 28448 21972 28500 21981
rect 29368 21972 29420 22024
rect 17224 21904 17276 21956
rect 10876 21836 10928 21888
rect 11152 21836 11204 21888
rect 12256 21879 12308 21888
rect 12256 21845 12265 21879
rect 12265 21845 12299 21879
rect 12299 21845 12308 21879
rect 12256 21836 12308 21845
rect 12440 21836 12492 21888
rect 23572 21904 23624 21956
rect 25688 21904 25740 21956
rect 31024 21904 31076 21956
rect 27896 21836 27948 21888
rect 8378 21734 8430 21786
rect 8442 21734 8494 21786
rect 8506 21734 8558 21786
rect 8570 21734 8622 21786
rect 8634 21734 8686 21786
rect 15806 21734 15858 21786
rect 15870 21734 15922 21786
rect 15934 21734 15986 21786
rect 15998 21734 16050 21786
rect 16062 21734 16114 21786
rect 23234 21734 23286 21786
rect 23298 21734 23350 21786
rect 23362 21734 23414 21786
rect 23426 21734 23478 21786
rect 23490 21734 23542 21786
rect 30662 21734 30714 21786
rect 30726 21734 30778 21786
rect 30790 21734 30842 21786
rect 30854 21734 30906 21786
rect 30918 21734 30970 21786
rect 9680 21632 9732 21684
rect 13084 21632 13136 21684
rect 4344 21607 4396 21616
rect 4344 21573 4353 21607
rect 4353 21573 4387 21607
rect 4387 21573 4396 21607
rect 4344 21564 4396 21573
rect 5724 21564 5776 21616
rect 8760 21564 8812 21616
rect 8024 21496 8076 21548
rect 11060 21564 11112 21616
rect 12440 21607 12492 21616
rect 12440 21573 12449 21607
rect 12449 21573 12483 21607
rect 12483 21573 12492 21607
rect 12440 21564 12492 21573
rect 12532 21607 12584 21616
rect 12532 21573 12541 21607
rect 12541 21573 12575 21607
rect 12575 21573 12584 21607
rect 12532 21564 12584 21573
rect 23020 21632 23072 21684
rect 25228 21632 25280 21684
rect 27620 21632 27672 21684
rect 28540 21632 28592 21684
rect 18420 21607 18472 21616
rect 18420 21573 18429 21607
rect 18429 21573 18463 21607
rect 18463 21573 18472 21607
rect 18420 21564 18472 21573
rect 22100 21564 22152 21616
rect 26240 21564 26292 21616
rect 27896 21607 27948 21616
rect 27896 21573 27905 21607
rect 27905 21573 27939 21607
rect 27939 21573 27948 21607
rect 27896 21564 27948 21573
rect 9312 21539 9364 21548
rect 9312 21505 9346 21539
rect 9346 21505 9364 21539
rect 9312 21496 9364 21505
rect 10416 21496 10468 21548
rect 12256 21539 12308 21548
rect 12256 21505 12266 21539
rect 12266 21505 12300 21539
rect 12300 21505 12308 21539
rect 12256 21496 12308 21505
rect 12624 21539 12676 21548
rect 12624 21505 12638 21539
rect 12638 21505 12672 21539
rect 12672 21505 12676 21539
rect 12624 21496 12676 21505
rect 14924 21496 14976 21548
rect 17224 21539 17276 21548
rect 17224 21505 17233 21539
rect 17233 21505 17267 21539
rect 17267 21505 17276 21539
rect 17224 21496 17276 21505
rect 17960 21496 18012 21548
rect 18328 21539 18380 21548
rect 18328 21505 18337 21539
rect 18337 21505 18371 21539
rect 18371 21505 18380 21539
rect 18328 21496 18380 21505
rect 23572 21496 23624 21548
rect 24584 21496 24636 21548
rect 25504 21496 25556 21548
rect 29000 21496 29052 21548
rect 2688 21471 2740 21480
rect 2688 21437 2697 21471
rect 2697 21437 2731 21471
rect 2731 21437 2740 21471
rect 2688 21428 2740 21437
rect 6092 21428 6144 21480
rect 7380 21428 7432 21480
rect 9036 21471 9088 21480
rect 9036 21437 9045 21471
rect 9045 21437 9079 21471
rect 9079 21437 9088 21471
rect 9036 21428 9088 21437
rect 6276 21292 6328 21344
rect 13176 21292 13228 21344
rect 17408 21471 17460 21480
rect 17408 21437 17417 21471
rect 17417 21437 17451 21471
rect 17451 21437 17460 21471
rect 17408 21428 17460 21437
rect 25136 21428 25188 21480
rect 25320 21428 25372 21480
rect 27620 21471 27672 21480
rect 27620 21437 27629 21471
rect 27629 21437 27663 21471
rect 27663 21437 27672 21471
rect 27620 21428 27672 21437
rect 24860 21360 24912 21412
rect 26148 21360 26200 21412
rect 26700 21360 26752 21412
rect 20168 21292 20220 21344
rect 22652 21292 22704 21344
rect 24676 21335 24728 21344
rect 24676 21301 24685 21335
rect 24685 21301 24719 21335
rect 24719 21301 24728 21335
rect 24676 21292 24728 21301
rect 4664 21190 4716 21242
rect 4728 21190 4780 21242
rect 4792 21190 4844 21242
rect 4856 21190 4908 21242
rect 4920 21190 4972 21242
rect 12092 21190 12144 21242
rect 12156 21190 12208 21242
rect 12220 21190 12272 21242
rect 12284 21190 12336 21242
rect 12348 21190 12400 21242
rect 19520 21190 19572 21242
rect 19584 21190 19636 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 26948 21190 27000 21242
rect 27012 21190 27064 21242
rect 27076 21190 27128 21242
rect 27140 21190 27192 21242
rect 27204 21190 27256 21242
rect 2964 21131 3016 21140
rect 2964 21097 2973 21131
rect 2973 21097 3007 21131
rect 3007 21097 3016 21131
rect 2964 21088 3016 21097
rect 3332 21131 3384 21140
rect 3332 21097 3341 21131
rect 3341 21097 3375 21131
rect 3375 21097 3384 21131
rect 3332 21088 3384 21097
rect 2688 20952 2740 21004
rect 13820 21088 13872 21140
rect 14556 21131 14608 21140
rect 14556 21097 14565 21131
rect 14565 21097 14599 21131
rect 14599 21097 14608 21131
rect 14556 21088 14608 21097
rect 15200 21088 15252 21140
rect 18052 21088 18104 21140
rect 8760 21020 8812 21072
rect 9312 21020 9364 21072
rect 12624 21020 12676 21072
rect 22192 21088 22244 21140
rect 20168 21063 20220 21072
rect 20168 21029 20177 21063
rect 20177 21029 20211 21063
rect 20211 21029 20220 21063
rect 20168 21020 20220 21029
rect 3056 20884 3108 20936
rect 3976 20927 4028 20936
rect 3976 20893 3985 20927
rect 3985 20893 4019 20927
rect 4019 20893 4028 20927
rect 3976 20884 4028 20893
rect 6276 20995 6328 21004
rect 6276 20961 6285 20995
rect 6285 20961 6319 20995
rect 6319 20961 6328 20995
rect 6276 20952 6328 20961
rect 9680 20952 9732 21004
rect 9956 20995 10008 21004
rect 9956 20961 9965 20995
rect 9965 20961 9999 20995
rect 9999 20961 10008 20995
rect 9956 20952 10008 20961
rect 5540 20927 5592 20936
rect 5540 20893 5549 20927
rect 5549 20893 5583 20927
rect 5583 20893 5592 20927
rect 5540 20884 5592 20893
rect 10600 20927 10652 20936
rect 10600 20893 10609 20927
rect 10609 20893 10643 20927
rect 10643 20893 10652 20927
rect 10600 20884 10652 20893
rect 10876 20927 10928 20936
rect 10876 20893 10910 20927
rect 10910 20893 10928 20927
rect 10876 20884 10928 20893
rect 7012 20816 7064 20868
rect 11704 20816 11756 20868
rect 12716 20884 12768 20936
rect 14740 20927 14792 20936
rect 14740 20893 14749 20927
rect 14749 20893 14783 20927
rect 14783 20893 14792 20927
rect 14740 20884 14792 20893
rect 15292 20927 15344 20936
rect 15292 20893 15301 20927
rect 15301 20893 15335 20927
rect 15335 20893 15344 20927
rect 15292 20884 15344 20893
rect 4160 20748 4212 20800
rect 11428 20748 11480 20800
rect 16488 20816 16540 20868
rect 17500 20927 17552 20936
rect 17500 20893 17509 20927
rect 17509 20893 17543 20927
rect 17543 20893 17552 20927
rect 17500 20884 17552 20893
rect 14924 20748 14976 20800
rect 15200 20791 15252 20800
rect 15200 20757 15209 20791
rect 15209 20757 15243 20791
rect 15243 20757 15252 20791
rect 15200 20748 15252 20757
rect 17868 20816 17920 20868
rect 18788 20927 18840 20936
rect 18788 20893 18797 20927
rect 18797 20893 18831 20927
rect 18831 20893 18840 20927
rect 18788 20884 18840 20893
rect 19432 20884 19484 20936
rect 19984 20927 20036 20936
rect 19984 20893 19993 20927
rect 19993 20893 20027 20927
rect 20027 20893 20036 20927
rect 19984 20884 20036 20893
rect 20904 20927 20956 20936
rect 20904 20893 20913 20927
rect 20913 20893 20947 20927
rect 20947 20893 20956 20927
rect 20904 20884 20956 20893
rect 24860 21088 24912 21140
rect 26240 21088 26292 21140
rect 27620 21088 27672 21140
rect 24584 20927 24636 20936
rect 24584 20893 24593 20927
rect 24593 20893 24627 20927
rect 24627 20893 24636 20927
rect 24584 20884 24636 20893
rect 24676 20884 24728 20936
rect 21272 20816 21324 20868
rect 22192 20816 22244 20868
rect 29828 21020 29880 21072
rect 28172 20995 28224 21004
rect 28172 20961 28181 20995
rect 28181 20961 28215 20995
rect 28215 20961 28224 20995
rect 28172 20952 28224 20961
rect 29000 20995 29052 21004
rect 29000 20961 29009 20995
rect 29009 20961 29043 20995
rect 29043 20961 29052 20995
rect 29000 20952 29052 20961
rect 17960 20748 18012 20800
rect 22376 20748 22428 20800
rect 23112 20748 23164 20800
rect 28448 20927 28500 20936
rect 28448 20893 28457 20927
rect 28457 20893 28491 20927
rect 28491 20893 28500 20927
rect 28448 20884 28500 20893
rect 8378 20646 8430 20698
rect 8442 20646 8494 20698
rect 8506 20646 8558 20698
rect 8570 20646 8622 20698
rect 8634 20646 8686 20698
rect 15806 20646 15858 20698
rect 15870 20646 15922 20698
rect 15934 20646 15986 20698
rect 15998 20646 16050 20698
rect 16062 20646 16114 20698
rect 23234 20646 23286 20698
rect 23298 20646 23350 20698
rect 23362 20646 23414 20698
rect 23426 20646 23478 20698
rect 23490 20646 23542 20698
rect 30662 20646 30714 20698
rect 30726 20646 30778 20698
rect 30790 20646 30842 20698
rect 30854 20646 30906 20698
rect 30918 20646 30970 20698
rect 5540 20544 5592 20596
rect 4068 20476 4120 20528
rect 10048 20544 10100 20596
rect 10140 20544 10192 20596
rect 15292 20544 15344 20596
rect 15660 20544 15712 20596
rect 7104 20476 7156 20528
rect 2504 20383 2556 20392
rect 2504 20349 2513 20383
rect 2513 20349 2547 20383
rect 2547 20349 2556 20383
rect 2504 20340 2556 20349
rect 3976 20340 4028 20392
rect 6552 20383 6604 20392
rect 6552 20349 6561 20383
rect 6561 20349 6595 20383
rect 6595 20349 6604 20383
rect 6552 20340 6604 20349
rect 7196 20340 7248 20392
rect 9312 20451 9364 20460
rect 9312 20417 9346 20451
rect 9346 20417 9364 20451
rect 9312 20408 9364 20417
rect 9956 20476 10008 20528
rect 15200 20476 15252 20528
rect 14648 20451 14700 20460
rect 14648 20417 14657 20451
rect 14657 20417 14691 20451
rect 14691 20417 14700 20451
rect 14648 20408 14700 20417
rect 15568 20451 15620 20460
rect 15568 20417 15577 20451
rect 15577 20417 15611 20451
rect 15611 20417 15620 20451
rect 15568 20408 15620 20417
rect 16488 20408 16540 20460
rect 17408 20408 17460 20460
rect 18420 20519 18472 20528
rect 18420 20485 18429 20519
rect 18429 20485 18463 20519
rect 18463 20485 18472 20519
rect 18420 20476 18472 20485
rect 18788 20544 18840 20596
rect 20904 20544 20956 20596
rect 23572 20476 23624 20528
rect 19984 20408 20036 20460
rect 20812 20451 20864 20460
rect 20812 20417 20821 20451
rect 20821 20417 20855 20451
rect 20855 20417 20864 20451
rect 20812 20408 20864 20417
rect 21088 20451 21140 20460
rect 21088 20417 21097 20451
rect 21097 20417 21131 20451
rect 21131 20417 21140 20451
rect 21088 20408 21140 20417
rect 22376 20408 22428 20460
rect 24584 20408 24636 20460
rect 9772 20204 9824 20256
rect 10600 20204 10652 20256
rect 17500 20340 17552 20392
rect 17684 20340 17736 20392
rect 19892 20340 19944 20392
rect 21364 20383 21416 20392
rect 21364 20349 21373 20383
rect 21373 20349 21407 20383
rect 21407 20349 21416 20383
rect 21364 20340 21416 20349
rect 17776 20272 17828 20324
rect 15660 20204 15712 20256
rect 18328 20204 18380 20256
rect 22100 20247 22152 20256
rect 22100 20213 22109 20247
rect 22109 20213 22143 20247
rect 22143 20213 22152 20247
rect 22100 20204 22152 20213
rect 25320 20204 25372 20256
rect 4664 20102 4716 20154
rect 4728 20102 4780 20154
rect 4792 20102 4844 20154
rect 4856 20102 4908 20154
rect 4920 20102 4972 20154
rect 12092 20102 12144 20154
rect 12156 20102 12208 20154
rect 12220 20102 12272 20154
rect 12284 20102 12336 20154
rect 12348 20102 12400 20154
rect 19520 20102 19572 20154
rect 19584 20102 19636 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 26948 20102 27000 20154
rect 27012 20102 27064 20154
rect 27076 20102 27128 20154
rect 27140 20102 27192 20154
rect 27204 20102 27256 20154
rect 2504 20000 2556 20052
rect 4068 20043 4120 20052
rect 4068 20009 4077 20043
rect 4077 20009 4111 20043
rect 4111 20009 4120 20043
rect 4068 20000 4120 20009
rect 9312 20000 9364 20052
rect 18512 20000 18564 20052
rect 27988 20000 28040 20052
rect 9956 19932 10008 19984
rect 7104 19907 7156 19916
rect 7104 19873 7113 19907
rect 7113 19873 7147 19907
rect 7147 19873 7156 19907
rect 7104 19864 7156 19873
rect 22376 19932 22428 19984
rect 14740 19864 14792 19916
rect 18972 19864 19024 19916
rect 3884 19796 3936 19848
rect 4160 19839 4212 19848
rect 4160 19805 4169 19839
rect 4169 19805 4203 19839
rect 4203 19805 4212 19839
rect 4160 19796 4212 19805
rect 5264 19839 5316 19848
rect 5264 19805 5273 19839
rect 5273 19805 5307 19839
rect 5307 19805 5316 19839
rect 5264 19796 5316 19805
rect 6092 19839 6144 19848
rect 6092 19805 6101 19839
rect 6101 19805 6135 19839
rect 6135 19805 6144 19839
rect 6092 19796 6144 19805
rect 6460 19796 6512 19848
rect 9864 19839 9916 19848
rect 9864 19805 9873 19839
rect 9873 19805 9907 19839
rect 9907 19805 9916 19839
rect 9864 19796 9916 19805
rect 10140 19796 10192 19848
rect 18328 19796 18380 19848
rect 19432 19796 19484 19848
rect 20352 19864 20404 19916
rect 22100 19864 22152 19916
rect 25412 19864 25464 19916
rect 26700 19864 26752 19916
rect 17224 19728 17276 19780
rect 17592 19728 17644 19780
rect 18420 19728 18472 19780
rect 2136 19660 2188 19712
rect 6184 19660 6236 19712
rect 6552 19660 6604 19712
rect 10876 19660 10928 19712
rect 21364 19728 21416 19780
rect 22008 19728 22060 19780
rect 28448 19728 28500 19780
rect 24676 19703 24728 19712
rect 24676 19669 24685 19703
rect 24685 19669 24719 19703
rect 24719 19669 24728 19703
rect 24676 19660 24728 19669
rect 25872 19660 25924 19712
rect 28632 19703 28684 19712
rect 28632 19669 28641 19703
rect 28641 19669 28675 19703
rect 28675 19669 28684 19703
rect 28632 19660 28684 19669
rect 8378 19558 8430 19610
rect 8442 19558 8494 19610
rect 8506 19558 8558 19610
rect 8570 19558 8622 19610
rect 8634 19558 8686 19610
rect 15806 19558 15858 19610
rect 15870 19558 15922 19610
rect 15934 19558 15986 19610
rect 15998 19558 16050 19610
rect 16062 19558 16114 19610
rect 23234 19558 23286 19610
rect 23298 19558 23350 19610
rect 23362 19558 23414 19610
rect 23426 19558 23478 19610
rect 23490 19558 23542 19610
rect 30662 19558 30714 19610
rect 30726 19558 30778 19610
rect 30790 19558 30842 19610
rect 30854 19558 30906 19610
rect 30918 19558 30970 19610
rect 18420 19499 18472 19508
rect 18420 19465 18429 19499
rect 18429 19465 18463 19499
rect 18463 19465 18472 19499
rect 18420 19456 18472 19465
rect 2136 19431 2188 19440
rect 2136 19397 2145 19431
rect 2145 19397 2179 19431
rect 2179 19397 2188 19431
rect 2136 19388 2188 19397
rect 3884 19431 3936 19440
rect 3884 19397 3893 19431
rect 3893 19397 3927 19431
rect 3927 19397 3936 19431
rect 3884 19388 3936 19397
rect 3240 19320 3292 19372
rect 10600 19320 10652 19372
rect 12900 19363 12952 19372
rect 12900 19329 12909 19363
rect 12909 19329 12943 19363
rect 12943 19329 12952 19363
rect 12900 19320 12952 19329
rect 12992 19320 13044 19372
rect 1860 19295 1912 19304
rect 1860 19261 1869 19295
rect 1869 19261 1903 19295
rect 1903 19261 1912 19295
rect 1860 19252 1912 19261
rect 15200 19388 15252 19440
rect 15384 19388 15436 19440
rect 17592 19388 17644 19440
rect 22008 19388 22060 19440
rect 24676 19388 24728 19440
rect 25872 19499 25924 19508
rect 25872 19465 25881 19499
rect 25881 19465 25915 19499
rect 25915 19465 25924 19499
rect 25872 19456 25924 19465
rect 27436 19456 27488 19508
rect 28632 19456 28684 19508
rect 27988 19431 28040 19440
rect 27988 19397 27997 19431
rect 27997 19397 28031 19431
rect 28031 19397 28040 19431
rect 27988 19388 28040 19397
rect 15660 19320 15712 19372
rect 18512 19363 18564 19372
rect 18512 19329 18521 19363
rect 18521 19329 18555 19363
rect 18555 19329 18564 19363
rect 18512 19320 18564 19329
rect 23572 19320 23624 19372
rect 23664 19363 23716 19372
rect 23664 19329 23673 19363
rect 23673 19329 23707 19363
rect 23707 19329 23716 19363
rect 29920 19388 29972 19440
rect 23664 19320 23716 19329
rect 29000 19363 29052 19372
rect 29000 19329 29009 19363
rect 29009 19329 29043 19363
rect 29043 19329 29052 19363
rect 29000 19320 29052 19329
rect 29184 19363 29236 19372
rect 29184 19329 29193 19363
rect 29193 19329 29227 19363
rect 29227 19329 29236 19363
rect 29184 19320 29236 19329
rect 14464 19184 14516 19236
rect 15292 19184 15344 19236
rect 14280 19159 14332 19168
rect 14280 19125 14289 19159
rect 14289 19125 14323 19159
rect 14323 19125 14332 19159
rect 16212 19252 16264 19304
rect 29368 19295 29420 19304
rect 29368 19261 29377 19295
rect 29377 19261 29411 19295
rect 29411 19261 29420 19295
rect 29368 19252 29420 19261
rect 27712 19184 27764 19236
rect 14280 19116 14332 19125
rect 29184 19116 29236 19168
rect 4664 19014 4716 19066
rect 4728 19014 4780 19066
rect 4792 19014 4844 19066
rect 4856 19014 4908 19066
rect 4920 19014 4972 19066
rect 12092 19014 12144 19066
rect 12156 19014 12208 19066
rect 12220 19014 12272 19066
rect 12284 19014 12336 19066
rect 12348 19014 12400 19066
rect 19520 19014 19572 19066
rect 19584 19014 19636 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 26948 19014 27000 19066
rect 27012 19014 27064 19066
rect 27076 19014 27128 19066
rect 27140 19014 27192 19066
rect 27204 19014 27256 19066
rect 1860 18912 1912 18964
rect 3240 18912 3292 18964
rect 12992 18955 13044 18964
rect 12992 18921 13001 18955
rect 13001 18921 13035 18955
rect 13035 18921 13044 18955
rect 12992 18912 13044 18921
rect 25412 18912 25464 18964
rect 28448 18955 28500 18964
rect 28448 18921 28457 18955
rect 28457 18921 28491 18955
rect 28491 18921 28500 18955
rect 28448 18912 28500 18921
rect 29000 18912 29052 18964
rect 2504 18751 2556 18760
rect 2504 18717 2513 18751
rect 2513 18717 2547 18751
rect 2547 18717 2556 18751
rect 2504 18708 2556 18717
rect 3424 18751 3476 18760
rect 3424 18717 3433 18751
rect 3433 18717 3467 18751
rect 3467 18717 3476 18751
rect 3424 18708 3476 18717
rect 4068 18708 4120 18760
rect 12348 18776 12400 18828
rect 14372 18776 14424 18828
rect 17132 18776 17184 18828
rect 5724 18640 5776 18692
rect 9220 18708 9272 18760
rect 11152 18708 11204 18760
rect 13820 18708 13872 18760
rect 15292 18708 15344 18760
rect 16304 18708 16356 18760
rect 22928 18776 22980 18828
rect 23664 18776 23716 18828
rect 24584 18819 24636 18828
rect 24584 18785 24593 18819
rect 24593 18785 24627 18819
rect 24627 18785 24636 18819
rect 24584 18776 24636 18785
rect 18420 18708 18472 18760
rect 19432 18751 19484 18760
rect 19432 18717 19441 18751
rect 19441 18717 19475 18751
rect 19475 18717 19484 18751
rect 19432 18708 19484 18717
rect 19892 18751 19944 18760
rect 19892 18717 19901 18751
rect 19901 18717 19935 18751
rect 19935 18717 19944 18751
rect 19892 18708 19944 18717
rect 20996 18708 21048 18760
rect 27436 18751 27488 18760
rect 27436 18717 27445 18751
rect 27445 18717 27479 18751
rect 27479 18717 27488 18751
rect 27436 18708 27488 18717
rect 27988 18844 28040 18896
rect 28632 18708 28684 18760
rect 29828 18776 29880 18828
rect 29920 18776 29972 18828
rect 29184 18751 29236 18760
rect 29184 18717 29193 18751
rect 29193 18717 29227 18751
rect 29227 18717 29236 18751
rect 29184 18708 29236 18717
rect 14280 18640 14332 18692
rect 17408 18683 17460 18692
rect 17408 18649 17417 18683
rect 17417 18649 17451 18683
rect 17451 18649 17460 18683
rect 17408 18640 17460 18649
rect 17500 18683 17552 18692
rect 17500 18649 17509 18683
rect 17509 18649 17543 18683
rect 17543 18649 17552 18683
rect 17500 18640 17552 18649
rect 18052 18683 18104 18692
rect 18052 18649 18061 18683
rect 18061 18649 18095 18683
rect 18095 18649 18104 18683
rect 18052 18640 18104 18649
rect 24860 18683 24912 18692
rect 24860 18649 24869 18683
rect 24869 18649 24903 18683
rect 24903 18649 24912 18683
rect 24860 18640 24912 18649
rect 25320 18640 25372 18692
rect 27712 18683 27764 18692
rect 27712 18649 27721 18683
rect 27721 18649 27755 18683
rect 27755 18649 27764 18683
rect 27712 18640 27764 18649
rect 7472 18572 7524 18624
rect 8760 18572 8812 18624
rect 9128 18572 9180 18624
rect 15200 18572 15252 18624
rect 15476 18572 15528 18624
rect 16396 18615 16448 18624
rect 16396 18581 16405 18615
rect 16405 18581 16439 18615
rect 16439 18581 16448 18615
rect 16396 18572 16448 18581
rect 18328 18572 18380 18624
rect 20628 18615 20680 18624
rect 20628 18581 20637 18615
rect 20637 18581 20671 18615
rect 20671 18581 20680 18615
rect 20628 18572 20680 18581
rect 22468 18572 22520 18624
rect 26332 18615 26384 18624
rect 26332 18581 26341 18615
rect 26341 18581 26375 18615
rect 26375 18581 26384 18615
rect 26332 18572 26384 18581
rect 8378 18470 8430 18522
rect 8442 18470 8494 18522
rect 8506 18470 8558 18522
rect 8570 18470 8622 18522
rect 8634 18470 8686 18522
rect 15806 18470 15858 18522
rect 15870 18470 15922 18522
rect 15934 18470 15986 18522
rect 15998 18470 16050 18522
rect 16062 18470 16114 18522
rect 23234 18470 23286 18522
rect 23298 18470 23350 18522
rect 23362 18470 23414 18522
rect 23426 18470 23478 18522
rect 23490 18470 23542 18522
rect 30662 18470 30714 18522
rect 30726 18470 30778 18522
rect 30790 18470 30842 18522
rect 30854 18470 30906 18522
rect 30918 18470 30970 18522
rect 2504 18368 2556 18420
rect 2780 18300 2832 18352
rect 6552 18368 6604 18420
rect 7472 18343 7524 18352
rect 7472 18309 7481 18343
rect 7481 18309 7515 18343
rect 7515 18309 7524 18343
rect 7472 18300 7524 18309
rect 8760 18300 8812 18352
rect 9220 18343 9272 18352
rect 9220 18309 9229 18343
rect 9229 18309 9263 18343
rect 9263 18309 9272 18343
rect 9220 18300 9272 18309
rect 11704 18300 11756 18352
rect 15476 18368 15528 18420
rect 17132 18411 17184 18420
rect 17132 18377 17141 18411
rect 17141 18377 17175 18411
rect 17175 18377 17184 18411
rect 17132 18368 17184 18377
rect 5724 18232 5776 18284
rect 6736 18232 6788 18284
rect 10876 18232 10928 18284
rect 12900 18232 12952 18284
rect 14280 18232 14332 18284
rect 14740 18300 14792 18352
rect 15660 18300 15712 18352
rect 17408 18300 17460 18352
rect 15200 18232 15252 18284
rect 15292 18232 15344 18284
rect 2044 18207 2096 18216
rect 2044 18173 2053 18207
rect 2053 18173 2087 18207
rect 2087 18173 2096 18207
rect 2044 18164 2096 18173
rect 2320 18207 2372 18216
rect 2320 18173 2329 18207
rect 2329 18173 2363 18207
rect 2363 18173 2372 18207
rect 2320 18164 2372 18173
rect 12440 18207 12492 18216
rect 12440 18173 12449 18207
rect 12449 18173 12483 18207
rect 12483 18173 12492 18207
rect 12440 18164 12492 18173
rect 6000 18096 6052 18148
rect 11888 18096 11940 18148
rect 12348 18096 12400 18148
rect 15384 18164 15436 18216
rect 16212 18232 16264 18284
rect 16488 18164 16540 18216
rect 18052 18368 18104 18420
rect 22192 18368 22244 18420
rect 24860 18411 24912 18420
rect 24860 18377 24869 18411
rect 24869 18377 24903 18411
rect 24903 18377 24912 18411
rect 24860 18368 24912 18377
rect 26332 18368 26384 18420
rect 17684 18343 17736 18352
rect 17684 18309 17693 18343
rect 17693 18309 17727 18343
rect 17727 18309 17736 18343
rect 17684 18300 17736 18309
rect 18328 18300 18380 18352
rect 18972 18275 19024 18284
rect 18972 18241 18981 18275
rect 18981 18241 19015 18275
rect 19015 18241 19024 18275
rect 18972 18232 19024 18241
rect 20628 18300 20680 18352
rect 5816 18071 5868 18080
rect 5816 18037 5825 18071
rect 5825 18037 5859 18071
rect 5859 18037 5868 18071
rect 5816 18028 5868 18037
rect 9772 18071 9824 18080
rect 9772 18037 9781 18071
rect 9781 18037 9815 18071
rect 9815 18037 9824 18071
rect 9772 18028 9824 18037
rect 11980 18071 12032 18080
rect 11980 18037 11989 18071
rect 11989 18037 12023 18071
rect 12023 18037 12032 18071
rect 11980 18028 12032 18037
rect 16304 18028 16356 18080
rect 18236 18164 18288 18216
rect 21456 18164 21508 18216
rect 25228 18275 25280 18284
rect 25228 18241 25237 18275
rect 25237 18241 25271 18275
rect 25271 18241 25280 18275
rect 25228 18232 25280 18241
rect 29828 18275 29880 18284
rect 29828 18241 29837 18275
rect 29837 18241 29871 18275
rect 29871 18241 29880 18275
rect 29828 18232 29880 18241
rect 22928 18164 22980 18216
rect 25412 18207 25464 18216
rect 25412 18173 25421 18207
rect 25421 18173 25455 18207
rect 25455 18173 25464 18207
rect 25412 18164 25464 18173
rect 31024 18164 31076 18216
rect 20076 18028 20128 18080
rect 20996 18028 21048 18080
rect 22008 18071 22060 18080
rect 22008 18037 22017 18071
rect 22017 18037 22051 18071
rect 22051 18037 22060 18071
rect 22008 18028 22060 18037
rect 4664 17926 4716 17978
rect 4728 17926 4780 17978
rect 4792 17926 4844 17978
rect 4856 17926 4908 17978
rect 4920 17926 4972 17978
rect 12092 17926 12144 17978
rect 12156 17926 12208 17978
rect 12220 17926 12272 17978
rect 12284 17926 12336 17978
rect 12348 17926 12400 17978
rect 19520 17926 19572 17978
rect 19584 17926 19636 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 26948 17926 27000 17978
rect 27012 17926 27064 17978
rect 27076 17926 27128 17978
rect 27140 17926 27192 17978
rect 27204 17926 27256 17978
rect 2320 17824 2372 17876
rect 2780 17824 2832 17876
rect 11060 17824 11112 17876
rect 12440 17824 12492 17876
rect 10876 17799 10928 17808
rect 10876 17765 10885 17799
rect 10885 17765 10919 17799
rect 10919 17765 10928 17799
rect 10876 17756 10928 17765
rect 9128 17731 9180 17740
rect 9128 17697 9137 17731
rect 9137 17697 9171 17731
rect 9171 17697 9180 17731
rect 9128 17688 9180 17697
rect 9772 17688 9824 17740
rect 11980 17688 12032 17740
rect 2504 17620 2556 17672
rect 3332 17620 3384 17672
rect 3976 17620 4028 17672
rect 5080 17663 5132 17672
rect 5080 17629 5089 17663
rect 5089 17629 5123 17663
rect 5123 17629 5132 17663
rect 5080 17620 5132 17629
rect 5724 17663 5776 17672
rect 5724 17629 5733 17663
rect 5733 17629 5767 17663
rect 5767 17629 5776 17663
rect 5724 17620 5776 17629
rect 6552 17620 6604 17672
rect 12440 17620 12492 17672
rect 12900 17620 12952 17672
rect 14280 17867 14332 17876
rect 14280 17833 14289 17867
rect 14289 17833 14323 17867
rect 14323 17833 14332 17867
rect 14280 17824 14332 17833
rect 21456 17867 21508 17876
rect 21456 17833 21465 17867
rect 21465 17833 21499 17867
rect 21499 17833 21508 17867
rect 21456 17824 21508 17833
rect 14372 17756 14424 17808
rect 14740 17731 14792 17740
rect 14740 17697 14749 17731
rect 14749 17697 14783 17731
rect 14783 17697 14792 17731
rect 14740 17688 14792 17697
rect 16304 17688 16356 17740
rect 15200 17620 15252 17672
rect 15660 17663 15712 17672
rect 15660 17629 15669 17663
rect 15669 17629 15703 17663
rect 15703 17629 15712 17663
rect 15660 17620 15712 17629
rect 16396 17620 16448 17672
rect 6736 17552 6788 17604
rect 7472 17552 7524 17604
rect 3332 17527 3384 17536
rect 3332 17493 3341 17527
rect 3341 17493 3375 17527
rect 3375 17493 3384 17527
rect 3332 17484 3384 17493
rect 6828 17484 6880 17536
rect 10968 17552 11020 17604
rect 15108 17552 15160 17604
rect 15476 17552 15528 17604
rect 18420 17663 18472 17672
rect 18420 17629 18429 17663
rect 18429 17629 18463 17663
rect 18463 17629 18472 17663
rect 18420 17620 18472 17629
rect 20076 17731 20128 17740
rect 20076 17697 20085 17731
rect 20085 17697 20119 17731
rect 20119 17697 20128 17731
rect 20076 17688 20128 17697
rect 17868 17552 17920 17604
rect 17960 17484 18012 17536
rect 18144 17552 18196 17604
rect 22008 17620 22060 17672
rect 22468 17595 22520 17604
rect 22468 17561 22502 17595
rect 22502 17561 22520 17595
rect 22468 17552 22520 17561
rect 22744 17620 22796 17672
rect 25228 17620 25280 17672
rect 27620 17620 27672 17672
rect 23664 17552 23716 17604
rect 23572 17527 23624 17536
rect 23572 17493 23581 17527
rect 23581 17493 23615 17527
rect 23615 17493 23624 17527
rect 23572 17484 23624 17493
rect 26424 17484 26476 17536
rect 8378 17382 8430 17434
rect 8442 17382 8494 17434
rect 8506 17382 8558 17434
rect 8570 17382 8622 17434
rect 8634 17382 8686 17434
rect 15806 17382 15858 17434
rect 15870 17382 15922 17434
rect 15934 17382 15986 17434
rect 15998 17382 16050 17434
rect 16062 17382 16114 17434
rect 23234 17382 23286 17434
rect 23298 17382 23350 17434
rect 23362 17382 23414 17434
rect 23426 17382 23478 17434
rect 23490 17382 23542 17434
rect 30662 17382 30714 17434
rect 30726 17382 30778 17434
rect 30790 17382 30842 17434
rect 30854 17382 30906 17434
rect 30918 17382 30970 17434
rect 5724 17280 5776 17332
rect 3976 17255 4028 17264
rect 3976 17221 3985 17255
rect 3985 17221 4019 17255
rect 4019 17221 4028 17255
rect 3976 17212 4028 17221
rect 5816 17212 5868 17264
rect 6828 17323 6880 17332
rect 6828 17289 6837 17323
rect 6837 17289 6871 17323
rect 6871 17289 6880 17323
rect 6828 17280 6880 17289
rect 7472 17323 7524 17332
rect 7472 17289 7481 17323
rect 7481 17289 7515 17323
rect 7515 17289 7524 17323
rect 7472 17280 7524 17289
rect 2872 17187 2924 17196
rect 2872 17153 2881 17187
rect 2881 17153 2915 17187
rect 2915 17153 2924 17187
rect 2872 17144 2924 17153
rect 3424 17144 3476 17196
rect 6000 17187 6052 17196
rect 6000 17153 6009 17187
rect 6009 17153 6043 17187
rect 6043 17153 6052 17187
rect 6000 17144 6052 17153
rect 6736 17187 6788 17196
rect 6736 17153 6745 17187
rect 6745 17153 6779 17187
rect 6779 17153 6788 17187
rect 6736 17144 6788 17153
rect 12440 17212 12492 17264
rect 13820 17280 13872 17332
rect 14648 17280 14700 17332
rect 16764 17280 16816 17332
rect 17776 17280 17828 17332
rect 14004 17255 14056 17264
rect 14004 17221 14013 17255
rect 14013 17221 14047 17255
rect 14047 17221 14056 17255
rect 14004 17212 14056 17221
rect 15292 17212 15344 17264
rect 15384 17212 15436 17264
rect 11796 17144 11848 17196
rect 5724 17119 5776 17128
rect 5724 17085 5733 17119
rect 5733 17085 5767 17119
rect 5767 17085 5776 17119
rect 5724 17076 5776 17085
rect 13084 17051 13136 17060
rect 13084 17017 13093 17051
rect 13093 17017 13127 17051
rect 13127 17017 13136 17051
rect 15200 17187 15252 17196
rect 15200 17153 15209 17187
rect 15209 17153 15243 17187
rect 15243 17153 15252 17187
rect 15200 17144 15252 17153
rect 15476 17187 15528 17196
rect 15476 17153 15485 17187
rect 15485 17153 15519 17187
rect 15519 17153 15528 17187
rect 15476 17144 15528 17153
rect 16212 17212 16264 17264
rect 18144 17212 18196 17264
rect 16120 17144 16172 17196
rect 16764 17144 16816 17196
rect 17500 17187 17552 17196
rect 17500 17153 17509 17187
rect 17509 17153 17543 17187
rect 17543 17153 17552 17187
rect 17500 17144 17552 17153
rect 18236 17187 18288 17196
rect 18236 17153 18245 17187
rect 18245 17153 18279 17187
rect 18279 17153 18288 17187
rect 18236 17144 18288 17153
rect 18328 17187 18380 17196
rect 18328 17153 18337 17187
rect 18337 17153 18371 17187
rect 18371 17153 18380 17187
rect 18328 17144 18380 17153
rect 19432 17280 19484 17332
rect 22468 17280 22520 17332
rect 27620 17280 27672 17332
rect 27436 17255 27488 17264
rect 27436 17221 27445 17255
rect 27445 17221 27479 17255
rect 27479 17221 27488 17255
rect 27436 17212 27488 17221
rect 14280 17076 14332 17128
rect 15752 17119 15804 17128
rect 15752 17085 15761 17119
rect 15761 17085 15795 17119
rect 15795 17085 15804 17119
rect 15752 17076 15804 17085
rect 16304 17076 16356 17128
rect 16580 17076 16632 17128
rect 13084 17008 13136 17017
rect 15384 17008 15436 17060
rect 15568 17051 15620 17060
rect 15568 17017 15577 17051
rect 15577 17017 15611 17051
rect 15611 17017 15620 17051
rect 22744 17187 22796 17196
rect 22744 17153 22753 17187
rect 22753 17153 22787 17187
rect 22787 17153 22796 17187
rect 22744 17144 22796 17153
rect 23572 17144 23624 17196
rect 19432 17119 19484 17128
rect 19432 17085 19441 17119
rect 19441 17085 19475 17119
rect 19475 17085 19484 17119
rect 19432 17076 19484 17085
rect 20996 17119 21048 17128
rect 20996 17085 21005 17119
rect 21005 17085 21039 17119
rect 21039 17085 21048 17119
rect 20996 17076 21048 17085
rect 22928 17119 22980 17128
rect 22928 17085 22937 17119
rect 22937 17085 22971 17119
rect 22971 17085 22980 17119
rect 22928 17076 22980 17085
rect 28356 17144 28408 17196
rect 27896 17076 27948 17128
rect 27988 17119 28040 17128
rect 27988 17085 27997 17119
rect 27997 17085 28031 17119
rect 28031 17085 28040 17119
rect 27988 17076 28040 17085
rect 29736 17119 29788 17128
rect 29736 17085 29745 17119
rect 29745 17085 29779 17119
rect 29779 17085 29788 17119
rect 29736 17076 29788 17085
rect 15568 17008 15620 17017
rect 18420 17008 18472 17060
rect 2964 16940 3016 16992
rect 3424 16983 3476 16992
rect 3424 16949 3433 16983
rect 3433 16949 3467 16983
rect 3467 16949 3476 16983
rect 3424 16940 3476 16949
rect 14280 16940 14332 16992
rect 15752 16940 15804 16992
rect 18052 16983 18104 16992
rect 18052 16949 18061 16983
rect 18061 16949 18095 16983
rect 18095 16949 18104 16983
rect 18052 16940 18104 16949
rect 21272 16983 21324 16992
rect 21272 16949 21281 16983
rect 21281 16949 21315 16983
rect 21315 16949 21324 16983
rect 21272 16940 21324 16949
rect 24952 16940 25004 16992
rect 26148 16983 26200 16992
rect 26148 16949 26157 16983
rect 26157 16949 26191 16983
rect 26191 16949 26200 16983
rect 26148 16940 26200 16949
rect 4664 16838 4716 16890
rect 4728 16838 4780 16890
rect 4792 16838 4844 16890
rect 4856 16838 4908 16890
rect 4920 16838 4972 16890
rect 12092 16838 12144 16890
rect 12156 16838 12208 16890
rect 12220 16838 12272 16890
rect 12284 16838 12336 16890
rect 12348 16838 12400 16890
rect 19520 16838 19572 16890
rect 19584 16838 19636 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 26948 16838 27000 16890
rect 27012 16838 27064 16890
rect 27076 16838 27128 16890
rect 27140 16838 27192 16890
rect 27204 16838 27256 16890
rect 11796 16779 11848 16788
rect 11796 16745 11805 16779
rect 11805 16745 11839 16779
rect 11839 16745 11848 16779
rect 11796 16736 11848 16745
rect 11888 16736 11940 16788
rect 12348 16736 12400 16788
rect 14372 16779 14424 16788
rect 14372 16745 14381 16779
rect 14381 16745 14415 16779
rect 14415 16745 14424 16779
rect 14372 16736 14424 16745
rect 2872 16668 2924 16720
rect 4712 16668 4764 16720
rect 2044 16532 2096 16584
rect 3976 16600 4028 16652
rect 9588 16600 9640 16652
rect 5724 16532 5776 16584
rect 6184 16575 6236 16584
rect 6184 16541 6193 16575
rect 6193 16541 6227 16575
rect 6227 16541 6236 16575
rect 6184 16532 6236 16541
rect 12348 16643 12400 16652
rect 12348 16609 12357 16643
rect 12357 16609 12391 16643
rect 12391 16609 12400 16643
rect 12348 16600 12400 16609
rect 13084 16600 13136 16652
rect 15568 16668 15620 16720
rect 16488 16668 16540 16720
rect 18420 16736 18472 16788
rect 27620 16736 27672 16788
rect 13544 16575 13596 16584
rect 13544 16541 13553 16575
rect 13553 16541 13587 16575
rect 13587 16541 13596 16575
rect 13544 16532 13596 16541
rect 13820 16600 13872 16652
rect 14280 16600 14332 16652
rect 6460 16507 6512 16516
rect 6460 16473 6469 16507
rect 6469 16473 6503 16507
rect 6503 16473 6512 16507
rect 6460 16464 6512 16473
rect 8300 16464 8352 16516
rect 9128 16439 9180 16448
rect 9128 16405 9137 16439
rect 9137 16405 9171 16439
rect 9171 16405 9180 16439
rect 9128 16396 9180 16405
rect 9496 16439 9548 16448
rect 9496 16405 9505 16439
rect 9505 16405 9539 16439
rect 9539 16405 9548 16439
rect 9496 16396 9548 16405
rect 15200 16600 15252 16652
rect 15476 16532 15528 16584
rect 16764 16600 16816 16652
rect 17040 16711 17092 16720
rect 17040 16677 17049 16711
rect 17049 16677 17083 16711
rect 17083 16677 17092 16711
rect 17040 16668 17092 16677
rect 17960 16668 18012 16720
rect 19432 16600 19484 16652
rect 19984 16643 20036 16652
rect 19984 16609 19993 16643
rect 19993 16609 20027 16643
rect 20027 16609 20036 16643
rect 19984 16600 20036 16609
rect 26148 16643 26200 16652
rect 26148 16609 26157 16643
rect 26157 16609 26191 16643
rect 26191 16609 26200 16643
rect 26148 16600 26200 16609
rect 26424 16643 26476 16652
rect 26424 16609 26433 16643
rect 26433 16609 26467 16643
rect 26467 16609 26476 16643
rect 26424 16600 26476 16609
rect 16212 16464 16264 16516
rect 16488 16464 16540 16516
rect 17868 16575 17920 16584
rect 17868 16541 17877 16575
rect 17877 16541 17911 16575
rect 17911 16541 17920 16575
rect 17868 16532 17920 16541
rect 22008 16532 22060 16584
rect 27896 16532 27948 16584
rect 28264 16532 28316 16584
rect 29644 16532 29696 16584
rect 23112 16464 23164 16516
rect 27436 16464 27488 16516
rect 15292 16396 15344 16448
rect 16120 16396 16172 16448
rect 18052 16396 18104 16448
rect 19432 16439 19484 16448
rect 19432 16405 19441 16439
rect 19441 16405 19475 16439
rect 19475 16405 19484 16439
rect 19432 16396 19484 16405
rect 19524 16396 19576 16448
rect 19892 16439 19944 16448
rect 19892 16405 19901 16439
rect 19901 16405 19935 16439
rect 19935 16405 19944 16439
rect 19892 16396 19944 16405
rect 28724 16396 28776 16448
rect 30012 16396 30064 16448
rect 8378 16294 8430 16346
rect 8442 16294 8494 16346
rect 8506 16294 8558 16346
rect 8570 16294 8622 16346
rect 8634 16294 8686 16346
rect 15806 16294 15858 16346
rect 15870 16294 15922 16346
rect 15934 16294 15986 16346
rect 15998 16294 16050 16346
rect 16062 16294 16114 16346
rect 23234 16294 23286 16346
rect 23298 16294 23350 16346
rect 23362 16294 23414 16346
rect 23426 16294 23478 16346
rect 23490 16294 23542 16346
rect 30662 16294 30714 16346
rect 30726 16294 30778 16346
rect 30790 16294 30842 16346
rect 30854 16294 30906 16346
rect 30918 16294 30970 16346
rect 2964 16167 3016 16176
rect 2964 16133 2973 16167
rect 2973 16133 3007 16167
rect 3007 16133 3016 16167
rect 2964 16124 3016 16133
rect 3424 16124 3476 16176
rect 4712 16167 4764 16176
rect 4712 16133 4721 16167
rect 4721 16133 4755 16167
rect 4755 16133 4764 16167
rect 4712 16124 4764 16133
rect 9128 16124 9180 16176
rect 10968 16235 11020 16244
rect 10968 16201 10977 16235
rect 10977 16201 11011 16235
rect 11011 16201 11020 16235
rect 10968 16192 11020 16201
rect 13544 16192 13596 16244
rect 15568 16192 15620 16244
rect 28264 16235 28316 16244
rect 28264 16201 28273 16235
rect 28273 16201 28307 16235
rect 28307 16201 28316 16235
rect 28264 16192 28316 16201
rect 11152 16124 11204 16176
rect 15660 16124 15712 16176
rect 19432 16124 19484 16176
rect 29736 16124 29788 16176
rect 3332 15988 3384 16040
rect 6184 15988 6236 16040
rect 9588 16056 9640 16108
rect 11612 16056 11664 16108
rect 15384 16099 15436 16108
rect 15384 16065 15393 16099
rect 15393 16065 15427 16099
rect 15427 16065 15436 16099
rect 15384 16056 15436 16065
rect 15568 16099 15620 16108
rect 15568 16065 15577 16099
rect 15577 16065 15611 16099
rect 15611 16065 15620 16099
rect 15568 16056 15620 16065
rect 16212 16099 16264 16108
rect 16212 16065 16221 16099
rect 16221 16065 16255 16099
rect 16255 16065 16264 16099
rect 16212 16056 16264 16065
rect 23756 16099 23808 16108
rect 23756 16065 23765 16099
rect 23765 16065 23799 16099
rect 23799 16065 23808 16099
rect 23756 16056 23808 16065
rect 24400 16056 24452 16108
rect 24768 16056 24820 16108
rect 30012 16099 30064 16108
rect 30012 16065 30021 16099
rect 30021 16065 30055 16099
rect 30055 16065 30064 16099
rect 30012 16056 30064 16065
rect 7288 15852 7340 15904
rect 8300 15895 8352 15904
rect 8300 15861 8309 15895
rect 8309 15861 8343 15895
rect 8343 15861 8352 15895
rect 8300 15852 8352 15861
rect 9312 15852 9364 15904
rect 11796 15988 11848 16040
rect 15108 15988 15160 16040
rect 16488 15988 16540 16040
rect 23664 15988 23716 16040
rect 24308 16031 24360 16040
rect 24308 15997 24317 16031
rect 24317 15997 24351 16031
rect 24351 15997 24360 16031
rect 24308 15988 24360 15997
rect 25964 15988 26016 16040
rect 28724 15988 28776 16040
rect 11888 15852 11940 15904
rect 13820 15920 13872 15972
rect 14004 15920 14056 15972
rect 14096 15852 14148 15904
rect 19892 15852 19944 15904
rect 24860 15852 24912 15904
rect 4664 15750 4716 15802
rect 4728 15750 4780 15802
rect 4792 15750 4844 15802
rect 4856 15750 4908 15802
rect 4920 15750 4972 15802
rect 12092 15750 12144 15802
rect 12156 15750 12208 15802
rect 12220 15750 12272 15802
rect 12284 15750 12336 15802
rect 12348 15750 12400 15802
rect 19520 15750 19572 15802
rect 19584 15750 19636 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 26948 15750 27000 15802
rect 27012 15750 27064 15802
rect 27076 15750 27128 15802
rect 27140 15750 27192 15802
rect 27204 15750 27256 15802
rect 6184 15691 6236 15700
rect 6184 15657 6193 15691
rect 6193 15657 6227 15691
rect 6227 15657 6236 15691
rect 6184 15648 6236 15657
rect 6460 15648 6512 15700
rect 6828 15648 6880 15700
rect 9128 15648 9180 15700
rect 9312 15648 9364 15700
rect 25964 15691 26016 15700
rect 25964 15657 25973 15691
rect 25973 15657 26007 15691
rect 26007 15657 26016 15691
rect 25964 15648 26016 15657
rect 11152 15580 11204 15632
rect 12624 15580 12676 15632
rect 5172 15444 5224 15496
rect 7288 15487 7340 15496
rect 7288 15453 7306 15487
rect 7306 15453 7340 15487
rect 7288 15444 7340 15453
rect 9036 15444 9088 15496
rect 12716 15512 12768 15564
rect 12808 15512 12860 15564
rect 15384 15580 15436 15632
rect 16580 15580 16632 15632
rect 19984 15580 20036 15632
rect 24308 15580 24360 15632
rect 9772 15376 9824 15428
rect 11980 15376 12032 15428
rect 13544 15444 13596 15496
rect 16212 15444 16264 15496
rect 16488 15444 16540 15496
rect 18604 15444 18656 15496
rect 13452 15376 13504 15428
rect 13820 15376 13872 15428
rect 16856 15419 16908 15428
rect 16856 15385 16890 15419
rect 16890 15385 16908 15419
rect 16856 15376 16908 15385
rect 18788 15376 18840 15428
rect 21456 15487 21508 15496
rect 21456 15453 21465 15487
rect 21465 15453 21499 15487
rect 21499 15453 21508 15487
rect 21456 15444 21508 15453
rect 22744 15444 22796 15496
rect 23756 15444 23808 15496
rect 24860 15487 24912 15496
rect 24860 15453 24894 15487
rect 24894 15453 24912 15487
rect 24860 15444 24912 15453
rect 29644 15512 29696 15564
rect 27988 15444 28040 15496
rect 28356 15444 28408 15496
rect 29184 15419 29236 15428
rect 29184 15385 29193 15419
rect 29193 15385 29227 15419
rect 29227 15385 29236 15419
rect 29184 15376 29236 15385
rect 4436 15308 4488 15360
rect 10232 15308 10284 15360
rect 12440 15308 12492 15360
rect 18604 15308 18656 15360
rect 20720 15308 20772 15360
rect 21088 15351 21140 15360
rect 21088 15317 21097 15351
rect 21097 15317 21131 15351
rect 21131 15317 21140 15351
rect 21088 15308 21140 15317
rect 21180 15308 21232 15360
rect 23572 15308 23624 15360
rect 24584 15308 24636 15360
rect 28172 15308 28224 15360
rect 8378 15206 8430 15258
rect 8442 15206 8494 15258
rect 8506 15206 8558 15258
rect 8570 15206 8622 15258
rect 8634 15206 8686 15258
rect 15806 15206 15858 15258
rect 15870 15206 15922 15258
rect 15934 15206 15986 15258
rect 15998 15206 16050 15258
rect 16062 15206 16114 15258
rect 23234 15206 23286 15258
rect 23298 15206 23350 15258
rect 23362 15206 23414 15258
rect 23426 15206 23478 15258
rect 23490 15206 23542 15258
rect 30662 15206 30714 15258
rect 30726 15206 30778 15258
rect 30790 15206 30842 15258
rect 30854 15206 30906 15258
rect 30918 15206 30970 15258
rect 8024 15147 8076 15156
rect 8024 15113 8033 15147
rect 8033 15113 8067 15147
rect 8067 15113 8076 15147
rect 8024 15104 8076 15113
rect 9772 15147 9824 15156
rect 9772 15113 9781 15147
rect 9781 15113 9815 15147
rect 9815 15113 9824 15147
rect 9772 15104 9824 15113
rect 10232 15147 10284 15156
rect 10232 15113 10241 15147
rect 10241 15113 10275 15147
rect 10275 15113 10284 15147
rect 10232 15104 10284 15113
rect 11060 15147 11112 15156
rect 11060 15113 11069 15147
rect 11069 15113 11103 15147
rect 11103 15113 11112 15147
rect 11060 15104 11112 15113
rect 11980 15104 12032 15156
rect 16856 15147 16908 15156
rect 16856 15113 16865 15147
rect 16865 15113 16899 15147
rect 16899 15113 16908 15147
rect 16856 15104 16908 15113
rect 22008 15104 22060 15156
rect 24584 15147 24636 15156
rect 24584 15113 24593 15147
rect 24593 15113 24627 15147
rect 24627 15113 24636 15147
rect 24584 15104 24636 15113
rect 29644 15147 29696 15156
rect 29644 15113 29653 15147
rect 29653 15113 29687 15147
rect 29687 15113 29696 15147
rect 29644 15104 29696 15113
rect 5264 15011 5316 15020
rect 5264 14977 5273 15011
rect 5273 14977 5307 15011
rect 5307 14977 5316 15011
rect 5264 14968 5316 14977
rect 6552 15011 6604 15020
rect 6552 14977 6561 15011
rect 6561 14977 6595 15011
rect 6595 14977 6604 15011
rect 6552 14968 6604 14977
rect 13176 15036 13228 15088
rect 14740 15036 14792 15088
rect 17132 15036 17184 15088
rect 18604 15079 18656 15088
rect 18604 15045 18613 15079
rect 18613 15045 18647 15079
rect 18647 15045 18656 15079
rect 18604 15036 18656 15045
rect 5356 14943 5408 14952
rect 5356 14909 5365 14943
rect 5365 14909 5399 14943
rect 5399 14909 5408 14943
rect 5356 14900 5408 14909
rect 5908 14943 5960 14952
rect 5908 14909 5917 14943
rect 5917 14909 5951 14943
rect 5951 14909 5960 14943
rect 5908 14900 5960 14909
rect 9588 14900 9640 14952
rect 11888 15011 11940 15020
rect 11888 14977 11897 15011
rect 11897 14977 11931 15011
rect 11931 14977 11940 15011
rect 11888 14968 11940 14977
rect 13452 14968 13504 15020
rect 13820 14900 13872 14952
rect 17224 15011 17276 15020
rect 17224 14977 17233 15011
rect 17233 14977 17267 15011
rect 17267 14977 17276 15011
rect 17224 14968 17276 14977
rect 17500 14968 17552 15020
rect 18788 15011 18840 15020
rect 18788 14977 18797 15011
rect 18797 14977 18831 15011
rect 18831 14977 18840 15011
rect 18788 14968 18840 14977
rect 20720 15079 20772 15088
rect 20720 15045 20729 15079
rect 20729 15045 20763 15079
rect 20763 15045 20772 15079
rect 20720 15036 20772 15045
rect 21088 15036 21140 15088
rect 23572 15036 23624 15088
rect 23664 15036 23716 15088
rect 28172 15079 28224 15088
rect 28172 15045 28181 15079
rect 28181 15045 28215 15079
rect 28215 15045 28224 15079
rect 28172 15036 28224 15045
rect 29184 15036 29236 15088
rect 15200 14900 15252 14952
rect 17040 14900 17092 14952
rect 17408 14943 17460 14952
rect 17408 14909 17417 14943
rect 17417 14909 17451 14943
rect 17451 14909 17460 14943
rect 17408 14900 17460 14909
rect 18604 14900 18656 14952
rect 19892 14900 19944 14952
rect 21180 14968 21232 15020
rect 21916 14968 21968 15020
rect 27804 14968 27856 15020
rect 11704 14764 11756 14816
rect 14648 14764 14700 14816
rect 14924 14764 14976 14816
rect 16212 14764 16264 14816
rect 20996 14832 21048 14884
rect 22468 14943 22520 14952
rect 22468 14909 22477 14943
rect 22477 14909 22511 14943
rect 22511 14909 22520 14943
rect 22468 14900 22520 14909
rect 25964 14900 26016 14952
rect 27896 14943 27948 14952
rect 27896 14909 27905 14943
rect 27905 14909 27939 14943
rect 27939 14909 27948 14943
rect 27896 14900 27948 14909
rect 17224 14764 17276 14816
rect 22744 14764 22796 14816
rect 25872 14764 25924 14816
rect 4664 14662 4716 14714
rect 4728 14662 4780 14714
rect 4792 14662 4844 14714
rect 4856 14662 4908 14714
rect 4920 14662 4972 14714
rect 12092 14662 12144 14714
rect 12156 14662 12208 14714
rect 12220 14662 12272 14714
rect 12284 14662 12336 14714
rect 12348 14662 12400 14714
rect 19520 14662 19572 14714
rect 19584 14662 19636 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 26948 14662 27000 14714
rect 27012 14662 27064 14714
rect 27076 14662 27128 14714
rect 27140 14662 27192 14714
rect 27204 14662 27256 14714
rect 6552 14560 6604 14612
rect 18512 14560 18564 14612
rect 20904 14560 20956 14612
rect 21272 14560 21324 14612
rect 21916 14603 21968 14612
rect 21916 14569 21925 14603
rect 21925 14569 21959 14603
rect 21959 14569 21968 14603
rect 21916 14560 21968 14569
rect 27896 14560 27948 14612
rect 10232 14492 10284 14544
rect 10968 14492 11020 14544
rect 10692 14424 10744 14476
rect 13176 14492 13228 14544
rect 13820 14492 13872 14544
rect 20996 14492 21048 14544
rect 14924 14467 14976 14476
rect 14924 14433 14933 14467
rect 14933 14433 14967 14467
rect 14967 14433 14976 14467
rect 14924 14424 14976 14433
rect 17132 14424 17184 14476
rect 4620 14399 4672 14408
rect 4620 14365 4629 14399
rect 4629 14365 4663 14399
rect 4663 14365 4672 14399
rect 4620 14356 4672 14365
rect 5908 14288 5960 14340
rect 6736 14288 6788 14340
rect 9404 14399 9456 14408
rect 9404 14365 9413 14399
rect 9413 14365 9447 14399
rect 9447 14365 9456 14399
rect 9404 14356 9456 14365
rect 11612 14356 11664 14408
rect 11796 14399 11848 14408
rect 11796 14365 11805 14399
rect 11805 14365 11839 14399
rect 11839 14365 11848 14399
rect 11796 14356 11848 14365
rect 11520 14263 11572 14272
rect 11520 14229 11529 14263
rect 11529 14229 11563 14263
rect 11563 14229 11572 14263
rect 11520 14220 11572 14229
rect 12440 14356 12492 14408
rect 14188 14356 14240 14408
rect 20904 14424 20956 14476
rect 24400 14424 24452 14476
rect 24584 14424 24636 14476
rect 25596 14424 25648 14476
rect 12072 14288 12124 14340
rect 15568 14288 15620 14340
rect 16764 14288 16816 14340
rect 19984 14288 20036 14340
rect 12440 14220 12492 14272
rect 16304 14263 16356 14272
rect 16304 14229 16313 14263
rect 16313 14229 16347 14263
rect 16347 14229 16356 14263
rect 16304 14220 16356 14229
rect 16488 14220 16540 14272
rect 20904 14220 20956 14272
rect 20996 14263 21048 14272
rect 20996 14229 21005 14263
rect 21005 14229 21039 14263
rect 21039 14229 21048 14263
rect 20996 14220 21048 14229
rect 21456 14331 21508 14340
rect 21456 14297 21465 14331
rect 21465 14297 21499 14331
rect 21499 14297 21508 14331
rect 21456 14288 21508 14297
rect 21548 14288 21600 14340
rect 21732 14399 21784 14408
rect 21732 14365 21741 14399
rect 21741 14365 21775 14399
rect 21775 14365 21784 14399
rect 21732 14356 21784 14365
rect 24768 14399 24820 14408
rect 24768 14365 24777 14399
rect 24777 14365 24811 14399
rect 24811 14365 24820 14399
rect 24768 14356 24820 14365
rect 27804 14356 27856 14408
rect 25688 14288 25740 14340
rect 28724 14399 28776 14408
rect 28724 14365 28733 14399
rect 28733 14365 28767 14399
rect 28767 14365 28776 14399
rect 28724 14356 28776 14365
rect 30288 14399 30340 14408
rect 30288 14365 30297 14399
rect 30297 14365 30331 14399
rect 30331 14365 30340 14399
rect 30288 14356 30340 14365
rect 29644 14288 29696 14340
rect 31024 14288 31076 14340
rect 23756 14220 23808 14272
rect 27528 14220 27580 14272
rect 28632 14263 28684 14272
rect 28632 14229 28641 14263
rect 28641 14229 28675 14263
rect 28675 14229 28684 14263
rect 28632 14220 28684 14229
rect 8378 14118 8430 14170
rect 8442 14118 8494 14170
rect 8506 14118 8558 14170
rect 8570 14118 8622 14170
rect 8634 14118 8686 14170
rect 15806 14118 15858 14170
rect 15870 14118 15922 14170
rect 15934 14118 15986 14170
rect 15998 14118 16050 14170
rect 16062 14118 16114 14170
rect 23234 14118 23286 14170
rect 23298 14118 23350 14170
rect 23362 14118 23414 14170
rect 23426 14118 23478 14170
rect 23490 14118 23542 14170
rect 30662 14118 30714 14170
rect 30726 14118 30778 14170
rect 30790 14118 30842 14170
rect 30854 14118 30906 14170
rect 30918 14118 30970 14170
rect 4620 14016 4672 14068
rect 5172 14016 5224 14068
rect 9404 14016 9456 14068
rect 14188 14059 14240 14068
rect 14188 14025 14197 14059
rect 14197 14025 14231 14059
rect 14231 14025 14240 14059
rect 14188 14016 14240 14025
rect 15568 14059 15620 14068
rect 15568 14025 15577 14059
rect 15577 14025 15611 14059
rect 15611 14025 15620 14059
rect 15568 14016 15620 14025
rect 16304 14016 16356 14068
rect 16396 14016 16448 14068
rect 17224 14059 17276 14068
rect 17224 14025 17233 14059
rect 17233 14025 17267 14059
rect 17267 14025 17276 14059
rect 17224 14016 17276 14025
rect 19984 14059 20036 14068
rect 19984 14025 19993 14059
rect 19993 14025 20027 14059
rect 20027 14025 20036 14059
rect 19984 14016 20036 14025
rect 20996 14016 21048 14068
rect 22468 14016 22520 14068
rect 29644 14016 29696 14068
rect 4436 13991 4488 14000
rect 4436 13957 4445 13991
rect 4445 13957 4479 13991
rect 4479 13957 4488 13991
rect 4436 13948 4488 13957
rect 5816 13948 5868 14000
rect 6736 13923 6788 13932
rect 6736 13889 6745 13923
rect 6745 13889 6779 13923
rect 6779 13889 6788 13923
rect 6736 13880 6788 13889
rect 11888 13880 11940 13932
rect 12532 13923 12584 13932
rect 12532 13889 12566 13923
rect 12566 13889 12584 13923
rect 12532 13880 12584 13889
rect 14096 13923 14148 13932
rect 14096 13889 14105 13923
rect 14105 13889 14139 13923
rect 14139 13889 14148 13923
rect 14096 13880 14148 13889
rect 14924 13880 14976 13932
rect 16488 13880 16540 13932
rect 17500 13880 17552 13932
rect 20444 13880 20496 13932
rect 21732 13880 21784 13932
rect 4160 13855 4212 13864
rect 4160 13821 4169 13855
rect 4169 13821 4203 13855
rect 4203 13821 4212 13855
rect 4160 13812 4212 13821
rect 6184 13812 6236 13864
rect 7196 13812 7248 13864
rect 17316 13855 17368 13864
rect 17316 13821 17325 13855
rect 17325 13821 17359 13855
rect 17359 13821 17368 13855
rect 17316 13812 17368 13821
rect 17408 13855 17460 13864
rect 17408 13821 17417 13855
rect 17417 13821 17451 13855
rect 17451 13821 17460 13855
rect 17408 13812 17460 13821
rect 23112 13948 23164 14000
rect 25596 13991 25648 14000
rect 25596 13957 25605 13991
rect 25605 13957 25639 13991
rect 25639 13957 25648 13991
rect 25596 13948 25648 13957
rect 23020 13880 23072 13932
rect 25872 13923 25924 13932
rect 25872 13889 25881 13923
rect 25881 13889 25915 13923
rect 25915 13889 25924 13923
rect 25872 13880 25924 13889
rect 13176 13676 13228 13728
rect 20076 13744 20128 13796
rect 24768 13744 24820 13796
rect 26516 13880 26568 13932
rect 28632 13948 28684 14000
rect 29736 13880 29788 13932
rect 28632 13855 28684 13864
rect 28632 13821 28641 13855
rect 28641 13821 28675 13855
rect 28675 13821 28684 13855
rect 28632 13812 28684 13821
rect 24584 13676 24636 13728
rect 24952 13676 25004 13728
rect 27344 13676 27396 13728
rect 4664 13574 4716 13626
rect 4728 13574 4780 13626
rect 4792 13574 4844 13626
rect 4856 13574 4908 13626
rect 4920 13574 4972 13626
rect 12092 13574 12144 13626
rect 12156 13574 12208 13626
rect 12220 13574 12272 13626
rect 12284 13574 12336 13626
rect 12348 13574 12400 13626
rect 19520 13574 19572 13626
rect 19584 13574 19636 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 26948 13574 27000 13626
rect 27012 13574 27064 13626
rect 27076 13574 27128 13626
rect 27140 13574 27192 13626
rect 27204 13574 27256 13626
rect 4160 13472 4212 13524
rect 12532 13472 12584 13524
rect 20444 13472 20496 13524
rect 21548 13472 21600 13524
rect 28632 13472 28684 13524
rect 28724 13447 28776 13456
rect 28724 13413 28733 13447
rect 28733 13413 28767 13447
rect 28767 13413 28776 13447
rect 28724 13404 28776 13413
rect 5264 13336 5316 13388
rect 9128 13379 9180 13388
rect 9128 13345 9137 13379
rect 9137 13345 9171 13379
rect 9171 13345 9180 13379
rect 9128 13336 9180 13345
rect 13176 13379 13228 13388
rect 13176 13345 13185 13379
rect 13185 13345 13219 13379
rect 13219 13345 13228 13379
rect 13176 13336 13228 13345
rect 13268 13336 13320 13388
rect 15108 13336 15160 13388
rect 17316 13336 17368 13388
rect 20996 13336 21048 13388
rect 27344 13336 27396 13388
rect 4988 13268 5040 13320
rect 8024 13268 8076 13320
rect 16212 13311 16264 13320
rect 16212 13277 16221 13311
rect 16221 13277 16255 13311
rect 16255 13277 16264 13311
rect 16212 13268 16264 13277
rect 18236 13311 18288 13320
rect 18236 13277 18245 13311
rect 18245 13277 18279 13311
rect 18279 13277 18288 13311
rect 18236 13268 18288 13277
rect 22928 13268 22980 13320
rect 24768 13268 24820 13320
rect 29644 13268 29696 13320
rect 9220 13200 9272 13252
rect 9496 13200 9548 13252
rect 9588 13132 9640 13184
rect 13360 13200 13412 13252
rect 16856 13200 16908 13252
rect 24584 13243 24636 13252
rect 24584 13209 24593 13243
rect 24593 13209 24627 13243
rect 24627 13209 24636 13243
rect 24584 13200 24636 13209
rect 27528 13200 27580 13252
rect 28264 13200 28316 13252
rect 17500 13132 17552 13184
rect 17592 13175 17644 13184
rect 17592 13141 17601 13175
rect 17601 13141 17635 13175
rect 17635 13141 17644 13175
rect 17592 13132 17644 13141
rect 25044 13132 25096 13184
rect 26056 13175 26108 13184
rect 26056 13141 26065 13175
rect 26065 13141 26099 13175
rect 26099 13141 26108 13175
rect 26056 13132 26108 13141
rect 8378 13030 8430 13082
rect 8442 13030 8494 13082
rect 8506 13030 8558 13082
rect 8570 13030 8622 13082
rect 8634 13030 8686 13082
rect 15806 13030 15858 13082
rect 15870 13030 15922 13082
rect 15934 13030 15986 13082
rect 15998 13030 16050 13082
rect 16062 13030 16114 13082
rect 23234 13030 23286 13082
rect 23298 13030 23350 13082
rect 23362 13030 23414 13082
rect 23426 13030 23478 13082
rect 23490 13030 23542 13082
rect 30662 13030 30714 13082
rect 30726 13030 30778 13082
rect 30790 13030 30842 13082
rect 30854 13030 30906 13082
rect 30918 13030 30970 13082
rect 5816 12971 5868 12980
rect 5816 12937 5825 12971
rect 5825 12937 5859 12971
rect 5859 12937 5868 12971
rect 5816 12928 5868 12937
rect 9220 12971 9272 12980
rect 9220 12937 9229 12971
rect 9229 12937 9263 12971
rect 9263 12937 9272 12971
rect 9220 12928 9272 12937
rect 9588 12928 9640 12980
rect 6920 12860 6972 12912
rect 5264 12792 5316 12844
rect 5356 12835 5408 12844
rect 5356 12801 5365 12835
rect 5365 12801 5399 12835
rect 5399 12801 5408 12835
rect 5356 12792 5408 12801
rect 7104 12792 7156 12844
rect 7656 12792 7708 12844
rect 9496 12792 9548 12844
rect 16856 12971 16908 12980
rect 16856 12937 16865 12971
rect 16865 12937 16899 12971
rect 16899 12937 16908 12971
rect 16856 12928 16908 12937
rect 26056 12928 26108 12980
rect 25044 12903 25096 12912
rect 25044 12869 25053 12903
rect 25053 12869 25087 12903
rect 25087 12869 25096 12903
rect 25044 12860 25096 12869
rect 5448 12724 5500 12776
rect 8300 12767 8352 12776
rect 8300 12733 8309 12767
rect 8309 12733 8343 12767
rect 8343 12733 8352 12767
rect 8300 12724 8352 12733
rect 9128 12656 9180 12708
rect 11888 12724 11940 12776
rect 14924 12792 14976 12844
rect 12808 12656 12860 12708
rect 17592 12792 17644 12844
rect 15108 12656 15160 12708
rect 17408 12767 17460 12776
rect 17408 12733 17417 12767
rect 17417 12733 17451 12767
rect 17451 12733 17460 12767
rect 17408 12724 17460 12733
rect 19892 12792 19944 12844
rect 22928 12835 22980 12844
rect 22928 12801 22937 12835
rect 22937 12801 22971 12835
rect 22971 12801 22980 12835
rect 22928 12792 22980 12801
rect 23112 12792 23164 12844
rect 21456 12724 21508 12776
rect 23940 12724 23992 12776
rect 26148 12792 26200 12844
rect 27436 12835 27488 12844
rect 27436 12801 27445 12835
rect 27445 12801 27479 12835
rect 27479 12801 27488 12835
rect 27436 12792 27488 12801
rect 28264 12860 28316 12912
rect 29736 12903 29788 12912
rect 29736 12869 29745 12903
rect 29745 12869 29779 12903
rect 29779 12869 29788 12903
rect 29736 12860 29788 12869
rect 28356 12792 28408 12844
rect 26516 12767 26568 12776
rect 26516 12733 26525 12767
rect 26525 12733 26559 12767
rect 26559 12733 26568 12767
rect 26516 12724 26568 12733
rect 27988 12724 28040 12776
rect 17776 12656 17828 12708
rect 19432 12656 19484 12708
rect 7840 12588 7892 12640
rect 10416 12588 10468 12640
rect 22468 12588 22520 12640
rect 23480 12631 23532 12640
rect 23480 12597 23489 12631
rect 23489 12597 23523 12631
rect 23523 12597 23532 12631
rect 23480 12588 23532 12597
rect 25044 12588 25096 12640
rect 4664 12486 4716 12538
rect 4728 12486 4780 12538
rect 4792 12486 4844 12538
rect 4856 12486 4908 12538
rect 4920 12486 4972 12538
rect 12092 12486 12144 12538
rect 12156 12486 12208 12538
rect 12220 12486 12272 12538
rect 12284 12486 12336 12538
rect 12348 12486 12400 12538
rect 19520 12486 19572 12538
rect 19584 12486 19636 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 26948 12486 27000 12538
rect 27012 12486 27064 12538
rect 27076 12486 27128 12538
rect 27140 12486 27192 12538
rect 27204 12486 27256 12538
rect 17316 12384 17368 12436
rect 4988 12223 5040 12232
rect 4988 12189 4997 12223
rect 4997 12189 5031 12223
rect 5031 12189 5040 12223
rect 4988 12180 5040 12189
rect 5172 12180 5224 12232
rect 6920 12223 6972 12232
rect 6920 12189 6929 12223
rect 6929 12189 6963 12223
rect 6963 12189 6972 12223
rect 6920 12180 6972 12189
rect 7104 12223 7156 12232
rect 7104 12189 7113 12223
rect 7113 12189 7147 12223
rect 7147 12189 7156 12223
rect 7104 12180 7156 12189
rect 7196 12180 7248 12232
rect 23480 12384 23532 12436
rect 23940 12427 23992 12436
rect 23940 12393 23949 12427
rect 23949 12393 23983 12427
rect 23983 12393 23992 12427
rect 23940 12384 23992 12393
rect 22468 12291 22520 12300
rect 22468 12257 22477 12291
rect 22477 12257 22511 12291
rect 22511 12257 22520 12291
rect 22468 12248 22520 12257
rect 22928 12248 22980 12300
rect 27436 12316 27488 12368
rect 26148 12291 26200 12300
rect 26148 12257 26157 12291
rect 26157 12257 26191 12291
rect 26191 12257 26200 12291
rect 26148 12248 26200 12257
rect 7840 12223 7892 12232
rect 7840 12189 7849 12223
rect 7849 12189 7883 12223
rect 7883 12189 7892 12223
rect 7840 12180 7892 12189
rect 8116 12180 8168 12232
rect 4160 12112 4212 12164
rect 7932 12155 7984 12164
rect 7932 12121 7941 12155
rect 7941 12121 7975 12155
rect 7975 12121 7984 12155
rect 7932 12112 7984 12121
rect 4436 12044 4488 12096
rect 11796 12180 11848 12232
rect 12440 12180 12492 12232
rect 16396 12180 16448 12232
rect 18236 12180 18288 12232
rect 26056 12180 26108 12232
rect 16212 12112 16264 12164
rect 23756 12112 23808 12164
rect 12532 12044 12584 12096
rect 17316 12044 17368 12096
rect 8378 11942 8430 11994
rect 8442 11942 8494 11994
rect 8506 11942 8558 11994
rect 8570 11942 8622 11994
rect 8634 11942 8686 11994
rect 15806 11942 15858 11994
rect 15870 11942 15922 11994
rect 15934 11942 15986 11994
rect 15998 11942 16050 11994
rect 16062 11942 16114 11994
rect 23234 11942 23286 11994
rect 23298 11942 23350 11994
rect 23362 11942 23414 11994
rect 23426 11942 23478 11994
rect 23490 11942 23542 11994
rect 30662 11942 30714 11994
rect 30726 11942 30778 11994
rect 30790 11942 30842 11994
rect 30854 11942 30906 11994
rect 30918 11942 30970 11994
rect 4436 11815 4488 11824
rect 4436 11781 4445 11815
rect 4445 11781 4479 11815
rect 4479 11781 4488 11815
rect 4436 11772 4488 11781
rect 5724 11772 5776 11824
rect 4160 11747 4212 11756
rect 4160 11713 4169 11747
rect 4169 11713 4203 11747
rect 4203 11713 4212 11747
rect 4160 11704 4212 11713
rect 4988 11636 5040 11688
rect 7656 11840 7708 11892
rect 7932 11840 7984 11892
rect 12624 11840 12676 11892
rect 12808 11840 12860 11892
rect 7564 11704 7616 11756
rect 7840 11704 7892 11756
rect 6828 11679 6880 11688
rect 6828 11645 6837 11679
rect 6837 11645 6871 11679
rect 6871 11645 6880 11679
rect 6828 11636 6880 11645
rect 8024 11568 8076 11620
rect 8944 11704 8996 11756
rect 9680 11704 9732 11756
rect 10692 11747 10744 11756
rect 10692 11713 10701 11747
rect 10701 11713 10735 11747
rect 10735 11713 10744 11747
rect 10692 11704 10744 11713
rect 18236 11772 18288 11824
rect 17776 11704 17828 11756
rect 18512 11747 18564 11756
rect 18512 11713 18521 11747
rect 18521 11713 18555 11747
rect 18555 11713 18564 11747
rect 18512 11704 18564 11713
rect 23756 11772 23808 11824
rect 19892 11747 19944 11756
rect 19892 11713 19901 11747
rect 19901 11713 19935 11747
rect 19935 11713 19944 11747
rect 19892 11704 19944 11713
rect 20444 11704 20496 11756
rect 9496 11679 9548 11688
rect 9496 11645 9505 11679
rect 9505 11645 9539 11679
rect 9539 11645 9548 11679
rect 9496 11636 9548 11645
rect 13084 11679 13136 11688
rect 13084 11645 13093 11679
rect 13093 11645 13127 11679
rect 13127 11645 13136 11679
rect 13084 11636 13136 11645
rect 13268 11679 13320 11688
rect 13268 11645 13277 11679
rect 13277 11645 13311 11679
rect 13311 11645 13320 11679
rect 13268 11636 13320 11645
rect 17868 11679 17920 11688
rect 17868 11645 17877 11679
rect 17877 11645 17911 11679
rect 17911 11645 17920 11679
rect 17868 11636 17920 11645
rect 22928 11747 22980 11756
rect 22928 11713 22937 11747
rect 22937 11713 22971 11747
rect 22971 11713 22980 11747
rect 22928 11704 22980 11713
rect 23020 11704 23072 11756
rect 23112 11568 23164 11620
rect 10416 11543 10468 11552
rect 10416 11509 10425 11543
rect 10425 11509 10459 11543
rect 10459 11509 10468 11543
rect 10416 11500 10468 11509
rect 11980 11500 12032 11552
rect 12624 11543 12676 11552
rect 12624 11509 12633 11543
rect 12633 11509 12667 11543
rect 12667 11509 12676 11543
rect 12624 11500 12676 11509
rect 19432 11500 19484 11552
rect 19892 11500 19944 11552
rect 21732 11500 21784 11552
rect 22008 11500 22060 11552
rect 4664 11398 4716 11450
rect 4728 11398 4780 11450
rect 4792 11398 4844 11450
rect 4856 11398 4908 11450
rect 4920 11398 4972 11450
rect 12092 11398 12144 11450
rect 12156 11398 12208 11450
rect 12220 11398 12272 11450
rect 12284 11398 12336 11450
rect 12348 11398 12400 11450
rect 19520 11398 19572 11450
rect 19584 11398 19636 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 26948 11398 27000 11450
rect 27012 11398 27064 11450
rect 27076 11398 27128 11450
rect 27140 11398 27192 11450
rect 27204 11398 27256 11450
rect 7564 11339 7616 11348
rect 7564 11305 7573 11339
rect 7573 11305 7607 11339
rect 7607 11305 7616 11339
rect 7564 11296 7616 11305
rect 12072 11296 12124 11348
rect 13084 11296 13136 11348
rect 18236 11296 18288 11348
rect 20444 11296 20496 11348
rect 23112 11296 23164 11348
rect 29000 11271 29052 11280
rect 29000 11237 29009 11271
rect 29009 11237 29043 11271
rect 29043 11237 29052 11271
rect 29000 11228 29052 11237
rect 30288 11271 30340 11280
rect 30288 11237 30297 11271
rect 30297 11237 30331 11271
rect 30331 11237 30340 11271
rect 30288 11228 30340 11237
rect 5172 11160 5224 11212
rect 5264 11203 5316 11212
rect 5264 11169 5273 11203
rect 5273 11169 5307 11203
rect 5307 11169 5316 11203
rect 5264 11160 5316 11169
rect 5540 11160 5592 11212
rect 5724 11203 5776 11212
rect 5724 11169 5733 11203
rect 5733 11169 5767 11203
rect 5767 11169 5776 11203
rect 5724 11160 5776 11169
rect 8024 11203 8076 11212
rect 8024 11169 8033 11203
rect 8033 11169 8067 11203
rect 8067 11169 8076 11203
rect 8024 11160 8076 11169
rect 8208 11203 8260 11212
rect 8208 11169 8217 11203
rect 8217 11169 8251 11203
rect 8251 11169 8260 11203
rect 8208 11160 8260 11169
rect 9128 11160 9180 11212
rect 11888 11160 11940 11212
rect 17316 11160 17368 11212
rect 19432 11203 19484 11212
rect 19432 11169 19441 11203
rect 19441 11169 19475 11203
rect 19475 11169 19484 11203
rect 19432 11160 19484 11169
rect 19800 11160 19852 11212
rect 21732 11203 21784 11212
rect 21732 11169 21741 11203
rect 21741 11169 21775 11203
rect 21775 11169 21784 11203
rect 21732 11160 21784 11169
rect 22008 11203 22060 11212
rect 22008 11169 22017 11203
rect 22017 11169 22051 11203
rect 22051 11169 22060 11203
rect 22008 11160 22060 11169
rect 23664 11160 23716 11212
rect 24768 11160 24820 11212
rect 4252 11135 4304 11144
rect 4252 11101 4261 11135
rect 4261 11101 4295 11135
rect 4295 11101 4304 11135
rect 4252 11092 4304 11101
rect 5448 11092 5500 11144
rect 5632 11092 5684 11144
rect 9864 11135 9916 11144
rect 9864 11101 9873 11135
rect 9873 11101 9907 11135
rect 9907 11101 9916 11135
rect 9864 11092 9916 11101
rect 12624 11092 12676 11144
rect 5724 11024 5776 11076
rect 14924 11024 14976 11076
rect 10048 10956 10100 11008
rect 23112 11092 23164 11144
rect 24676 11135 24728 11144
rect 24676 11101 24685 11135
rect 24685 11101 24719 11135
rect 24719 11101 24728 11135
rect 24676 11092 24728 11101
rect 25412 11160 25464 11212
rect 25688 11135 25740 11144
rect 25688 11101 25697 11135
rect 25697 11101 25731 11135
rect 25731 11101 25740 11135
rect 25688 11092 25740 11101
rect 29828 11203 29880 11212
rect 29828 11169 29837 11203
rect 29837 11169 29871 11203
rect 29871 11169 29880 11203
rect 29828 11160 29880 11169
rect 17960 11024 18012 11076
rect 20720 11024 20772 11076
rect 26516 11024 26568 11076
rect 28724 11067 28776 11076
rect 28724 11033 28733 11067
rect 28733 11033 28767 11067
rect 28767 11033 28776 11067
rect 28724 11024 28776 11033
rect 16304 10956 16356 11008
rect 18604 10956 18656 11008
rect 24860 10999 24912 11008
rect 24860 10965 24869 10999
rect 24869 10965 24903 10999
rect 24903 10965 24912 10999
rect 24860 10956 24912 10965
rect 25320 10999 25372 11008
rect 25320 10965 25329 10999
rect 25329 10965 25363 10999
rect 25363 10965 25372 10999
rect 25320 10956 25372 10965
rect 8378 10854 8430 10906
rect 8442 10854 8494 10906
rect 8506 10854 8558 10906
rect 8570 10854 8622 10906
rect 8634 10854 8686 10906
rect 15806 10854 15858 10906
rect 15870 10854 15922 10906
rect 15934 10854 15986 10906
rect 15998 10854 16050 10906
rect 16062 10854 16114 10906
rect 23234 10854 23286 10906
rect 23298 10854 23350 10906
rect 23362 10854 23414 10906
rect 23426 10854 23478 10906
rect 23490 10854 23542 10906
rect 30662 10854 30714 10906
rect 30726 10854 30778 10906
rect 30790 10854 30842 10906
rect 30854 10854 30906 10906
rect 30918 10854 30970 10906
rect 4252 10795 4304 10804
rect 4252 10761 4261 10795
rect 4261 10761 4295 10795
rect 4295 10761 4304 10795
rect 4252 10752 4304 10761
rect 8116 10752 8168 10804
rect 12440 10752 12492 10804
rect 18604 10795 18656 10804
rect 18604 10761 18613 10795
rect 18613 10761 18647 10795
rect 18647 10761 18656 10795
rect 18604 10752 18656 10761
rect 24860 10752 24912 10804
rect 4988 10684 5040 10736
rect 5724 10727 5776 10736
rect 5724 10693 5733 10727
rect 5733 10693 5767 10727
rect 5767 10693 5776 10727
rect 5724 10684 5776 10693
rect 7840 10684 7892 10736
rect 8024 10684 8076 10736
rect 11520 10684 11572 10736
rect 11980 10684 12032 10736
rect 18144 10684 18196 10736
rect 20720 10684 20772 10736
rect 23112 10727 23164 10736
rect 23112 10693 23121 10727
rect 23121 10693 23155 10727
rect 23155 10693 23164 10727
rect 23112 10684 23164 10693
rect 25320 10684 25372 10736
rect 27436 10684 27488 10736
rect 27988 10684 28040 10736
rect 29828 10752 29880 10804
rect 11152 10659 11204 10668
rect 11152 10625 11161 10659
rect 11161 10625 11195 10659
rect 11195 10625 11204 10659
rect 11152 10616 11204 10625
rect 12900 10616 12952 10668
rect 14280 10616 14332 10668
rect 16304 10659 16356 10668
rect 16304 10625 16313 10659
rect 16313 10625 16347 10659
rect 16347 10625 16356 10659
rect 16304 10616 16356 10625
rect 16764 10616 16816 10668
rect 19984 10616 20036 10668
rect 23020 10616 23072 10668
rect 24768 10659 24820 10668
rect 24768 10625 24777 10659
rect 24777 10625 24811 10659
rect 24811 10625 24820 10659
rect 24768 10616 24820 10625
rect 28172 10616 28224 10668
rect 29000 10684 29052 10736
rect 29920 10684 29972 10736
rect 28724 10659 28776 10668
rect 28724 10625 28733 10659
rect 28733 10625 28767 10659
rect 28767 10625 28776 10659
rect 28724 10616 28776 10625
rect 9864 10548 9916 10600
rect 12532 10548 12584 10600
rect 12716 10548 12768 10600
rect 17868 10548 17920 10600
rect 22928 10548 22980 10600
rect 26516 10591 26568 10600
rect 26516 10557 26525 10591
rect 26525 10557 26559 10591
rect 26559 10557 26568 10591
rect 26516 10548 26568 10557
rect 27712 10548 27764 10600
rect 28908 10659 28960 10668
rect 28908 10625 28917 10659
rect 28917 10625 28951 10659
rect 28951 10625 28960 10659
rect 28908 10616 28960 10625
rect 29736 10548 29788 10600
rect 9220 10455 9272 10464
rect 9220 10421 9229 10455
rect 9229 10421 9263 10455
rect 9263 10421 9272 10455
rect 9220 10412 9272 10421
rect 9772 10412 9824 10464
rect 12440 10455 12492 10464
rect 12440 10421 12449 10455
rect 12449 10421 12483 10455
rect 12483 10421 12492 10455
rect 12440 10412 12492 10421
rect 14556 10455 14608 10464
rect 14556 10421 14565 10455
rect 14565 10421 14599 10455
rect 14599 10421 14608 10455
rect 14556 10412 14608 10421
rect 4664 10310 4716 10362
rect 4728 10310 4780 10362
rect 4792 10310 4844 10362
rect 4856 10310 4908 10362
rect 4920 10310 4972 10362
rect 12092 10310 12144 10362
rect 12156 10310 12208 10362
rect 12220 10310 12272 10362
rect 12284 10310 12336 10362
rect 12348 10310 12400 10362
rect 19520 10310 19572 10362
rect 19584 10310 19636 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 26948 10310 27000 10362
rect 27012 10310 27064 10362
rect 27076 10310 27128 10362
rect 27140 10310 27192 10362
rect 27204 10310 27256 10362
rect 5540 10251 5592 10260
rect 5540 10217 5549 10251
rect 5549 10217 5583 10251
rect 5583 10217 5592 10251
rect 5540 10208 5592 10217
rect 9864 10208 9916 10260
rect 12072 10208 12124 10260
rect 12532 10251 12584 10260
rect 12532 10217 12541 10251
rect 12541 10217 12575 10251
rect 12575 10217 12584 10251
rect 12532 10208 12584 10217
rect 14280 10251 14332 10260
rect 14280 10217 14289 10251
rect 14289 10217 14323 10251
rect 14323 10217 14332 10251
rect 14280 10208 14332 10217
rect 17868 10208 17920 10260
rect 19984 10208 20036 10260
rect 23020 10208 23072 10260
rect 28724 10208 28776 10260
rect 29736 10251 29788 10260
rect 29736 10217 29745 10251
rect 29745 10217 29779 10251
rect 29779 10217 29788 10251
rect 29736 10208 29788 10217
rect 8208 10115 8260 10124
rect 8208 10081 8217 10115
rect 8217 10081 8251 10115
rect 8251 10081 8260 10115
rect 8208 10072 8260 10081
rect 9772 10115 9824 10124
rect 9772 10081 9781 10115
rect 9781 10081 9815 10115
rect 9815 10081 9824 10115
rect 9772 10072 9824 10081
rect 10048 10115 10100 10124
rect 10048 10081 10057 10115
rect 10057 10081 10091 10115
rect 10091 10081 10100 10115
rect 10048 10072 10100 10081
rect 14556 10072 14608 10124
rect 15108 10072 15160 10124
rect 17960 10072 18012 10124
rect 9220 9936 9272 9988
rect 11336 10004 11388 10056
rect 12532 10004 12584 10056
rect 14648 10047 14700 10056
rect 14648 10013 14657 10047
rect 14657 10013 14691 10047
rect 14691 10013 14700 10047
rect 14648 10004 14700 10013
rect 17592 10004 17644 10056
rect 30012 10140 30064 10192
rect 25412 10072 25464 10124
rect 24584 10004 24636 10056
rect 25044 10004 25096 10056
rect 27988 10004 28040 10056
rect 28172 10047 28224 10056
rect 28172 10013 28181 10047
rect 28181 10013 28215 10047
rect 28215 10013 28224 10047
rect 28172 10004 28224 10013
rect 7656 9911 7708 9920
rect 7656 9877 7665 9911
rect 7665 9877 7699 9911
rect 7699 9877 7708 9911
rect 7656 9868 7708 9877
rect 8300 9868 8352 9920
rect 11060 9936 11112 9988
rect 27712 9936 27764 9988
rect 12808 9868 12860 9920
rect 24860 9868 24912 9920
rect 26056 9868 26108 9920
rect 27436 9868 27488 9920
rect 30196 9979 30248 9988
rect 30196 9945 30205 9979
rect 30205 9945 30239 9979
rect 30239 9945 30248 9979
rect 30196 9936 30248 9945
rect 29000 9911 29052 9920
rect 29000 9877 29009 9911
rect 29009 9877 29043 9911
rect 29043 9877 29052 9911
rect 29000 9868 29052 9877
rect 8378 9766 8430 9818
rect 8442 9766 8494 9818
rect 8506 9766 8558 9818
rect 8570 9766 8622 9818
rect 8634 9766 8686 9818
rect 15806 9766 15858 9818
rect 15870 9766 15922 9818
rect 15934 9766 15986 9818
rect 15998 9766 16050 9818
rect 16062 9766 16114 9818
rect 23234 9766 23286 9818
rect 23298 9766 23350 9818
rect 23362 9766 23414 9818
rect 23426 9766 23478 9818
rect 23490 9766 23542 9818
rect 30662 9766 30714 9818
rect 30726 9766 30778 9818
rect 30790 9766 30842 9818
rect 30854 9766 30906 9818
rect 30918 9766 30970 9818
rect 8300 9664 8352 9716
rect 8392 9707 8444 9716
rect 8392 9673 8401 9707
rect 8401 9673 8435 9707
rect 8435 9673 8444 9707
rect 8392 9664 8444 9673
rect 14648 9664 14700 9716
rect 4988 9596 5040 9648
rect 7656 9596 7708 9648
rect 11060 9596 11112 9648
rect 24768 9664 24820 9716
rect 26056 9707 26108 9716
rect 26056 9673 26065 9707
rect 26065 9673 26099 9707
rect 26099 9673 26108 9707
rect 26056 9664 26108 9673
rect 5632 9571 5684 9580
rect 5632 9537 5641 9571
rect 5641 9537 5675 9571
rect 5675 9537 5684 9571
rect 5632 9528 5684 9537
rect 6828 9528 6880 9580
rect 8300 9528 8352 9580
rect 9588 9528 9640 9580
rect 5540 9503 5592 9512
rect 5540 9469 5549 9503
rect 5549 9469 5583 9503
rect 5583 9469 5592 9503
rect 5540 9460 5592 9469
rect 9496 9460 9548 9512
rect 12072 9571 12124 9580
rect 12072 9537 12081 9571
rect 12081 9537 12115 9571
rect 12115 9537 12124 9571
rect 12072 9528 12124 9537
rect 16396 9528 16448 9580
rect 16580 9528 16632 9580
rect 17592 9528 17644 9580
rect 21916 9528 21968 9580
rect 22836 9528 22888 9580
rect 24860 9596 24912 9648
rect 25044 9596 25096 9648
rect 28172 9664 28224 9716
rect 27896 9596 27948 9648
rect 29000 9596 29052 9648
rect 31024 9664 31076 9716
rect 29828 9571 29880 9580
rect 29828 9537 29837 9571
rect 29837 9537 29871 9571
rect 29871 9537 29880 9571
rect 29828 9528 29880 9537
rect 11980 9503 12032 9512
rect 11980 9469 11989 9503
rect 11989 9469 12023 9503
rect 12023 9469 12032 9503
rect 11980 9460 12032 9469
rect 12440 9503 12492 9512
rect 12440 9469 12449 9503
rect 12449 9469 12483 9503
rect 12483 9469 12492 9503
rect 12440 9460 12492 9469
rect 14464 9460 14516 9512
rect 15384 9503 15436 9512
rect 15384 9469 15393 9503
rect 15393 9469 15427 9503
rect 15427 9469 15436 9503
rect 15384 9460 15436 9469
rect 18144 9460 18196 9512
rect 29368 9503 29420 9512
rect 29368 9469 29377 9503
rect 29377 9469 29411 9503
rect 29411 9469 29420 9503
rect 29368 9460 29420 9469
rect 14832 9367 14884 9376
rect 14832 9333 14841 9367
rect 14841 9333 14875 9367
rect 14875 9333 14884 9367
rect 14832 9324 14884 9333
rect 23848 9324 23900 9376
rect 4664 9222 4716 9274
rect 4728 9222 4780 9274
rect 4792 9222 4844 9274
rect 4856 9222 4908 9274
rect 4920 9222 4972 9274
rect 12092 9222 12144 9274
rect 12156 9222 12208 9274
rect 12220 9222 12272 9274
rect 12284 9222 12336 9274
rect 12348 9222 12400 9274
rect 19520 9222 19572 9274
rect 19584 9222 19636 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 26948 9222 27000 9274
rect 27012 9222 27064 9274
rect 27076 9222 27128 9274
rect 27140 9222 27192 9274
rect 27204 9222 27256 9274
rect 9680 9163 9732 9172
rect 9680 9129 9689 9163
rect 9689 9129 9723 9163
rect 9723 9129 9732 9163
rect 9680 9120 9732 9129
rect 14464 9163 14516 9172
rect 14464 9129 14473 9163
rect 14473 9129 14507 9163
rect 14507 9129 14516 9163
rect 14464 9120 14516 9129
rect 22836 9163 22888 9172
rect 22836 9129 22845 9163
rect 22845 9129 22879 9163
rect 22879 9129 22888 9163
rect 22836 9120 22888 9129
rect 25044 9120 25096 9172
rect 29828 9163 29880 9172
rect 29828 9129 29837 9163
rect 29837 9129 29871 9163
rect 29871 9129 29880 9163
rect 29828 9120 29880 9129
rect 8392 8984 8444 9036
rect 30012 9027 30064 9036
rect 30012 8993 30021 9027
rect 30021 8993 30055 9027
rect 30055 8993 30064 9027
rect 30012 8984 30064 8993
rect 5632 8916 5684 8968
rect 8300 8916 8352 8968
rect 9312 8959 9364 8968
rect 9312 8925 9321 8959
rect 9321 8925 9355 8959
rect 9355 8925 9364 8959
rect 9312 8916 9364 8925
rect 12256 8916 12308 8968
rect 14832 8916 14884 8968
rect 16212 8916 16264 8968
rect 19892 8959 19944 8968
rect 19892 8925 19901 8959
rect 19901 8925 19935 8959
rect 19935 8925 19944 8959
rect 19892 8916 19944 8925
rect 21456 8916 21508 8968
rect 23848 8916 23900 8968
rect 9496 8848 9548 8900
rect 12992 8891 13044 8900
rect 12992 8857 13001 8891
rect 13001 8857 13035 8891
rect 13035 8857 13044 8891
rect 12992 8848 13044 8857
rect 22284 8848 22336 8900
rect 24676 8916 24728 8968
rect 24768 8959 24820 8968
rect 24768 8925 24777 8959
rect 24777 8925 24811 8959
rect 24811 8925 24820 8959
rect 24768 8916 24820 8925
rect 27528 8916 27580 8968
rect 28908 8959 28960 8968
rect 28908 8925 28917 8959
rect 28917 8925 28951 8959
rect 28951 8925 28960 8959
rect 28908 8916 28960 8925
rect 30196 8916 30248 8968
rect 27712 8891 27764 8900
rect 27712 8857 27721 8891
rect 27721 8857 27755 8891
rect 27755 8857 27764 8891
rect 27712 8848 27764 8857
rect 27804 8848 27856 8900
rect 8760 8780 8812 8832
rect 13084 8780 13136 8832
rect 19984 8823 20036 8832
rect 19984 8789 19993 8823
rect 19993 8789 20027 8823
rect 20027 8789 20036 8823
rect 19984 8780 20036 8789
rect 27896 8823 27948 8832
rect 27896 8789 27905 8823
rect 27905 8789 27939 8823
rect 27939 8789 27948 8823
rect 27896 8780 27948 8789
rect 27988 8823 28040 8832
rect 27988 8789 27997 8823
rect 27997 8789 28031 8823
rect 28031 8789 28040 8823
rect 27988 8780 28040 8789
rect 8378 8678 8430 8730
rect 8442 8678 8494 8730
rect 8506 8678 8558 8730
rect 8570 8678 8622 8730
rect 8634 8678 8686 8730
rect 15806 8678 15858 8730
rect 15870 8678 15922 8730
rect 15934 8678 15986 8730
rect 15998 8678 16050 8730
rect 16062 8678 16114 8730
rect 23234 8678 23286 8730
rect 23298 8678 23350 8730
rect 23362 8678 23414 8730
rect 23426 8678 23478 8730
rect 23490 8678 23542 8730
rect 30662 8678 30714 8730
rect 30726 8678 30778 8730
rect 30790 8678 30842 8730
rect 30854 8678 30906 8730
rect 30918 8678 30970 8730
rect 8300 8619 8352 8628
rect 8300 8585 8309 8619
rect 8309 8585 8343 8619
rect 8343 8585 8352 8619
rect 8300 8576 8352 8585
rect 12900 8619 12952 8628
rect 12900 8585 12909 8619
rect 12909 8585 12943 8619
rect 12943 8585 12952 8619
rect 12900 8576 12952 8585
rect 19064 8576 19116 8628
rect 9220 8508 9272 8560
rect 19432 8576 19484 8628
rect 27436 8576 27488 8628
rect 29368 8576 29420 8628
rect 19984 8508 20036 8560
rect 5356 8440 5408 8492
rect 9312 8440 9364 8492
rect 11152 8483 11204 8492
rect 11152 8449 11161 8483
rect 11161 8449 11195 8483
rect 11195 8449 11204 8483
rect 11152 8440 11204 8449
rect 11244 8440 11296 8492
rect 12256 8483 12308 8492
rect 12256 8449 12265 8483
rect 12265 8449 12299 8483
rect 12299 8449 12308 8483
rect 12256 8440 12308 8449
rect 12992 8440 13044 8492
rect 13084 8483 13136 8492
rect 13084 8449 13093 8483
rect 13093 8449 13127 8483
rect 13127 8449 13136 8483
rect 13084 8440 13136 8449
rect 13452 8483 13504 8492
rect 13452 8449 13461 8483
rect 13461 8449 13495 8483
rect 13495 8449 13504 8483
rect 13452 8440 13504 8449
rect 13912 8483 13964 8492
rect 13912 8449 13921 8483
rect 13921 8449 13955 8483
rect 13955 8449 13964 8483
rect 13912 8440 13964 8449
rect 14464 8440 14516 8492
rect 19156 8440 19208 8492
rect 21456 8440 21508 8492
rect 24768 8508 24820 8560
rect 27528 8508 27580 8560
rect 22284 8440 22336 8492
rect 23848 8483 23900 8492
rect 23848 8449 23857 8483
rect 23857 8449 23891 8483
rect 23891 8449 23900 8483
rect 23848 8440 23900 8449
rect 5448 8372 5500 8424
rect 8300 8372 8352 8424
rect 6920 8304 6972 8356
rect 5724 8279 5776 8288
rect 5724 8245 5733 8279
rect 5733 8245 5767 8279
rect 5767 8245 5776 8279
rect 5724 8236 5776 8245
rect 11060 8279 11112 8288
rect 11060 8245 11069 8279
rect 11069 8245 11103 8279
rect 11103 8245 11112 8279
rect 11060 8236 11112 8245
rect 16672 8236 16724 8288
rect 17132 8415 17184 8424
rect 17132 8381 17141 8415
rect 17141 8381 17175 8415
rect 17175 8381 17184 8415
rect 17132 8372 17184 8381
rect 18972 8372 19024 8424
rect 27712 8440 27764 8492
rect 27896 8483 27948 8492
rect 27896 8449 27905 8483
rect 27905 8449 27939 8483
rect 27939 8449 27948 8483
rect 27896 8440 27948 8449
rect 27988 8483 28040 8492
rect 27988 8449 28033 8483
rect 28033 8449 28040 8483
rect 28540 8483 28592 8492
rect 27988 8440 28040 8449
rect 28540 8449 28549 8483
rect 28549 8449 28583 8483
rect 28583 8449 28592 8483
rect 28540 8440 28592 8449
rect 27804 8415 27856 8424
rect 27804 8381 27813 8415
rect 27813 8381 27847 8415
rect 27847 8381 27856 8415
rect 27804 8372 27856 8381
rect 18604 8236 18656 8288
rect 20812 8236 20864 8288
rect 22100 8279 22152 8288
rect 22100 8245 22109 8279
rect 22109 8245 22143 8279
rect 22143 8245 22152 8279
rect 22100 8236 22152 8245
rect 4664 8134 4716 8186
rect 4728 8134 4780 8186
rect 4792 8134 4844 8186
rect 4856 8134 4908 8186
rect 4920 8134 4972 8186
rect 12092 8134 12144 8186
rect 12156 8134 12208 8186
rect 12220 8134 12272 8186
rect 12284 8134 12336 8186
rect 12348 8134 12400 8186
rect 19520 8134 19572 8186
rect 19584 8134 19636 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 26948 8134 27000 8186
rect 27012 8134 27064 8186
rect 27076 8134 27128 8186
rect 27140 8134 27192 8186
rect 27204 8134 27256 8186
rect 12532 8075 12584 8084
rect 12532 8041 12541 8075
rect 12541 8041 12575 8075
rect 12575 8041 12584 8075
rect 12532 8032 12584 8041
rect 13452 8032 13504 8084
rect 16672 8032 16724 8084
rect 17132 8032 17184 8084
rect 19432 8032 19484 8084
rect 27528 8032 27580 8084
rect 5724 7896 5776 7948
rect 11060 7939 11112 7948
rect 11060 7905 11069 7939
rect 11069 7905 11103 7939
rect 11103 7905 11112 7939
rect 11060 7896 11112 7905
rect 18604 7939 18656 7948
rect 18604 7905 18613 7939
rect 18613 7905 18647 7939
rect 18647 7905 18656 7939
rect 18604 7896 18656 7905
rect 18972 7896 19024 7948
rect 20812 7939 20864 7948
rect 20812 7905 20821 7939
rect 20821 7905 20855 7939
rect 20855 7905 20864 7939
rect 20812 7896 20864 7905
rect 6092 7760 6144 7812
rect 6644 7692 6696 7744
rect 7104 7735 7156 7744
rect 7104 7701 7113 7735
rect 7113 7701 7147 7735
rect 7147 7701 7156 7735
rect 7840 7828 7892 7880
rect 9312 7871 9364 7880
rect 9312 7837 9321 7871
rect 9321 7837 9355 7871
rect 9355 7837 9364 7871
rect 9312 7828 9364 7837
rect 10784 7871 10836 7880
rect 10784 7837 10793 7871
rect 10793 7837 10827 7871
rect 10827 7837 10836 7871
rect 10784 7828 10836 7837
rect 14464 7828 14516 7880
rect 15200 7828 15252 7880
rect 18512 7828 18564 7880
rect 11704 7760 11756 7812
rect 7104 7692 7156 7701
rect 7748 7735 7800 7744
rect 7748 7701 7757 7735
rect 7757 7701 7791 7735
rect 7791 7701 7800 7735
rect 7748 7692 7800 7701
rect 8024 7692 8076 7744
rect 11060 7692 11112 7744
rect 13912 7760 13964 7812
rect 17408 7760 17460 7812
rect 17684 7692 17736 7744
rect 19616 7871 19668 7880
rect 19616 7837 19625 7871
rect 19625 7837 19659 7871
rect 19659 7837 19668 7871
rect 19616 7828 19668 7837
rect 19892 7828 19944 7880
rect 20444 7828 20496 7880
rect 23848 7828 23900 7880
rect 24308 7828 24360 7880
rect 28540 7871 28592 7880
rect 28540 7837 28549 7871
rect 28549 7837 28583 7871
rect 28583 7837 28592 7871
rect 28540 7828 28592 7837
rect 22100 7760 22152 7812
rect 22192 7692 22244 7744
rect 28448 7735 28500 7744
rect 28448 7701 28457 7735
rect 28457 7701 28491 7735
rect 28491 7701 28500 7735
rect 28448 7692 28500 7701
rect 8378 7590 8430 7642
rect 8442 7590 8494 7642
rect 8506 7590 8558 7642
rect 8570 7590 8622 7642
rect 8634 7590 8686 7642
rect 15806 7590 15858 7642
rect 15870 7590 15922 7642
rect 15934 7590 15986 7642
rect 15998 7590 16050 7642
rect 16062 7590 16114 7642
rect 23234 7590 23286 7642
rect 23298 7590 23350 7642
rect 23362 7590 23414 7642
rect 23426 7590 23478 7642
rect 23490 7590 23542 7642
rect 30662 7590 30714 7642
rect 30726 7590 30778 7642
rect 30790 7590 30842 7642
rect 30854 7590 30906 7642
rect 30918 7590 30970 7642
rect 6092 7488 6144 7540
rect 6644 7531 6696 7540
rect 6644 7497 6653 7531
rect 6653 7497 6687 7531
rect 6687 7497 6696 7531
rect 6644 7488 6696 7497
rect 10784 7531 10836 7540
rect 10784 7497 10793 7531
rect 10793 7497 10827 7531
rect 10827 7497 10836 7531
rect 10784 7488 10836 7497
rect 11704 7531 11756 7540
rect 11704 7497 11713 7531
rect 11713 7497 11747 7531
rect 11747 7497 11756 7531
rect 11704 7488 11756 7497
rect 5264 7352 5316 7404
rect 5632 7420 5684 7472
rect 8024 7463 8076 7472
rect 8024 7429 8033 7463
rect 8033 7429 8067 7463
rect 8067 7429 8076 7463
rect 8024 7420 8076 7429
rect 8760 7420 8812 7472
rect 5448 7395 5500 7404
rect 5448 7361 5457 7395
rect 5457 7361 5491 7395
rect 5491 7361 5500 7395
rect 5448 7352 5500 7361
rect 7104 7352 7156 7404
rect 7748 7395 7800 7404
rect 7748 7361 7757 7395
rect 7757 7361 7791 7395
rect 7791 7361 7800 7395
rect 7748 7352 7800 7361
rect 9312 7284 9364 7336
rect 11244 7352 11296 7404
rect 13360 7488 13412 7540
rect 16396 7488 16448 7540
rect 18512 7488 18564 7540
rect 28540 7488 28592 7540
rect 12440 7327 12492 7336
rect 12440 7293 12449 7327
rect 12449 7293 12483 7327
rect 12483 7293 12492 7327
rect 12440 7284 12492 7293
rect 16672 7352 16724 7404
rect 16764 7352 16816 7404
rect 21456 7395 21508 7404
rect 21456 7361 21465 7395
rect 21465 7361 21499 7395
rect 21499 7361 21508 7395
rect 21456 7352 21508 7361
rect 22284 7420 22336 7472
rect 28448 7420 28500 7472
rect 16212 7284 16264 7336
rect 17132 7327 17184 7336
rect 17132 7293 17141 7327
rect 17141 7293 17175 7327
rect 17175 7293 17184 7327
rect 17132 7284 17184 7293
rect 17500 7284 17552 7336
rect 19616 7284 19668 7336
rect 25964 7352 26016 7404
rect 27620 7395 27672 7404
rect 27620 7361 27629 7395
rect 27629 7361 27663 7395
rect 27663 7361 27672 7395
rect 27620 7352 27672 7361
rect 17684 7148 17736 7200
rect 21364 7191 21416 7200
rect 21364 7157 21373 7191
rect 21373 7157 21407 7191
rect 21407 7157 21416 7191
rect 21364 7148 21416 7157
rect 22652 7148 22704 7200
rect 22836 7148 22888 7200
rect 25320 7191 25372 7200
rect 25320 7157 25329 7191
rect 25329 7157 25363 7191
rect 25363 7157 25372 7191
rect 25320 7148 25372 7157
rect 4664 7046 4716 7098
rect 4728 7046 4780 7098
rect 4792 7046 4844 7098
rect 4856 7046 4908 7098
rect 4920 7046 4972 7098
rect 12092 7046 12144 7098
rect 12156 7046 12208 7098
rect 12220 7046 12272 7098
rect 12284 7046 12336 7098
rect 12348 7046 12400 7098
rect 19520 7046 19572 7098
rect 19584 7046 19636 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 26948 7046 27000 7098
rect 27012 7046 27064 7098
rect 27076 7046 27128 7098
rect 27140 7046 27192 7098
rect 27204 7046 27256 7098
rect 6920 6987 6972 6996
rect 6920 6953 6941 6987
rect 6941 6953 6972 6987
rect 6920 6944 6972 6953
rect 25964 6987 26016 6996
rect 25964 6953 25973 6987
rect 25973 6953 26007 6987
rect 26007 6953 26016 6987
rect 25964 6944 26016 6953
rect 5356 6808 5408 6860
rect 9956 6808 10008 6860
rect 7196 6783 7248 6792
rect 7196 6749 7205 6783
rect 7205 6749 7239 6783
rect 7239 6749 7248 6783
rect 7196 6740 7248 6749
rect 8760 6740 8812 6792
rect 5908 6672 5960 6724
rect 9404 6715 9456 6724
rect 9404 6681 9413 6715
rect 9413 6681 9447 6715
rect 9447 6681 9456 6715
rect 9404 6672 9456 6681
rect 10048 6672 10100 6724
rect 8300 6604 8352 6656
rect 11060 6604 11112 6656
rect 13544 6604 13596 6656
rect 14648 6783 14700 6792
rect 14648 6749 14657 6783
rect 14657 6749 14691 6783
rect 14691 6749 14700 6783
rect 14648 6740 14700 6749
rect 17132 6808 17184 6860
rect 17408 6808 17460 6860
rect 20444 6851 20496 6860
rect 20444 6817 20453 6851
rect 20453 6817 20487 6851
rect 20487 6817 20496 6851
rect 20444 6808 20496 6817
rect 22192 6808 22244 6860
rect 27712 6808 27764 6860
rect 30012 6808 30064 6860
rect 16672 6740 16724 6792
rect 17500 6783 17552 6792
rect 17500 6749 17509 6783
rect 17509 6749 17543 6783
rect 17543 6749 17552 6783
rect 17500 6740 17552 6749
rect 17684 6783 17736 6792
rect 17684 6749 17693 6783
rect 17693 6749 17727 6783
rect 17727 6749 17736 6783
rect 17684 6740 17736 6749
rect 24584 6783 24636 6792
rect 24584 6749 24593 6783
rect 24593 6749 24627 6783
rect 24627 6749 24636 6783
rect 24584 6740 24636 6749
rect 25320 6740 25372 6792
rect 25964 6740 26016 6792
rect 28816 6783 28868 6792
rect 28816 6749 28825 6783
rect 28825 6749 28859 6783
rect 28859 6749 28868 6783
rect 28816 6740 28868 6749
rect 28908 6783 28960 6792
rect 28908 6749 28917 6783
rect 28917 6749 28951 6783
rect 28951 6749 28960 6783
rect 28908 6740 28960 6749
rect 16488 6672 16540 6724
rect 21364 6672 21416 6724
rect 27896 6672 27948 6724
rect 14372 6604 14424 6656
rect 16856 6604 16908 6656
rect 22376 6604 22428 6656
rect 27344 6604 27396 6656
rect 28448 6647 28500 6656
rect 28448 6613 28457 6647
rect 28457 6613 28491 6647
rect 28491 6613 28500 6647
rect 28448 6604 28500 6613
rect 8378 6502 8430 6554
rect 8442 6502 8494 6554
rect 8506 6502 8558 6554
rect 8570 6502 8622 6554
rect 8634 6502 8686 6554
rect 15806 6502 15858 6554
rect 15870 6502 15922 6554
rect 15934 6502 15986 6554
rect 15998 6502 16050 6554
rect 16062 6502 16114 6554
rect 23234 6502 23286 6554
rect 23298 6502 23350 6554
rect 23362 6502 23414 6554
rect 23426 6502 23478 6554
rect 23490 6502 23542 6554
rect 30662 6502 30714 6554
rect 30726 6502 30778 6554
rect 30790 6502 30842 6554
rect 30854 6502 30906 6554
rect 30918 6502 30970 6554
rect 5908 6400 5960 6452
rect 7196 6400 7248 6452
rect 9404 6400 9456 6452
rect 5080 6332 5132 6384
rect 9956 6400 10008 6452
rect 10048 6443 10100 6452
rect 10048 6409 10057 6443
rect 10057 6409 10091 6443
rect 10091 6409 10100 6443
rect 10048 6400 10100 6409
rect 12624 6400 12676 6452
rect 24584 6400 24636 6452
rect 27620 6400 27672 6452
rect 28356 6400 28408 6452
rect 11980 6332 12032 6384
rect 22744 6332 22796 6384
rect 28908 6332 28960 6384
rect 5264 6307 5316 6316
rect 5264 6273 5273 6307
rect 5273 6273 5307 6307
rect 5307 6273 5316 6307
rect 5264 6264 5316 6273
rect 5448 6307 5500 6316
rect 5448 6273 5457 6307
rect 5457 6273 5491 6307
rect 5491 6273 5500 6307
rect 5448 6264 5500 6273
rect 8300 6307 8352 6316
rect 8300 6273 8309 6307
rect 8309 6273 8343 6307
rect 8343 6273 8352 6307
rect 8300 6264 8352 6273
rect 9404 6307 9456 6316
rect 9404 6273 9413 6307
rect 9413 6273 9447 6307
rect 9447 6273 9456 6307
rect 9404 6264 9456 6273
rect 9588 6264 9640 6316
rect 8760 6196 8812 6248
rect 13544 6307 13596 6316
rect 13544 6273 13553 6307
rect 13553 6273 13587 6307
rect 13587 6273 13596 6307
rect 13544 6264 13596 6273
rect 22376 6307 22428 6316
rect 22376 6273 22385 6307
rect 22385 6273 22419 6307
rect 22419 6273 22428 6307
rect 22376 6264 22428 6273
rect 24308 6307 24360 6316
rect 24308 6273 24317 6307
rect 24317 6273 24351 6307
rect 24351 6273 24360 6307
rect 24308 6264 24360 6273
rect 21456 6196 21508 6248
rect 25964 6264 26016 6316
rect 29092 6264 29144 6316
rect 21732 6060 21784 6112
rect 28816 6196 28868 6248
rect 28448 6128 28500 6180
rect 27436 6060 27488 6112
rect 29828 6060 29880 6112
rect 4664 5958 4716 6010
rect 4728 5958 4780 6010
rect 4792 5958 4844 6010
rect 4856 5958 4908 6010
rect 4920 5958 4972 6010
rect 12092 5958 12144 6010
rect 12156 5958 12208 6010
rect 12220 5958 12272 6010
rect 12284 5958 12336 6010
rect 12348 5958 12400 6010
rect 19520 5958 19572 6010
rect 19584 5958 19636 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 26948 5958 27000 6010
rect 27012 5958 27064 6010
rect 27076 5958 27128 6010
rect 27140 5958 27192 6010
rect 27204 5958 27256 6010
rect 14648 5856 14700 5908
rect 28908 5856 28960 5908
rect 29092 5899 29144 5908
rect 29092 5865 29101 5899
rect 29101 5865 29135 5899
rect 29135 5865 29144 5899
rect 29092 5856 29144 5865
rect 9588 5720 9640 5772
rect 9404 5652 9456 5704
rect 11980 5720 12032 5772
rect 16856 5720 16908 5772
rect 19708 5763 19760 5772
rect 19708 5729 19717 5763
rect 19717 5729 19751 5763
rect 19751 5729 19760 5763
rect 19708 5720 19760 5729
rect 19984 5763 20036 5772
rect 19984 5729 19993 5763
rect 19993 5729 20027 5763
rect 20027 5729 20036 5763
rect 19984 5720 20036 5729
rect 20444 5720 20496 5772
rect 20812 5720 20864 5772
rect 21456 5763 21508 5772
rect 21456 5729 21465 5763
rect 21465 5729 21499 5763
rect 21499 5729 21508 5763
rect 21456 5720 21508 5729
rect 21732 5763 21784 5772
rect 21732 5729 21741 5763
rect 21741 5729 21775 5763
rect 21775 5729 21784 5763
rect 21732 5720 21784 5729
rect 24308 5720 24360 5772
rect 12440 5652 12492 5704
rect 19432 5584 19484 5636
rect 17960 5516 18012 5568
rect 22836 5652 22888 5704
rect 25964 5652 26016 5704
rect 27896 5788 27948 5840
rect 28724 5720 28776 5772
rect 31024 5720 31076 5772
rect 27344 5652 27396 5704
rect 27712 5652 27764 5704
rect 27896 5584 27948 5636
rect 28356 5695 28408 5704
rect 28356 5661 28365 5695
rect 28365 5661 28399 5695
rect 28399 5661 28408 5695
rect 28356 5652 28408 5661
rect 29828 5695 29880 5704
rect 29828 5661 29837 5695
rect 29837 5661 29871 5695
rect 29871 5661 29880 5695
rect 29828 5652 29880 5661
rect 27436 5516 27488 5568
rect 8378 5414 8430 5466
rect 8442 5414 8494 5466
rect 8506 5414 8558 5466
rect 8570 5414 8622 5466
rect 8634 5414 8686 5466
rect 15806 5414 15858 5466
rect 15870 5414 15922 5466
rect 15934 5414 15986 5466
rect 15998 5414 16050 5466
rect 16062 5414 16114 5466
rect 23234 5414 23286 5466
rect 23298 5414 23350 5466
rect 23362 5414 23414 5466
rect 23426 5414 23478 5466
rect 23490 5414 23542 5466
rect 30662 5414 30714 5466
rect 30726 5414 30778 5466
rect 30790 5414 30842 5466
rect 30854 5414 30906 5466
rect 30918 5414 30970 5466
rect 19708 5312 19760 5364
rect 27896 5312 27948 5364
rect 14556 5176 14608 5228
rect 17224 5219 17276 5228
rect 17224 5185 17258 5219
rect 17258 5185 17276 5219
rect 17224 5176 17276 5185
rect 28356 5244 28408 5296
rect 18604 5176 18656 5228
rect 27436 5219 27488 5228
rect 27436 5185 27445 5219
rect 27445 5185 27479 5219
rect 27479 5185 27488 5219
rect 27436 5176 27488 5185
rect 27712 5176 27764 5228
rect 28724 5219 28776 5228
rect 28724 5185 28733 5219
rect 28733 5185 28767 5219
rect 28767 5185 28776 5219
rect 28724 5176 28776 5185
rect 28816 5176 28868 5228
rect 14372 5151 14424 5160
rect 14372 5117 14381 5151
rect 14381 5117 14415 5151
rect 14415 5117 14424 5151
rect 14372 5108 14424 5117
rect 28448 5040 28500 5092
rect 14004 4972 14056 5024
rect 28724 5015 28776 5024
rect 28724 4981 28733 5015
rect 28733 4981 28767 5015
rect 28767 4981 28776 5015
rect 28724 4972 28776 4981
rect 4664 4870 4716 4922
rect 4728 4870 4780 4922
rect 4792 4870 4844 4922
rect 4856 4870 4908 4922
rect 4920 4870 4972 4922
rect 12092 4870 12144 4922
rect 12156 4870 12208 4922
rect 12220 4870 12272 4922
rect 12284 4870 12336 4922
rect 12348 4870 12400 4922
rect 19520 4870 19572 4922
rect 19584 4870 19636 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 26948 4870 27000 4922
rect 27012 4870 27064 4922
rect 27076 4870 27128 4922
rect 27140 4870 27192 4922
rect 27204 4870 27256 4922
rect 17224 4811 17276 4820
rect 17224 4777 17233 4811
rect 17233 4777 17267 4811
rect 17267 4777 17276 4811
rect 17224 4768 17276 4777
rect 19432 4811 19484 4820
rect 19432 4777 19441 4811
rect 19441 4777 19475 4811
rect 19475 4777 19484 4811
rect 19432 4768 19484 4777
rect 14372 4700 14424 4752
rect 14648 4675 14700 4684
rect 14648 4641 14657 4675
rect 14657 4641 14691 4675
rect 14691 4641 14700 4675
rect 14648 4632 14700 4641
rect 14556 4607 14608 4616
rect 14556 4573 14565 4607
rect 14565 4573 14599 4607
rect 14599 4573 14608 4607
rect 14556 4564 14608 4573
rect 20812 4675 20864 4684
rect 20812 4641 20821 4675
rect 20821 4641 20855 4675
rect 20855 4641 20864 4675
rect 20812 4632 20864 4641
rect 17960 4564 18012 4616
rect 19984 4564 20036 4616
rect 8378 4326 8430 4378
rect 8442 4326 8494 4378
rect 8506 4326 8558 4378
rect 8570 4326 8622 4378
rect 8634 4326 8686 4378
rect 15806 4326 15858 4378
rect 15870 4326 15922 4378
rect 15934 4326 15986 4378
rect 15998 4326 16050 4378
rect 16062 4326 16114 4378
rect 23234 4326 23286 4378
rect 23298 4326 23350 4378
rect 23362 4326 23414 4378
rect 23426 4326 23478 4378
rect 23490 4326 23542 4378
rect 30662 4326 30714 4378
rect 30726 4326 30778 4378
rect 30790 4326 30842 4378
rect 30854 4326 30906 4378
rect 30918 4326 30970 4378
rect 14648 4224 14700 4276
rect 14372 4156 14424 4208
rect 14004 4131 14056 4140
rect 14004 4097 14038 4131
rect 14038 4097 14056 4131
rect 14004 4088 14056 4097
rect 4664 3782 4716 3834
rect 4728 3782 4780 3834
rect 4792 3782 4844 3834
rect 4856 3782 4908 3834
rect 4920 3782 4972 3834
rect 12092 3782 12144 3834
rect 12156 3782 12208 3834
rect 12220 3782 12272 3834
rect 12284 3782 12336 3834
rect 12348 3782 12400 3834
rect 19520 3782 19572 3834
rect 19584 3782 19636 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 26948 3782 27000 3834
rect 27012 3782 27064 3834
rect 27076 3782 27128 3834
rect 27140 3782 27192 3834
rect 27204 3782 27256 3834
rect 8378 3238 8430 3290
rect 8442 3238 8494 3290
rect 8506 3238 8558 3290
rect 8570 3238 8622 3290
rect 8634 3238 8686 3290
rect 15806 3238 15858 3290
rect 15870 3238 15922 3290
rect 15934 3238 15986 3290
rect 15998 3238 16050 3290
rect 16062 3238 16114 3290
rect 23234 3238 23286 3290
rect 23298 3238 23350 3290
rect 23362 3238 23414 3290
rect 23426 3238 23478 3290
rect 23490 3238 23542 3290
rect 30662 3238 30714 3290
rect 30726 3238 30778 3290
rect 30790 3238 30842 3290
rect 30854 3238 30906 3290
rect 30918 3238 30970 3290
rect 4664 2694 4716 2746
rect 4728 2694 4780 2746
rect 4792 2694 4844 2746
rect 4856 2694 4908 2746
rect 4920 2694 4972 2746
rect 12092 2694 12144 2746
rect 12156 2694 12208 2746
rect 12220 2694 12272 2746
rect 12284 2694 12336 2746
rect 12348 2694 12400 2746
rect 19520 2694 19572 2746
rect 19584 2694 19636 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 26948 2694 27000 2746
rect 27012 2694 27064 2746
rect 27076 2694 27128 2746
rect 27140 2694 27192 2746
rect 27204 2694 27256 2746
rect 28724 2388 28776 2440
rect 31024 2320 31076 2372
rect 8378 2150 8430 2202
rect 8442 2150 8494 2202
rect 8506 2150 8558 2202
rect 8570 2150 8622 2202
rect 8634 2150 8686 2202
rect 15806 2150 15858 2202
rect 15870 2150 15922 2202
rect 15934 2150 15986 2202
rect 15998 2150 16050 2202
rect 16062 2150 16114 2202
rect 23234 2150 23286 2202
rect 23298 2150 23350 2202
rect 23362 2150 23414 2202
rect 23426 2150 23478 2202
rect 23490 2150 23542 2202
rect 30662 2150 30714 2202
rect 30726 2150 30778 2202
rect 30790 2150 30842 2202
rect 30854 2150 30906 2202
rect 30918 2150 30970 2202
<< metal2 >>
rect 2134 31200 2190 32000
rect 6090 31200 6146 32000
rect 10046 31362 10102 32000
rect 10046 31334 10272 31362
rect 10046 31200 10102 31334
rect 2148 28762 2176 31200
rect 6104 29238 6132 31200
rect 8378 29404 8686 29413
rect 8378 29402 8384 29404
rect 8440 29402 8464 29404
rect 8520 29402 8544 29404
rect 8600 29402 8624 29404
rect 8680 29402 8686 29404
rect 8440 29350 8442 29402
rect 8622 29350 8624 29402
rect 8378 29348 8384 29350
rect 8440 29348 8464 29350
rect 8520 29348 8544 29350
rect 8600 29348 8624 29350
rect 8680 29348 8686 29350
rect 8378 29339 8686 29348
rect 6092 29232 6144 29238
rect 6092 29174 6144 29180
rect 10244 29170 10272 31334
rect 14002 31200 14058 32000
rect 17958 31362 18014 32000
rect 21914 31362 21970 32000
rect 25870 31362 25926 32000
rect 17958 31334 18184 31362
rect 17958 31200 18014 31334
rect 14016 29170 14044 31200
rect 15806 29404 16114 29413
rect 15806 29402 15812 29404
rect 15868 29402 15892 29404
rect 15948 29402 15972 29404
rect 16028 29402 16052 29404
rect 16108 29402 16114 29404
rect 15868 29350 15870 29402
rect 16050 29350 16052 29402
rect 15806 29348 15812 29350
rect 15868 29348 15892 29350
rect 15948 29348 15972 29350
rect 16028 29348 16052 29350
rect 16108 29348 16114 29350
rect 15806 29339 16114 29348
rect 18156 29238 18184 31334
rect 21914 31334 22048 31362
rect 21914 31200 21970 31334
rect 15384 29232 15436 29238
rect 15384 29174 15436 29180
rect 18144 29232 18196 29238
rect 18144 29174 18196 29180
rect 3240 29164 3292 29170
rect 3240 29106 3292 29112
rect 10232 29164 10284 29170
rect 10232 29106 10284 29112
rect 14004 29164 14056 29170
rect 14004 29106 14056 29112
rect 3056 29096 3108 29102
rect 3056 29038 3108 29044
rect 2136 28756 2188 28762
rect 2136 28698 2188 28704
rect 3068 28490 3096 29038
rect 3148 28688 3200 28694
rect 3148 28630 3200 28636
rect 3056 28484 3108 28490
rect 3056 28426 3108 28432
rect 2872 28144 2924 28150
rect 2872 28086 2924 28092
rect 2320 27328 2372 27334
rect 2320 27270 2372 27276
rect 2332 26450 2360 27270
rect 2884 26994 2912 28086
rect 2964 28076 3016 28082
rect 2964 28018 3016 28024
rect 2976 27674 3004 28018
rect 2964 27668 3016 27674
rect 2964 27610 3016 27616
rect 2872 26988 2924 26994
rect 2872 26930 2924 26936
rect 2320 26444 2372 26450
rect 2320 26386 2372 26392
rect 2884 26042 2912 26930
rect 3068 26314 3096 28426
rect 3160 27470 3188 28630
rect 3252 28558 3280 29106
rect 14464 29096 14516 29102
rect 14464 29038 14516 29044
rect 4528 29028 4580 29034
rect 4528 28970 4580 28976
rect 7196 29028 7248 29034
rect 7196 28970 7248 28976
rect 3516 28756 3568 28762
rect 3516 28698 3568 28704
rect 3240 28552 3292 28558
rect 3240 28494 3292 28500
rect 3252 27538 3280 28494
rect 3240 27532 3292 27538
rect 3240 27474 3292 27480
rect 3148 27464 3200 27470
rect 3148 27406 3200 27412
rect 3424 27328 3476 27334
rect 3424 27270 3476 27276
rect 3332 27124 3384 27130
rect 3332 27066 3384 27072
rect 3344 26518 3372 27066
rect 3436 26994 3464 27270
rect 3424 26988 3476 26994
rect 3424 26930 3476 26936
rect 3332 26512 3384 26518
rect 3332 26454 3384 26460
rect 3436 26382 3464 26930
rect 3424 26376 3476 26382
rect 3424 26318 3476 26324
rect 3056 26308 3108 26314
rect 3056 26250 3108 26256
rect 2872 26036 2924 26042
rect 2924 25996 3096 26024
rect 2872 25978 2924 25984
rect 2872 25152 2924 25158
rect 2872 25094 2924 25100
rect 2320 24200 2372 24206
rect 2320 24142 2372 24148
rect 2332 23798 2360 24142
rect 2884 23798 2912 25094
rect 3068 24818 3096 25996
rect 3148 25288 3200 25294
rect 3148 25230 3200 25236
rect 3240 25288 3292 25294
rect 3240 25230 3292 25236
rect 2964 24812 3016 24818
rect 2964 24754 3016 24760
rect 3056 24812 3108 24818
rect 3056 24754 3108 24760
rect 2976 24410 3004 24754
rect 2964 24404 3016 24410
rect 2964 24346 3016 24352
rect 3160 24342 3188 25230
rect 3252 24410 3280 25230
rect 3528 24818 3556 28698
rect 3884 28552 3936 28558
rect 3884 28494 3936 28500
rect 3896 27878 3924 28494
rect 4540 28150 4568 28970
rect 4664 28860 4972 28869
rect 4664 28858 4670 28860
rect 4726 28858 4750 28860
rect 4806 28858 4830 28860
rect 4886 28858 4910 28860
rect 4966 28858 4972 28860
rect 4726 28806 4728 28858
rect 4908 28806 4910 28858
rect 4664 28804 4670 28806
rect 4726 28804 4750 28806
rect 4806 28804 4830 28806
rect 4886 28804 4910 28806
rect 4966 28804 4972 28806
rect 4664 28795 4972 28804
rect 7208 28558 7236 28970
rect 12092 28860 12400 28869
rect 12092 28858 12098 28860
rect 12154 28858 12178 28860
rect 12234 28858 12258 28860
rect 12314 28858 12338 28860
rect 12394 28858 12400 28860
rect 12154 28806 12156 28858
rect 12336 28806 12338 28858
rect 12092 28804 12098 28806
rect 12154 28804 12178 28806
rect 12234 28804 12258 28806
rect 12314 28804 12338 28806
rect 12394 28804 12400 28806
rect 12092 28795 12400 28804
rect 7196 28552 7248 28558
rect 7196 28494 7248 28500
rect 8760 28552 8812 28558
rect 8760 28494 8812 28500
rect 10324 28552 10376 28558
rect 10324 28494 10376 28500
rect 11060 28552 11112 28558
rect 11060 28494 11112 28500
rect 11704 28552 11756 28558
rect 11704 28494 11756 28500
rect 12716 28552 12768 28558
rect 12716 28494 12768 28500
rect 13728 28552 13780 28558
rect 13728 28494 13780 28500
rect 7012 28416 7064 28422
rect 7012 28358 7064 28364
rect 4528 28144 4580 28150
rect 4528 28086 4580 28092
rect 6920 28076 6972 28082
rect 6920 28018 6972 28024
rect 3976 28008 4028 28014
rect 3976 27950 4028 27956
rect 3884 27872 3936 27878
rect 3884 27814 3936 27820
rect 3896 27690 3924 27814
rect 3804 27674 3924 27690
rect 3804 27668 3936 27674
rect 3804 27662 3884 27668
rect 3608 27396 3660 27402
rect 3608 27338 3660 27344
rect 3620 26586 3648 27338
rect 3608 26580 3660 26586
rect 3608 26522 3660 26528
rect 3804 26382 3832 27662
rect 3884 27610 3936 27616
rect 3988 27538 4016 27950
rect 5908 27872 5960 27878
rect 5908 27814 5960 27820
rect 4664 27772 4972 27781
rect 4664 27770 4670 27772
rect 4726 27770 4750 27772
rect 4806 27770 4830 27772
rect 4886 27770 4910 27772
rect 4966 27770 4972 27772
rect 4726 27718 4728 27770
rect 4908 27718 4910 27770
rect 4664 27716 4670 27718
rect 4726 27716 4750 27718
rect 4806 27716 4830 27718
rect 4886 27716 4910 27718
rect 4966 27716 4972 27718
rect 4664 27707 4972 27716
rect 5816 27600 5868 27606
rect 5816 27542 5868 27548
rect 3884 27532 3936 27538
rect 3884 27474 3936 27480
rect 3976 27532 4028 27538
rect 3976 27474 4028 27480
rect 3896 26586 3924 27474
rect 5828 27130 5856 27542
rect 5920 27470 5948 27814
rect 5908 27464 5960 27470
rect 5908 27406 5960 27412
rect 6644 27464 6696 27470
rect 6644 27406 6696 27412
rect 6656 27130 6684 27406
rect 5816 27124 5868 27130
rect 5816 27066 5868 27072
rect 6644 27124 6696 27130
rect 6644 27066 6696 27072
rect 4988 26988 5040 26994
rect 4988 26930 5040 26936
rect 4252 26852 4304 26858
rect 4252 26794 4304 26800
rect 3884 26580 3936 26586
rect 3884 26522 3936 26528
rect 4264 26382 4292 26794
rect 4664 26684 4972 26693
rect 4664 26682 4670 26684
rect 4726 26682 4750 26684
rect 4806 26682 4830 26684
rect 4886 26682 4910 26684
rect 4966 26682 4972 26684
rect 4726 26630 4728 26682
rect 4908 26630 4910 26682
rect 4664 26628 4670 26630
rect 4726 26628 4750 26630
rect 4806 26628 4830 26630
rect 4886 26628 4910 26630
rect 4966 26628 4972 26630
rect 4664 26619 4972 26628
rect 3792 26376 3844 26382
rect 3792 26318 3844 26324
rect 4252 26376 4304 26382
rect 4252 26318 4304 26324
rect 3976 26308 4028 26314
rect 3976 26250 4028 26256
rect 3988 26194 4016 26250
rect 4160 26240 4212 26246
rect 3988 26166 4108 26194
rect 4160 26182 4212 26188
rect 4080 25294 4108 26166
rect 4172 25294 4200 26182
rect 4344 25900 4396 25906
rect 4344 25842 4396 25848
rect 4068 25288 4120 25294
rect 4068 25230 4120 25236
rect 4160 25288 4212 25294
rect 4160 25230 4212 25236
rect 3516 24812 3568 24818
rect 3516 24754 3568 24760
rect 3424 24608 3476 24614
rect 3424 24550 3476 24556
rect 3240 24404 3292 24410
rect 3240 24346 3292 24352
rect 3148 24336 3200 24342
rect 3148 24278 3200 24284
rect 3436 24274 3464 24550
rect 3976 24404 4028 24410
rect 3976 24346 4028 24352
rect 3424 24268 3476 24274
rect 3424 24210 3476 24216
rect 3988 23866 4016 24346
rect 3976 23860 4028 23866
rect 3976 23802 4028 23808
rect 4080 23798 4108 25230
rect 4172 24206 4200 25230
rect 4356 24614 4384 25842
rect 4664 25596 4972 25605
rect 4664 25594 4670 25596
rect 4726 25594 4750 25596
rect 4806 25594 4830 25596
rect 4886 25594 4910 25596
rect 4966 25594 4972 25596
rect 4726 25542 4728 25594
rect 4908 25542 4910 25594
rect 4664 25540 4670 25542
rect 4726 25540 4750 25542
rect 4806 25540 4830 25542
rect 4886 25540 4910 25542
rect 4966 25540 4972 25542
rect 4664 25531 4972 25540
rect 5000 25498 5028 26930
rect 6736 26784 6788 26790
rect 6736 26726 6788 26732
rect 6748 25974 6776 26726
rect 6932 26382 6960 28018
rect 7024 27674 7052 28358
rect 7012 27668 7064 27674
rect 7012 27610 7064 27616
rect 6920 26376 6972 26382
rect 6920 26318 6972 26324
rect 6736 25968 6788 25974
rect 6736 25910 6788 25916
rect 6552 25832 6604 25838
rect 6552 25774 6604 25780
rect 4988 25492 5040 25498
rect 4988 25434 5040 25440
rect 5264 25220 5316 25226
rect 5264 25162 5316 25168
rect 4344 24608 4396 24614
rect 4344 24550 4396 24556
rect 4160 24200 4212 24206
rect 4160 24142 4212 24148
rect 4172 24070 4200 24142
rect 4160 24064 4212 24070
rect 4160 24006 4212 24012
rect 2320 23792 2372 23798
rect 2320 23734 2372 23740
rect 2872 23792 2924 23798
rect 2872 23734 2924 23740
rect 4068 23792 4120 23798
rect 4068 23734 4120 23740
rect 2332 23186 2360 23734
rect 2688 23724 2740 23730
rect 2688 23666 2740 23672
rect 2320 23180 2372 23186
rect 2320 23122 2372 23128
rect 1860 23112 1912 23118
rect 2332 23066 2360 23122
rect 1860 23054 1912 23060
rect 1872 22710 1900 23054
rect 2240 23038 2360 23066
rect 1860 22704 1912 22710
rect 1860 22646 1912 22652
rect 2240 22642 2268 23038
rect 2320 22976 2372 22982
rect 2320 22918 2372 22924
rect 2228 22636 2280 22642
rect 2228 22578 2280 22584
rect 2332 21962 2360 22918
rect 2700 22574 2728 23666
rect 4252 23316 4304 23322
rect 4252 23258 4304 23264
rect 3700 23112 3752 23118
rect 3700 23054 3752 23060
rect 3332 22704 3384 22710
rect 3332 22646 3384 22652
rect 2964 22636 3016 22642
rect 2964 22578 3016 22584
rect 2688 22568 2740 22574
rect 2688 22510 2740 22516
rect 2700 22030 2728 22510
rect 2688 22024 2740 22030
rect 2688 21966 2740 21972
rect 2320 21956 2372 21962
rect 2320 21898 2372 21904
rect 2700 21486 2728 21966
rect 2688 21480 2740 21486
rect 2688 21422 2740 21428
rect 2700 21010 2728 21422
rect 2976 21146 3004 22578
rect 3056 22432 3108 22438
rect 3056 22374 3108 22380
rect 2964 21140 3016 21146
rect 2964 21082 3016 21088
rect 2688 21004 2740 21010
rect 2688 20946 2740 20952
rect 3068 20942 3096 22374
rect 3344 21146 3372 22646
rect 3712 22506 3740 23054
rect 4160 22976 4212 22982
rect 4160 22918 4212 22924
rect 4068 22772 4120 22778
rect 4068 22714 4120 22720
rect 3700 22500 3752 22506
rect 3700 22442 3752 22448
rect 3712 22234 3740 22442
rect 3700 22228 3752 22234
rect 3700 22170 3752 22176
rect 4080 22094 4108 22714
rect 4172 22438 4200 22918
rect 4264 22642 4292 23258
rect 4252 22636 4304 22642
rect 4252 22578 4304 22584
rect 4160 22432 4212 22438
rect 4160 22374 4212 22380
rect 4080 22066 4200 22094
rect 4172 21962 4200 22066
rect 4160 21956 4212 21962
rect 4160 21898 4212 21904
rect 3332 21140 3384 21146
rect 3332 21082 3384 21088
rect 3056 20936 3108 20942
rect 3056 20878 3108 20884
rect 3976 20936 4028 20942
rect 3976 20878 4028 20884
rect 3988 20398 4016 20878
rect 4172 20806 4200 21898
rect 4356 21622 4384 24550
rect 4664 24508 4972 24517
rect 4664 24506 4670 24508
rect 4726 24506 4750 24508
rect 4806 24506 4830 24508
rect 4886 24506 4910 24508
rect 4966 24506 4972 24508
rect 4726 24454 4728 24506
rect 4908 24454 4910 24506
rect 4664 24452 4670 24454
rect 4726 24452 4750 24454
rect 4806 24452 4830 24454
rect 4886 24452 4910 24454
rect 4966 24452 4972 24454
rect 4664 24443 4972 24452
rect 5172 24336 5224 24342
rect 5172 24278 5224 24284
rect 5184 23730 5212 24278
rect 5276 23866 5304 25162
rect 6564 24954 6592 25774
rect 6828 25288 6880 25294
rect 6828 25230 6880 25236
rect 6552 24948 6604 24954
rect 6552 24890 6604 24896
rect 6736 24812 6788 24818
rect 6736 24754 6788 24760
rect 5264 23860 5316 23866
rect 5264 23802 5316 23808
rect 4988 23724 5040 23730
rect 4988 23666 5040 23672
rect 5172 23724 5224 23730
rect 5172 23666 5224 23672
rect 4528 23520 4580 23526
rect 4528 23462 4580 23468
rect 4540 23118 4568 23462
rect 4664 23420 4972 23429
rect 4664 23418 4670 23420
rect 4726 23418 4750 23420
rect 4806 23418 4830 23420
rect 4886 23418 4910 23420
rect 4966 23418 4972 23420
rect 4726 23366 4728 23418
rect 4908 23366 4910 23418
rect 4664 23364 4670 23366
rect 4726 23364 4750 23366
rect 4806 23364 4830 23366
rect 4886 23364 4910 23366
rect 4966 23364 4972 23366
rect 4664 23355 4972 23364
rect 5000 23322 5028 23666
rect 5080 23656 5132 23662
rect 5080 23598 5132 23604
rect 4988 23316 5040 23322
rect 4988 23258 5040 23264
rect 4528 23112 4580 23118
rect 4528 23054 4580 23060
rect 4988 22568 5040 22574
rect 4988 22510 5040 22516
rect 5000 22438 5028 22510
rect 4988 22432 5040 22438
rect 4988 22374 5040 22380
rect 4664 22332 4972 22341
rect 4664 22330 4670 22332
rect 4726 22330 4750 22332
rect 4806 22330 4830 22332
rect 4886 22330 4910 22332
rect 4966 22330 4972 22332
rect 4726 22278 4728 22330
rect 4908 22278 4910 22330
rect 4664 22276 4670 22278
rect 4726 22276 4750 22278
rect 4806 22276 4830 22278
rect 4886 22276 4910 22278
rect 4966 22276 4972 22278
rect 4664 22267 4972 22276
rect 5000 22030 5028 22374
rect 4988 22024 5040 22030
rect 4988 21966 5040 21972
rect 4344 21616 4396 21622
rect 4344 21558 4396 21564
rect 4664 21244 4972 21253
rect 4664 21242 4670 21244
rect 4726 21242 4750 21244
rect 4806 21242 4830 21244
rect 4886 21242 4910 21244
rect 4966 21242 4972 21244
rect 4726 21190 4728 21242
rect 4908 21190 4910 21242
rect 4664 21188 4670 21190
rect 4726 21188 4750 21190
rect 4806 21188 4830 21190
rect 4886 21188 4910 21190
rect 4966 21188 4972 21190
rect 4664 21179 4972 21188
rect 4160 20800 4212 20806
rect 4160 20742 4212 20748
rect 4068 20528 4120 20534
rect 4068 20470 4120 20476
rect 2504 20392 2556 20398
rect 2504 20334 2556 20340
rect 3976 20392 4028 20398
rect 3976 20334 4028 20340
rect 2516 20058 2544 20334
rect 4080 20058 4108 20470
rect 2504 20052 2556 20058
rect 2504 19994 2556 20000
rect 4068 20052 4120 20058
rect 4068 19994 4120 20000
rect 4172 19854 4200 20742
rect 4664 20156 4972 20165
rect 4664 20154 4670 20156
rect 4726 20154 4750 20156
rect 4806 20154 4830 20156
rect 4886 20154 4910 20156
rect 4966 20154 4972 20156
rect 4726 20102 4728 20154
rect 4908 20102 4910 20154
rect 4664 20100 4670 20102
rect 4726 20100 4750 20102
rect 4806 20100 4830 20102
rect 4886 20100 4910 20102
rect 4966 20100 4972 20102
rect 4664 20091 4972 20100
rect 3884 19848 3936 19854
rect 3884 19790 3936 19796
rect 4160 19848 4212 19854
rect 4160 19790 4212 19796
rect 2136 19712 2188 19718
rect 2136 19654 2188 19660
rect 2148 19446 2176 19654
rect 3896 19446 3924 19790
rect 2136 19440 2188 19446
rect 2136 19382 2188 19388
rect 3884 19440 3936 19446
rect 4172 19394 4200 19790
rect 3884 19382 3936 19388
rect 3240 19372 3292 19378
rect 3240 19314 3292 19320
rect 4080 19366 4200 19394
rect 1860 19304 1912 19310
rect 1860 19246 1912 19252
rect 1872 18970 1900 19246
rect 3252 18970 3280 19314
rect 1860 18964 1912 18970
rect 1860 18906 1912 18912
rect 3240 18964 3292 18970
rect 3240 18906 3292 18912
rect 4080 18766 4108 19366
rect 4664 19068 4972 19077
rect 4664 19066 4670 19068
rect 4726 19066 4750 19068
rect 4806 19066 4830 19068
rect 4886 19066 4910 19068
rect 4966 19066 4972 19068
rect 4726 19014 4728 19066
rect 4908 19014 4910 19066
rect 4664 19012 4670 19014
rect 4726 19012 4750 19014
rect 4806 19012 4830 19014
rect 4886 19012 4910 19014
rect 4966 19012 4972 19014
rect 4664 19003 4972 19012
rect 2504 18760 2556 18766
rect 2504 18702 2556 18708
rect 3424 18760 3476 18766
rect 3424 18702 3476 18708
rect 4068 18760 4120 18766
rect 4068 18702 4120 18708
rect 2516 18426 2544 18702
rect 2504 18420 2556 18426
rect 2504 18362 2556 18368
rect 2044 18216 2096 18222
rect 2044 18158 2096 18164
rect 2320 18216 2372 18222
rect 2320 18158 2372 18164
rect 2056 16590 2084 18158
rect 2332 17882 2360 18158
rect 2320 17876 2372 17882
rect 2320 17818 2372 17824
rect 2516 17678 2544 18362
rect 2780 18352 2832 18358
rect 2780 18294 2832 18300
rect 2792 17882 2820 18294
rect 2780 17876 2832 17882
rect 2780 17818 2832 17824
rect 2504 17672 2556 17678
rect 2504 17614 2556 17620
rect 3332 17672 3384 17678
rect 3436 17660 3464 18702
rect 4664 17980 4972 17989
rect 4664 17978 4670 17980
rect 4726 17978 4750 17980
rect 4806 17978 4830 17980
rect 4886 17978 4910 17980
rect 4966 17978 4972 17980
rect 4726 17926 4728 17978
rect 4908 17926 4910 17978
rect 4664 17924 4670 17926
rect 4726 17924 4750 17926
rect 4806 17924 4830 17926
rect 4886 17924 4910 17926
rect 4966 17924 4972 17926
rect 4664 17915 4972 17924
rect 5092 17678 5120 23598
rect 5184 23254 5212 23666
rect 6748 23322 6776 24754
rect 6736 23316 6788 23322
rect 6736 23258 6788 23264
rect 5172 23248 5224 23254
rect 5172 23190 5224 23196
rect 5184 22642 5212 23190
rect 5816 23112 5868 23118
rect 5816 23054 5868 23060
rect 5172 22636 5224 22642
rect 5172 22578 5224 22584
rect 5264 22568 5316 22574
rect 5264 22510 5316 22516
rect 5276 22166 5304 22510
rect 5828 22234 5856 23054
rect 6092 23044 6144 23050
rect 6092 22986 6144 22992
rect 6104 22778 6132 22986
rect 6092 22772 6144 22778
rect 6092 22714 6144 22720
rect 6748 22642 6776 23258
rect 6840 22642 6868 25230
rect 6932 24206 6960 26318
rect 7012 25220 7064 25226
rect 7012 25162 7064 25168
rect 7024 24954 7052 25162
rect 7012 24948 7064 24954
rect 7012 24890 7064 24896
rect 6920 24200 6972 24206
rect 6920 24142 6972 24148
rect 6932 23798 6960 24142
rect 7104 24064 7156 24070
rect 7104 24006 7156 24012
rect 6920 23792 6972 23798
rect 6920 23734 6972 23740
rect 6736 22636 6788 22642
rect 6736 22578 6788 22584
rect 6828 22636 6880 22642
rect 6828 22578 6880 22584
rect 6840 22438 6868 22578
rect 6828 22432 6880 22438
rect 6828 22374 6880 22380
rect 5816 22228 5868 22234
rect 5816 22170 5868 22176
rect 5264 22160 5316 22166
rect 5264 22102 5316 22108
rect 5276 19854 5304 22102
rect 6828 22094 6880 22098
rect 6932 22094 6960 23734
rect 7116 23050 7144 24006
rect 7104 23044 7156 23050
rect 7104 22986 7156 22992
rect 6828 22092 6960 22094
rect 6880 22066 6960 22092
rect 6828 22034 6880 22040
rect 5724 22024 5776 22030
rect 5724 21966 5776 21972
rect 6092 22024 6144 22030
rect 6092 21966 6144 21972
rect 6460 22024 6512 22030
rect 6460 21966 6512 21972
rect 5736 21622 5764 21966
rect 5724 21616 5776 21622
rect 5724 21558 5776 21564
rect 6104 21486 6132 21966
rect 6092 21480 6144 21486
rect 6092 21422 6144 21428
rect 5540 20936 5592 20942
rect 5540 20878 5592 20884
rect 5552 20602 5580 20878
rect 5540 20596 5592 20602
rect 5540 20538 5592 20544
rect 6104 19854 6132 21422
rect 6276 21344 6328 21350
rect 6276 21286 6328 21292
rect 6288 21010 6316 21286
rect 6276 21004 6328 21010
rect 6276 20946 6328 20952
rect 6472 19854 6500 21966
rect 7012 21956 7064 21962
rect 7012 21898 7064 21904
rect 7024 20874 7052 21898
rect 7012 20868 7064 20874
rect 7012 20810 7064 20816
rect 7104 20528 7156 20534
rect 7104 20470 7156 20476
rect 6552 20392 6604 20398
rect 6552 20334 6604 20340
rect 5264 19848 5316 19854
rect 5264 19790 5316 19796
rect 6092 19848 6144 19854
rect 6092 19790 6144 19796
rect 6460 19848 6512 19854
rect 6460 19790 6512 19796
rect 6564 19718 6592 20334
rect 7116 19922 7144 20470
rect 7208 20398 7236 28494
rect 8300 28416 8352 28422
rect 8300 28358 8352 28364
rect 8312 28082 8340 28358
rect 8378 28316 8686 28325
rect 8378 28314 8384 28316
rect 8440 28314 8464 28316
rect 8520 28314 8544 28316
rect 8600 28314 8624 28316
rect 8680 28314 8686 28316
rect 8440 28262 8442 28314
rect 8622 28262 8624 28314
rect 8378 28260 8384 28262
rect 8440 28260 8464 28262
rect 8520 28260 8544 28262
rect 8600 28260 8624 28262
rect 8680 28260 8686 28262
rect 8378 28251 8686 28260
rect 8300 28076 8352 28082
rect 8300 28018 8352 28024
rect 7380 28008 7432 28014
rect 7380 27950 7432 27956
rect 7656 28008 7708 28014
rect 7656 27950 7708 27956
rect 7392 27538 7420 27950
rect 7380 27532 7432 27538
rect 7380 27474 7432 27480
rect 7392 26518 7420 27474
rect 7668 27402 7696 27950
rect 7656 27396 7708 27402
rect 7656 27338 7708 27344
rect 8772 27334 8800 28494
rect 8852 28416 8904 28422
rect 8852 28358 8904 28364
rect 8864 28150 8892 28358
rect 8852 28144 8904 28150
rect 8852 28086 8904 28092
rect 9680 28076 9732 28082
rect 9680 28018 9732 28024
rect 9692 27606 9720 28018
rect 10336 27946 10364 28494
rect 10876 28416 10928 28422
rect 10876 28358 10928 28364
rect 10324 27940 10376 27946
rect 10324 27882 10376 27888
rect 9680 27600 9732 27606
rect 9680 27542 9732 27548
rect 10888 27470 10916 28358
rect 11072 27690 11100 28494
rect 11152 27872 11204 27878
rect 11152 27814 11204 27820
rect 10980 27674 11100 27690
rect 11164 27674 11192 27814
rect 10968 27668 11100 27674
rect 11020 27662 11100 27668
rect 10968 27610 11020 27616
rect 10876 27464 10928 27470
rect 10876 27406 10928 27412
rect 11072 27334 11100 27662
rect 11152 27668 11204 27674
rect 11152 27610 11204 27616
rect 11716 27538 11744 28494
rect 11796 28484 11848 28490
rect 11796 28426 11848 28432
rect 11704 27532 11756 27538
rect 11704 27474 11756 27480
rect 8760 27328 8812 27334
rect 8760 27270 8812 27276
rect 9312 27328 9364 27334
rect 9312 27270 9364 27276
rect 11060 27328 11112 27334
rect 11060 27270 11112 27276
rect 8378 27228 8686 27237
rect 8378 27226 8384 27228
rect 8440 27226 8464 27228
rect 8520 27226 8544 27228
rect 8600 27226 8624 27228
rect 8680 27226 8686 27228
rect 8440 27174 8442 27226
rect 8622 27174 8624 27226
rect 8378 27172 8384 27174
rect 8440 27172 8464 27174
rect 8520 27172 8544 27174
rect 8600 27172 8624 27174
rect 8680 27172 8686 27174
rect 8378 27163 8686 27172
rect 8300 26988 8352 26994
rect 8300 26930 8352 26936
rect 7380 26512 7432 26518
rect 7380 26454 7432 26460
rect 7288 26308 7340 26314
rect 7288 26250 7340 26256
rect 7300 25974 7328 26250
rect 7288 25968 7340 25974
rect 7288 25910 7340 25916
rect 7392 24274 7420 26454
rect 8024 26444 8076 26450
rect 8024 26386 8076 26392
rect 8036 25498 8064 26386
rect 8312 26382 8340 26930
rect 9324 26382 9352 27270
rect 11716 27062 11744 27474
rect 11808 27402 11836 28426
rect 12072 28416 12124 28422
rect 12072 28358 12124 28364
rect 12084 28082 12112 28358
rect 12728 28218 12756 28494
rect 12716 28212 12768 28218
rect 12716 28154 12768 28160
rect 12072 28076 12124 28082
rect 12072 28018 12124 28024
rect 11888 27940 11940 27946
rect 11888 27882 11940 27888
rect 11796 27396 11848 27402
rect 11796 27338 11848 27344
rect 11704 27056 11756 27062
rect 11704 26998 11756 27004
rect 11900 26994 11928 27882
rect 12092 27772 12400 27781
rect 12092 27770 12098 27772
rect 12154 27770 12178 27772
rect 12234 27770 12258 27772
rect 12314 27770 12338 27772
rect 12394 27770 12400 27772
rect 12154 27718 12156 27770
rect 12336 27718 12338 27770
rect 12092 27716 12098 27718
rect 12154 27716 12178 27718
rect 12234 27716 12258 27718
rect 12314 27716 12338 27718
rect 12394 27716 12400 27718
rect 12092 27707 12400 27716
rect 12728 27334 12756 28154
rect 13360 28144 13412 28150
rect 13360 28086 13412 28092
rect 12716 27328 12768 27334
rect 12716 27270 12768 27276
rect 11888 26988 11940 26994
rect 11888 26930 11940 26936
rect 11796 26920 11848 26926
rect 11796 26862 11848 26868
rect 11808 26586 11836 26862
rect 12092 26684 12400 26693
rect 12092 26682 12098 26684
rect 12154 26682 12178 26684
rect 12234 26682 12258 26684
rect 12314 26682 12338 26684
rect 12394 26682 12400 26684
rect 12154 26630 12156 26682
rect 12336 26630 12338 26682
rect 12092 26628 12098 26630
rect 12154 26628 12178 26630
rect 12234 26628 12258 26630
rect 12314 26628 12338 26630
rect 12394 26628 12400 26630
rect 12092 26619 12400 26628
rect 11796 26580 11848 26586
rect 11796 26522 11848 26528
rect 12164 26580 12216 26586
rect 12164 26522 12216 26528
rect 9680 26444 9732 26450
rect 9680 26386 9732 26392
rect 8300 26376 8352 26382
rect 8300 26318 8352 26324
rect 9312 26376 9364 26382
rect 9312 26318 9364 26324
rect 8312 26042 8340 26318
rect 8378 26140 8686 26149
rect 8378 26138 8384 26140
rect 8440 26138 8464 26140
rect 8520 26138 8544 26140
rect 8600 26138 8624 26140
rect 8680 26138 8686 26140
rect 8440 26086 8442 26138
rect 8622 26086 8624 26138
rect 8378 26084 8384 26086
rect 8440 26084 8464 26086
rect 8520 26084 8544 26086
rect 8600 26084 8624 26086
rect 8680 26084 8686 26086
rect 8378 26075 8686 26084
rect 8300 26036 8352 26042
rect 8300 25978 8352 25984
rect 9496 25900 9548 25906
rect 9496 25842 9548 25848
rect 9128 25696 9180 25702
rect 9128 25638 9180 25644
rect 8024 25492 8076 25498
rect 8024 25434 8076 25440
rect 8036 24954 8064 25434
rect 8378 25052 8686 25061
rect 8378 25050 8384 25052
rect 8440 25050 8464 25052
rect 8520 25050 8544 25052
rect 8600 25050 8624 25052
rect 8680 25050 8686 25052
rect 8440 24998 8442 25050
rect 8622 24998 8624 25050
rect 8378 24996 8384 24998
rect 8440 24996 8464 24998
rect 8520 24996 8544 24998
rect 8600 24996 8624 24998
rect 8680 24996 8686 24998
rect 8378 24987 8686 24996
rect 8024 24948 8076 24954
rect 8024 24890 8076 24896
rect 8760 24812 8812 24818
rect 8760 24754 8812 24760
rect 8116 24608 8168 24614
rect 8116 24550 8168 24556
rect 7380 24268 7432 24274
rect 7380 24210 7432 24216
rect 7392 21486 7420 24210
rect 8128 22710 8156 24550
rect 8378 23964 8686 23973
rect 8378 23962 8384 23964
rect 8440 23962 8464 23964
rect 8520 23962 8544 23964
rect 8600 23962 8624 23964
rect 8680 23962 8686 23964
rect 8440 23910 8442 23962
rect 8622 23910 8624 23962
rect 8378 23908 8384 23910
rect 8440 23908 8464 23910
rect 8520 23908 8544 23910
rect 8600 23908 8624 23910
rect 8680 23908 8686 23910
rect 8378 23899 8686 23908
rect 8772 23186 8800 24754
rect 8760 23180 8812 23186
rect 8760 23122 8812 23128
rect 8378 22876 8686 22885
rect 8378 22874 8384 22876
rect 8440 22874 8464 22876
rect 8520 22874 8544 22876
rect 8600 22874 8624 22876
rect 8680 22874 8686 22876
rect 8440 22822 8442 22874
rect 8622 22822 8624 22874
rect 8378 22820 8384 22822
rect 8440 22820 8464 22822
rect 8520 22820 8544 22822
rect 8600 22820 8624 22822
rect 8680 22820 8686 22822
rect 8378 22811 8686 22820
rect 8772 22778 8800 23122
rect 8760 22772 8812 22778
rect 8760 22714 8812 22720
rect 8116 22704 8168 22710
rect 8116 22646 8168 22652
rect 8760 22636 8812 22642
rect 8760 22578 8812 22584
rect 8378 21788 8686 21797
rect 8378 21786 8384 21788
rect 8440 21786 8464 21788
rect 8520 21786 8544 21788
rect 8600 21786 8624 21788
rect 8680 21786 8686 21788
rect 8440 21734 8442 21786
rect 8622 21734 8624 21786
rect 8378 21732 8384 21734
rect 8440 21732 8464 21734
rect 8520 21732 8544 21734
rect 8600 21732 8624 21734
rect 8680 21732 8686 21734
rect 8378 21723 8686 21732
rect 8772 21622 8800 22578
rect 9140 22166 9168 25638
rect 9508 25498 9536 25842
rect 9496 25492 9548 25498
rect 9496 25434 9548 25440
rect 9692 23662 9720 26386
rect 10232 26376 10284 26382
rect 10232 26318 10284 26324
rect 11152 26376 11204 26382
rect 11152 26318 11204 26324
rect 10244 26042 10272 26318
rect 10232 26036 10284 26042
rect 10232 25978 10284 25984
rect 10244 25294 10272 25978
rect 11164 25430 11192 26318
rect 11704 26308 11756 26314
rect 11704 26250 11756 26256
rect 11716 26042 11744 26250
rect 12176 26042 12204 26522
rect 11704 26036 11756 26042
rect 11704 25978 11756 25984
rect 12164 26036 12216 26042
rect 12164 25978 12216 25984
rect 11704 25900 11756 25906
rect 11704 25842 11756 25848
rect 11152 25424 11204 25430
rect 11152 25366 11204 25372
rect 10232 25288 10284 25294
rect 10232 25230 10284 25236
rect 10784 25220 10836 25226
rect 10784 25162 10836 25168
rect 9864 25152 9916 25158
rect 9864 25094 9916 25100
rect 9680 23656 9732 23662
rect 9680 23598 9732 23604
rect 9772 22704 9824 22710
rect 9772 22646 9824 22652
rect 9680 22568 9732 22574
rect 9680 22510 9732 22516
rect 9128 22160 9180 22166
rect 9128 22102 9180 22108
rect 8760 21616 8812 21622
rect 8760 21558 8812 21564
rect 8024 21548 8076 21554
rect 8024 21490 8076 21496
rect 7380 21480 7432 21486
rect 7380 21422 7432 21428
rect 7196 20392 7248 20398
rect 7196 20334 7248 20340
rect 7104 19916 7156 19922
rect 7104 19858 7156 19864
rect 6184 19712 6236 19718
rect 6184 19654 6236 19660
rect 6552 19712 6604 19718
rect 6552 19654 6604 19660
rect 5724 18692 5776 18698
rect 5724 18634 5776 18640
rect 5736 18290 5764 18634
rect 5724 18284 5776 18290
rect 5724 18226 5776 18232
rect 5736 17678 5764 18226
rect 6000 18148 6052 18154
rect 6000 18090 6052 18096
rect 5816 18080 5868 18086
rect 5816 18022 5868 18028
rect 3384 17632 3464 17660
rect 3332 17614 3384 17620
rect 3332 17536 3384 17542
rect 3332 17478 3384 17484
rect 2872 17196 2924 17202
rect 2872 17138 2924 17144
rect 2884 16726 2912 17138
rect 2964 16992 3016 16998
rect 2964 16934 3016 16940
rect 2872 16720 2924 16726
rect 2872 16662 2924 16668
rect 2044 16584 2096 16590
rect 2044 16526 2096 16532
rect 2976 16182 3004 16934
rect 2964 16176 3016 16182
rect 2964 16118 3016 16124
rect 3344 16046 3372 17478
rect 3436 17202 3464 17632
rect 3976 17672 4028 17678
rect 3976 17614 4028 17620
rect 5080 17672 5132 17678
rect 5080 17614 5132 17620
rect 5724 17672 5776 17678
rect 5724 17614 5776 17620
rect 3988 17270 4016 17614
rect 3976 17264 4028 17270
rect 3976 17206 4028 17212
rect 3424 17196 3476 17202
rect 3424 17138 3476 17144
rect 3424 16992 3476 16998
rect 3424 16934 3476 16940
rect 3436 16182 3464 16934
rect 3988 16658 4016 17206
rect 4664 16892 4972 16901
rect 4664 16890 4670 16892
rect 4726 16890 4750 16892
rect 4806 16890 4830 16892
rect 4886 16890 4910 16892
rect 4966 16890 4972 16892
rect 4726 16838 4728 16890
rect 4908 16838 4910 16890
rect 4664 16836 4670 16838
rect 4726 16836 4750 16838
rect 4806 16836 4830 16838
rect 4886 16836 4910 16838
rect 4966 16836 4972 16838
rect 4664 16827 4972 16836
rect 4712 16720 4764 16726
rect 4712 16662 4764 16668
rect 3976 16652 4028 16658
rect 3976 16594 4028 16600
rect 4724 16182 4752 16662
rect 3424 16176 3476 16182
rect 3424 16118 3476 16124
rect 4712 16176 4764 16182
rect 4712 16118 4764 16124
rect 3332 16040 3384 16046
rect 3332 15982 3384 15988
rect 4664 15804 4972 15813
rect 4664 15802 4670 15804
rect 4726 15802 4750 15804
rect 4806 15802 4830 15804
rect 4886 15802 4910 15804
rect 4966 15802 4972 15804
rect 4726 15750 4728 15802
rect 4908 15750 4910 15802
rect 4664 15748 4670 15750
rect 4726 15748 4750 15750
rect 4806 15748 4830 15750
rect 4886 15748 4910 15750
rect 4966 15748 4972 15750
rect 4664 15739 4972 15748
rect 4436 15360 4488 15366
rect 4436 15302 4488 15308
rect 4448 14006 4476 15302
rect 4664 14716 4972 14725
rect 4664 14714 4670 14716
rect 4726 14714 4750 14716
rect 4806 14714 4830 14716
rect 4886 14714 4910 14716
rect 4966 14714 4972 14716
rect 4726 14662 4728 14714
rect 4908 14662 4910 14714
rect 4664 14660 4670 14662
rect 4726 14660 4750 14662
rect 4806 14660 4830 14662
rect 4886 14660 4910 14662
rect 4966 14660 4972 14662
rect 4664 14651 4972 14660
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 4632 14074 4660 14350
rect 4620 14068 4672 14074
rect 4620 14010 4672 14016
rect 4436 14000 4488 14006
rect 4436 13942 4488 13948
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 4172 13530 4200 13806
rect 4664 13628 4972 13637
rect 4664 13626 4670 13628
rect 4726 13626 4750 13628
rect 4806 13626 4830 13628
rect 4886 13626 4910 13628
rect 4966 13626 4972 13628
rect 4726 13574 4728 13626
rect 4908 13574 4910 13626
rect 4664 13572 4670 13574
rect 4726 13572 4750 13574
rect 4806 13572 4830 13574
rect 4886 13572 4910 13574
rect 4966 13572 4972 13574
rect 4664 13563 4972 13572
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 4988 13320 5040 13326
rect 4988 13262 5040 13268
rect 4664 12540 4972 12549
rect 4664 12538 4670 12540
rect 4726 12538 4750 12540
rect 4806 12538 4830 12540
rect 4886 12538 4910 12540
rect 4966 12538 4972 12540
rect 4726 12486 4728 12538
rect 4908 12486 4910 12538
rect 4664 12484 4670 12486
rect 4726 12484 4750 12486
rect 4806 12484 4830 12486
rect 4886 12484 4910 12486
rect 4966 12484 4972 12486
rect 4664 12475 4972 12484
rect 5000 12238 5028 13262
rect 4988 12232 5040 12238
rect 4988 12174 5040 12180
rect 4160 12164 4212 12170
rect 4160 12106 4212 12112
rect 4172 11762 4200 12106
rect 4436 12096 4488 12102
rect 4436 12038 4488 12044
rect 4448 11830 4476 12038
rect 4436 11824 4488 11830
rect 4436 11766 4488 11772
rect 4160 11756 4212 11762
rect 4160 11698 4212 11704
rect 5000 11694 5028 12174
rect 4988 11688 5040 11694
rect 4988 11630 5040 11636
rect 4664 11452 4972 11461
rect 4664 11450 4670 11452
rect 4726 11450 4750 11452
rect 4806 11450 4830 11452
rect 4886 11450 4910 11452
rect 4966 11450 4972 11452
rect 4726 11398 4728 11450
rect 4908 11398 4910 11450
rect 4664 11396 4670 11398
rect 4726 11396 4750 11398
rect 4806 11396 4830 11398
rect 4886 11396 4910 11398
rect 4966 11396 4972 11398
rect 4664 11387 4972 11396
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 4264 10810 4292 11086
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 4988 10736 5040 10742
rect 4988 10678 5040 10684
rect 4664 10364 4972 10373
rect 4664 10362 4670 10364
rect 4726 10362 4750 10364
rect 4806 10362 4830 10364
rect 4886 10362 4910 10364
rect 4966 10362 4972 10364
rect 4726 10310 4728 10362
rect 4908 10310 4910 10362
rect 4664 10308 4670 10310
rect 4726 10308 4750 10310
rect 4806 10308 4830 10310
rect 4886 10308 4910 10310
rect 4966 10308 4972 10310
rect 4664 10299 4972 10308
rect 5000 9654 5028 10678
rect 4988 9648 5040 9654
rect 4988 9590 5040 9596
rect 4664 9276 4972 9285
rect 4664 9274 4670 9276
rect 4726 9274 4750 9276
rect 4806 9274 4830 9276
rect 4886 9274 4910 9276
rect 4966 9274 4972 9276
rect 4726 9222 4728 9274
rect 4908 9222 4910 9274
rect 4664 9220 4670 9222
rect 4726 9220 4750 9222
rect 4806 9220 4830 9222
rect 4886 9220 4910 9222
rect 4966 9220 4972 9222
rect 4664 9211 4972 9220
rect 4664 8188 4972 8197
rect 4664 8186 4670 8188
rect 4726 8186 4750 8188
rect 4806 8186 4830 8188
rect 4886 8186 4910 8188
rect 4966 8186 4972 8188
rect 4726 8134 4728 8186
rect 4908 8134 4910 8186
rect 4664 8132 4670 8134
rect 4726 8132 4750 8134
rect 4806 8132 4830 8134
rect 4886 8132 4910 8134
rect 4966 8132 4972 8134
rect 4664 8123 4972 8132
rect 4664 7100 4972 7109
rect 4664 7098 4670 7100
rect 4726 7098 4750 7100
rect 4806 7098 4830 7100
rect 4886 7098 4910 7100
rect 4966 7098 4972 7100
rect 4726 7046 4728 7098
rect 4908 7046 4910 7098
rect 4664 7044 4670 7046
rect 4726 7044 4750 7046
rect 4806 7044 4830 7046
rect 4886 7044 4910 7046
rect 4966 7044 4972 7046
rect 4664 7035 4972 7044
rect 5092 6390 5120 17614
rect 5736 17338 5764 17614
rect 5724 17332 5776 17338
rect 5724 17274 5776 17280
rect 5828 17270 5856 18022
rect 5816 17264 5868 17270
rect 5816 17206 5868 17212
rect 6012 17202 6040 18090
rect 6000 17196 6052 17202
rect 6000 17138 6052 17144
rect 5724 17128 5776 17134
rect 5724 17070 5776 17076
rect 5736 16590 5764 17070
rect 6196 16590 6224 19654
rect 6564 18426 6592 19654
rect 7472 18624 7524 18630
rect 7472 18566 7524 18572
rect 6552 18420 6604 18426
rect 6552 18362 6604 18368
rect 7484 18358 7512 18566
rect 7472 18352 7524 18358
rect 7472 18294 7524 18300
rect 6736 18284 6788 18290
rect 6736 18226 6788 18232
rect 6552 17672 6604 17678
rect 6552 17614 6604 17620
rect 5724 16584 5776 16590
rect 5724 16526 5776 16532
rect 6184 16584 6236 16590
rect 6184 16526 6236 16532
rect 6460 16516 6512 16522
rect 6460 16458 6512 16464
rect 6184 16040 6236 16046
rect 6184 15982 6236 15988
rect 6196 15706 6224 15982
rect 6472 15706 6500 16458
rect 6184 15700 6236 15706
rect 6184 15642 6236 15648
rect 6460 15700 6512 15706
rect 6460 15642 6512 15648
rect 5172 15496 5224 15502
rect 5172 15438 5224 15444
rect 5184 14074 5212 15438
rect 5264 15020 5316 15026
rect 5264 14962 5316 14968
rect 5172 14068 5224 14074
rect 5172 14010 5224 14016
rect 5276 13394 5304 14962
rect 5356 14952 5408 14958
rect 5356 14894 5408 14900
rect 5908 14952 5960 14958
rect 5908 14894 5960 14900
rect 5264 13388 5316 13394
rect 5264 13330 5316 13336
rect 5276 12850 5304 13330
rect 5368 12850 5396 14894
rect 5920 14346 5948 14894
rect 5908 14340 5960 14346
rect 5908 14282 5960 14288
rect 5816 14000 5868 14006
rect 5816 13942 5868 13948
rect 5828 12986 5856 13942
rect 6196 13870 6224 15642
rect 6564 15026 6592 17614
rect 6748 17610 6776 18226
rect 6736 17604 6788 17610
rect 6736 17546 6788 17552
rect 7472 17604 7524 17610
rect 7472 17546 7524 17552
rect 6748 17202 6776 17546
rect 6828 17536 6880 17542
rect 6828 17478 6880 17484
rect 6840 17338 6868 17478
rect 7484 17338 7512 17546
rect 6828 17332 6880 17338
rect 6828 17274 6880 17280
rect 7472 17332 7524 17338
rect 7472 17274 7524 17280
rect 6736 17196 6788 17202
rect 6736 17138 6788 17144
rect 7288 15904 7340 15910
rect 7288 15846 7340 15852
rect 6828 15700 6880 15706
rect 6828 15642 6880 15648
rect 6552 15020 6604 15026
rect 6552 14962 6604 14968
rect 6564 14618 6592 14962
rect 6552 14612 6604 14618
rect 6552 14554 6604 14560
rect 6736 14340 6788 14346
rect 6736 14282 6788 14288
rect 6748 13938 6776 14282
rect 6736 13932 6788 13938
rect 6736 13874 6788 13880
rect 6184 13864 6236 13870
rect 6184 13806 6236 13812
rect 5816 12980 5868 12986
rect 5816 12922 5868 12928
rect 5264 12844 5316 12850
rect 5264 12786 5316 12792
rect 5356 12844 5408 12850
rect 5356 12786 5408 12792
rect 5368 12434 5396 12786
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 5276 12406 5396 12434
rect 5172 12232 5224 12238
rect 5172 12174 5224 12180
rect 5184 11218 5212 12174
rect 5276 11218 5304 12406
rect 5172 11212 5224 11218
rect 5172 11154 5224 11160
rect 5264 11212 5316 11218
rect 5264 11154 5316 11160
rect 5460 11150 5488 12718
rect 5724 11824 5776 11830
rect 5724 11766 5776 11772
rect 5736 11218 5764 11766
rect 6840 11694 6868 15642
rect 7300 15502 7328 15846
rect 7288 15496 7340 15502
rect 7288 15438 7340 15444
rect 8036 15162 8064 21490
rect 8772 21078 8800 21558
rect 9036 21480 9088 21486
rect 9140 21468 9168 22102
rect 9692 21690 9720 22510
rect 9680 21684 9732 21690
rect 9680 21626 9732 21632
rect 9312 21548 9364 21554
rect 9312 21490 9364 21496
rect 9088 21440 9168 21468
rect 9036 21422 9088 21428
rect 8760 21072 8812 21078
rect 8760 21014 8812 21020
rect 8378 20700 8686 20709
rect 8378 20698 8384 20700
rect 8440 20698 8464 20700
rect 8520 20698 8544 20700
rect 8600 20698 8624 20700
rect 8680 20698 8686 20700
rect 8440 20646 8442 20698
rect 8622 20646 8624 20698
rect 8378 20644 8384 20646
rect 8440 20644 8464 20646
rect 8520 20644 8544 20646
rect 8600 20644 8624 20646
rect 8680 20644 8686 20646
rect 8378 20635 8686 20644
rect 8378 19612 8686 19621
rect 8378 19610 8384 19612
rect 8440 19610 8464 19612
rect 8520 19610 8544 19612
rect 8600 19610 8624 19612
rect 8680 19610 8686 19612
rect 8440 19558 8442 19610
rect 8622 19558 8624 19610
rect 8378 19556 8384 19558
rect 8440 19556 8464 19558
rect 8520 19556 8544 19558
rect 8600 19556 8624 19558
rect 8680 19556 8686 19558
rect 8378 19547 8686 19556
rect 8760 18624 8812 18630
rect 8760 18566 8812 18572
rect 8378 18524 8686 18533
rect 8378 18522 8384 18524
rect 8440 18522 8464 18524
rect 8520 18522 8544 18524
rect 8600 18522 8624 18524
rect 8680 18522 8686 18524
rect 8440 18470 8442 18522
rect 8622 18470 8624 18522
rect 8378 18468 8384 18470
rect 8440 18468 8464 18470
rect 8520 18468 8544 18470
rect 8600 18468 8624 18470
rect 8680 18468 8686 18470
rect 8378 18459 8686 18468
rect 8772 18358 8800 18566
rect 8760 18352 8812 18358
rect 8760 18294 8812 18300
rect 8378 17436 8686 17445
rect 8378 17434 8384 17436
rect 8440 17434 8464 17436
rect 8520 17434 8544 17436
rect 8600 17434 8624 17436
rect 8680 17434 8686 17436
rect 8440 17382 8442 17434
rect 8622 17382 8624 17434
rect 8378 17380 8384 17382
rect 8440 17380 8464 17382
rect 8520 17380 8544 17382
rect 8600 17380 8624 17382
rect 8680 17380 8686 17382
rect 8378 17371 8686 17380
rect 8300 16516 8352 16522
rect 8300 16458 8352 16464
rect 8312 15910 8340 16458
rect 8378 16348 8686 16357
rect 8378 16346 8384 16348
rect 8440 16346 8464 16348
rect 8520 16346 8544 16348
rect 8600 16346 8624 16348
rect 8680 16346 8686 16348
rect 8440 16294 8442 16346
rect 8622 16294 8624 16346
rect 8378 16292 8384 16294
rect 8440 16292 8464 16294
rect 8520 16292 8544 16294
rect 8600 16292 8624 16294
rect 8680 16292 8686 16294
rect 8378 16283 8686 16292
rect 8300 15904 8352 15910
rect 8300 15846 8352 15852
rect 8024 15156 8076 15162
rect 8024 15098 8076 15104
rect 7196 13864 7248 13870
rect 7196 13806 7248 13812
rect 6920 12912 6972 12918
rect 6920 12854 6972 12860
rect 6932 12238 6960 12854
rect 7104 12844 7156 12850
rect 7104 12786 7156 12792
rect 7116 12238 7144 12786
rect 7208 12238 7236 13806
rect 8036 13326 8064 15098
rect 8024 13320 8076 13326
rect 8024 13262 8076 13268
rect 7656 12844 7708 12850
rect 7656 12786 7708 12792
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 7104 12232 7156 12238
rect 7104 12174 7156 12180
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 7668 11898 7696 12786
rect 8312 12782 8340 15846
rect 9048 15502 9076 21422
rect 9324 21078 9352 21490
rect 9312 21072 9364 21078
rect 9312 21014 9364 21020
rect 9692 21010 9720 21626
rect 9680 21004 9732 21010
rect 9680 20946 9732 20952
rect 9312 20460 9364 20466
rect 9312 20402 9364 20408
rect 9324 20058 9352 20402
rect 9784 20262 9812 22646
rect 9772 20256 9824 20262
rect 9772 20198 9824 20204
rect 9312 20052 9364 20058
rect 9312 19994 9364 20000
rect 9876 19854 9904 25094
rect 9956 24744 10008 24750
rect 9956 24686 10008 24692
rect 9968 21010 9996 24686
rect 10796 23798 10824 25162
rect 11716 24954 11744 25842
rect 11980 25832 12032 25838
rect 11980 25774 12032 25780
rect 11992 25362 12020 25774
rect 12092 25596 12400 25605
rect 12092 25594 12098 25596
rect 12154 25594 12178 25596
rect 12234 25594 12258 25596
rect 12314 25594 12338 25596
rect 12394 25594 12400 25596
rect 12154 25542 12156 25594
rect 12336 25542 12338 25594
rect 12092 25540 12098 25542
rect 12154 25540 12178 25542
rect 12234 25540 12258 25542
rect 12314 25540 12338 25542
rect 12394 25540 12400 25542
rect 12092 25531 12400 25540
rect 11796 25356 11848 25362
rect 11796 25298 11848 25304
rect 11980 25356 12032 25362
rect 11980 25298 12032 25304
rect 11152 24948 11204 24954
rect 11152 24890 11204 24896
rect 11704 24948 11756 24954
rect 11704 24890 11756 24896
rect 10784 23792 10836 23798
rect 10784 23734 10836 23740
rect 10416 23724 10468 23730
rect 10416 23666 10468 23672
rect 10140 23520 10192 23526
rect 10140 23462 10192 23468
rect 10152 23322 10180 23462
rect 10140 23316 10192 23322
rect 10140 23258 10192 23264
rect 10428 22574 10456 23666
rect 10796 23118 10824 23734
rect 11060 23724 11112 23730
rect 11060 23666 11112 23672
rect 10784 23112 10836 23118
rect 10784 23054 10836 23060
rect 10416 22568 10468 22574
rect 10416 22510 10468 22516
rect 10140 22092 10192 22098
rect 10140 22034 10192 22040
rect 10416 22092 10468 22098
rect 10416 22034 10468 22040
rect 10048 22024 10100 22030
rect 10048 21966 10100 21972
rect 9956 21004 10008 21010
rect 9956 20946 10008 20952
rect 9968 20534 9996 20946
rect 10060 20602 10088 21966
rect 10152 20602 10180 22034
rect 10428 21554 10456 22034
rect 10876 21888 10928 21894
rect 10876 21830 10928 21836
rect 10416 21548 10468 21554
rect 10416 21490 10468 21496
rect 10888 20942 10916 21830
rect 11072 21622 11100 23666
rect 11164 22574 11192 24890
rect 11336 24676 11388 24682
rect 11336 24618 11388 24624
rect 11348 24274 11376 24618
rect 11612 24608 11664 24614
rect 11612 24550 11664 24556
rect 11624 24274 11652 24550
rect 11336 24268 11388 24274
rect 11336 24210 11388 24216
rect 11612 24268 11664 24274
rect 11612 24210 11664 24216
rect 11244 23656 11296 23662
rect 11244 23598 11296 23604
rect 11256 23254 11284 23598
rect 11520 23520 11572 23526
rect 11520 23462 11572 23468
rect 11244 23248 11296 23254
rect 11244 23190 11296 23196
rect 11532 22710 11560 23462
rect 11520 22704 11572 22710
rect 11520 22646 11572 22652
rect 11428 22636 11480 22642
rect 11428 22578 11480 22584
rect 11152 22568 11204 22574
rect 11152 22510 11204 22516
rect 11164 22094 11192 22510
rect 11440 22098 11468 22578
rect 11164 22066 11284 22094
rect 11152 21888 11204 21894
rect 11256 21876 11284 22066
rect 11428 22092 11480 22098
rect 11428 22034 11480 22040
rect 11204 21848 11284 21876
rect 11152 21830 11204 21836
rect 11060 21616 11112 21622
rect 11060 21558 11112 21564
rect 10600 20936 10652 20942
rect 10600 20878 10652 20884
rect 10876 20936 10928 20942
rect 10876 20878 10928 20884
rect 10048 20596 10100 20602
rect 10048 20538 10100 20544
rect 10140 20596 10192 20602
rect 10140 20538 10192 20544
rect 9956 20528 10008 20534
rect 9956 20470 10008 20476
rect 9968 19990 9996 20470
rect 9956 19984 10008 19990
rect 9956 19926 10008 19932
rect 10152 19854 10180 20538
rect 10612 20262 10640 20878
rect 10600 20256 10652 20262
rect 10600 20198 10652 20204
rect 9864 19848 9916 19854
rect 9864 19790 9916 19796
rect 10140 19848 10192 19854
rect 10140 19790 10192 19796
rect 10612 19378 10640 20198
rect 10876 19712 10928 19718
rect 10876 19654 10928 19660
rect 10600 19372 10652 19378
rect 10600 19314 10652 19320
rect 9220 18760 9272 18766
rect 9220 18702 9272 18708
rect 9128 18624 9180 18630
rect 9128 18566 9180 18572
rect 9140 17746 9168 18566
rect 9232 18358 9260 18702
rect 9220 18352 9272 18358
rect 9220 18294 9272 18300
rect 10888 18290 10916 19654
rect 11164 18766 11192 21830
rect 11440 20806 11468 22034
rect 11716 20874 11744 24890
rect 11808 22166 11836 25298
rect 12092 24508 12400 24517
rect 12092 24506 12098 24508
rect 12154 24506 12178 24508
rect 12234 24506 12258 24508
rect 12314 24506 12338 24508
rect 12394 24506 12400 24508
rect 12154 24454 12156 24506
rect 12336 24454 12338 24506
rect 12092 24452 12098 24454
rect 12154 24452 12178 24454
rect 12234 24452 12258 24454
rect 12314 24452 12338 24454
rect 12394 24452 12400 24454
rect 12092 24443 12400 24452
rect 12624 24132 12676 24138
rect 12624 24074 12676 24080
rect 12636 23798 12664 24074
rect 11980 23792 12032 23798
rect 11980 23734 12032 23740
rect 12624 23792 12676 23798
rect 12624 23734 12676 23740
rect 11992 23322 12020 23734
rect 12092 23420 12400 23429
rect 12092 23418 12098 23420
rect 12154 23418 12178 23420
rect 12234 23418 12258 23420
rect 12314 23418 12338 23420
rect 12394 23418 12400 23420
rect 12154 23366 12156 23418
rect 12336 23366 12338 23418
rect 12092 23364 12098 23366
rect 12154 23364 12178 23366
rect 12234 23364 12258 23366
rect 12314 23364 12338 23366
rect 12394 23364 12400 23366
rect 12092 23355 12400 23364
rect 11980 23316 12032 23322
rect 11980 23258 12032 23264
rect 12728 22642 12756 27270
rect 13372 27062 13400 28086
rect 13636 28008 13688 28014
rect 13636 27950 13688 27956
rect 13648 27606 13676 27950
rect 13740 27946 13768 28494
rect 13820 28212 13872 28218
rect 13820 28154 13872 28160
rect 13728 27940 13780 27946
rect 13728 27882 13780 27888
rect 13636 27600 13688 27606
rect 13636 27542 13688 27548
rect 13360 27056 13412 27062
rect 13360 26998 13412 27004
rect 12900 26784 12952 26790
rect 12900 26726 12952 26732
rect 12912 25974 12940 26726
rect 12992 26376 13044 26382
rect 12992 26318 13044 26324
rect 12900 25968 12952 25974
rect 12900 25910 12952 25916
rect 13004 25838 13032 26318
rect 12992 25832 13044 25838
rect 12992 25774 13044 25780
rect 13176 25696 13228 25702
rect 13176 25638 13228 25644
rect 12992 23656 13044 23662
rect 12992 23598 13044 23604
rect 12716 22636 12768 22642
rect 12716 22578 12768 22584
rect 12532 22432 12584 22438
rect 12532 22374 12584 22380
rect 12092 22332 12400 22341
rect 12092 22330 12098 22332
rect 12154 22330 12178 22332
rect 12234 22330 12258 22332
rect 12314 22330 12338 22332
rect 12394 22330 12400 22332
rect 12154 22278 12156 22330
rect 12336 22278 12338 22330
rect 12092 22276 12098 22278
rect 12154 22276 12178 22278
rect 12234 22276 12258 22278
rect 12314 22276 12338 22278
rect 12394 22276 12400 22278
rect 12092 22267 12400 22276
rect 11796 22160 11848 22166
rect 11796 22102 11848 22108
rect 12256 21888 12308 21894
rect 12256 21830 12308 21836
rect 12440 21888 12492 21894
rect 12440 21830 12492 21836
rect 12268 21554 12296 21830
rect 12452 21622 12480 21830
rect 12544 21622 12572 22374
rect 12440 21616 12492 21622
rect 12440 21558 12492 21564
rect 12532 21616 12584 21622
rect 12532 21558 12584 21564
rect 12256 21548 12308 21554
rect 12256 21490 12308 21496
rect 12624 21548 12676 21554
rect 12624 21490 12676 21496
rect 12092 21244 12400 21253
rect 12092 21242 12098 21244
rect 12154 21242 12178 21244
rect 12234 21242 12258 21244
rect 12314 21242 12338 21244
rect 12394 21242 12400 21244
rect 12154 21190 12156 21242
rect 12336 21190 12338 21242
rect 12092 21188 12098 21190
rect 12154 21188 12178 21190
rect 12234 21188 12258 21190
rect 12314 21188 12338 21190
rect 12394 21188 12400 21190
rect 12092 21179 12400 21188
rect 12636 21078 12664 21490
rect 12624 21072 12676 21078
rect 12624 21014 12676 21020
rect 12728 20942 12756 22578
rect 13004 22030 13032 23598
rect 13188 22642 13216 25638
rect 13360 24744 13412 24750
rect 13360 24686 13412 24692
rect 13372 24274 13400 24686
rect 13360 24268 13412 24274
rect 13360 24210 13412 24216
rect 13372 23118 13400 24210
rect 13452 24200 13504 24206
rect 13452 24142 13504 24148
rect 13464 23866 13492 24142
rect 13452 23860 13504 23866
rect 13452 23802 13504 23808
rect 13740 23730 13768 27882
rect 13832 27470 13860 28154
rect 13820 27464 13872 27470
rect 13820 27406 13872 27412
rect 14096 27464 14148 27470
rect 14096 27406 14148 27412
rect 14108 26994 14136 27406
rect 14096 26988 14148 26994
rect 14096 26930 14148 26936
rect 14108 24818 14136 26930
rect 14004 24812 14056 24818
rect 14004 24754 14056 24760
rect 14096 24812 14148 24818
rect 14096 24754 14148 24760
rect 14016 23730 14044 24754
rect 14096 24132 14148 24138
rect 14096 24074 14148 24080
rect 14108 23866 14136 24074
rect 14096 23860 14148 23866
rect 14096 23802 14148 23808
rect 13728 23724 13780 23730
rect 13728 23666 13780 23672
rect 14004 23724 14056 23730
rect 14004 23666 14056 23672
rect 13360 23112 13412 23118
rect 13360 23054 13412 23060
rect 13176 22636 13228 22642
rect 13176 22578 13228 22584
rect 13084 22500 13136 22506
rect 13084 22442 13136 22448
rect 12992 22024 13044 22030
rect 12992 21966 13044 21972
rect 13096 21690 13124 22442
rect 13176 21956 13228 21962
rect 13176 21898 13228 21904
rect 13084 21684 13136 21690
rect 13084 21626 13136 21632
rect 13188 21350 13216 21898
rect 13176 21344 13228 21350
rect 13176 21286 13228 21292
rect 13820 21140 13872 21146
rect 13820 21082 13872 21088
rect 12716 20936 12768 20942
rect 12716 20878 12768 20884
rect 11704 20868 11756 20874
rect 11704 20810 11756 20816
rect 11428 20800 11480 20806
rect 11428 20742 11480 20748
rect 12092 20156 12400 20165
rect 12092 20154 12098 20156
rect 12154 20154 12178 20156
rect 12234 20154 12258 20156
rect 12314 20154 12338 20156
rect 12394 20154 12400 20156
rect 12154 20102 12156 20154
rect 12336 20102 12338 20154
rect 12092 20100 12098 20102
rect 12154 20100 12178 20102
rect 12234 20100 12258 20102
rect 12314 20100 12338 20102
rect 12394 20100 12400 20102
rect 12092 20091 12400 20100
rect 12900 19372 12952 19378
rect 12900 19314 12952 19320
rect 12992 19372 13044 19378
rect 12992 19314 13044 19320
rect 12092 19068 12400 19077
rect 12092 19066 12098 19068
rect 12154 19066 12178 19068
rect 12234 19066 12258 19068
rect 12314 19066 12338 19068
rect 12394 19066 12400 19068
rect 12154 19014 12156 19066
rect 12336 19014 12338 19066
rect 12092 19012 12098 19014
rect 12154 19012 12178 19014
rect 12234 19012 12258 19014
rect 12314 19012 12338 19014
rect 12394 19012 12400 19014
rect 12092 19003 12400 19012
rect 12348 18828 12400 18834
rect 12348 18770 12400 18776
rect 11152 18760 11204 18766
rect 11152 18702 11204 18708
rect 10876 18284 10928 18290
rect 10876 18226 10928 18232
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 9784 17746 9812 18022
rect 10888 17814 10916 18226
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 10876 17808 10928 17814
rect 10876 17750 10928 17756
rect 9128 17740 9180 17746
rect 9128 17682 9180 17688
rect 9772 17740 9824 17746
rect 9772 17682 9824 17688
rect 10968 17604 11020 17610
rect 10968 17546 11020 17552
rect 9588 16652 9640 16658
rect 9588 16594 9640 16600
rect 9128 16448 9180 16454
rect 9128 16390 9180 16396
rect 9496 16448 9548 16454
rect 9496 16390 9548 16396
rect 9140 16182 9168 16390
rect 9128 16176 9180 16182
rect 9128 16118 9180 16124
rect 9312 15904 9364 15910
rect 9312 15846 9364 15852
rect 9324 15706 9352 15846
rect 9128 15700 9180 15706
rect 9128 15642 9180 15648
rect 9312 15700 9364 15706
rect 9312 15642 9364 15648
rect 9036 15496 9088 15502
rect 9036 15438 9088 15444
rect 8378 15260 8686 15269
rect 8378 15258 8384 15260
rect 8440 15258 8464 15260
rect 8520 15258 8544 15260
rect 8600 15258 8624 15260
rect 8680 15258 8686 15260
rect 8440 15206 8442 15258
rect 8622 15206 8624 15258
rect 8378 15204 8384 15206
rect 8440 15204 8464 15206
rect 8520 15204 8544 15206
rect 8600 15204 8624 15206
rect 8680 15204 8686 15206
rect 8378 15195 8686 15204
rect 8378 14172 8686 14181
rect 8378 14170 8384 14172
rect 8440 14170 8464 14172
rect 8520 14170 8544 14172
rect 8600 14170 8624 14172
rect 8680 14170 8686 14172
rect 8440 14118 8442 14170
rect 8622 14118 8624 14170
rect 8378 14116 8384 14118
rect 8440 14116 8464 14118
rect 8520 14116 8544 14118
rect 8600 14116 8624 14118
rect 8680 14116 8686 14118
rect 8378 14107 8686 14116
rect 9140 13394 9168 15642
rect 9404 14408 9456 14414
rect 9404 14350 9456 14356
rect 9416 14074 9444 14350
rect 9404 14068 9456 14074
rect 9404 14010 9456 14016
rect 9128 13388 9180 13394
rect 9128 13330 9180 13336
rect 9508 13258 9536 16390
rect 9600 16114 9628 16594
rect 10980 16250 11008 17546
rect 10968 16244 11020 16250
rect 10968 16186 11020 16192
rect 9588 16108 9640 16114
rect 9588 16050 9640 16056
rect 9600 14958 9628 16050
rect 9772 15428 9824 15434
rect 9772 15370 9824 15376
rect 9784 15162 9812 15370
rect 10232 15360 10284 15366
rect 10232 15302 10284 15308
rect 10244 15162 10272 15302
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 10232 15156 10284 15162
rect 10232 15098 10284 15104
rect 9588 14952 9640 14958
rect 9588 14894 9640 14900
rect 10244 14550 10272 15098
rect 10980 14550 11008 16186
rect 11072 15162 11100 17818
rect 11164 16182 11192 18702
rect 11704 18352 11756 18358
rect 11704 18294 11756 18300
rect 11152 16176 11204 16182
rect 11152 16118 11204 16124
rect 11164 15638 11192 16118
rect 11612 16108 11664 16114
rect 11612 16050 11664 16056
rect 11152 15632 11204 15638
rect 11152 15574 11204 15580
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 10232 14544 10284 14550
rect 10232 14486 10284 14492
rect 10968 14544 11020 14550
rect 10968 14486 11020 14492
rect 10692 14476 10744 14482
rect 10692 14418 10744 14424
rect 9220 13252 9272 13258
rect 9220 13194 9272 13200
rect 9496 13252 9548 13258
rect 9496 13194 9548 13200
rect 8378 13084 8686 13093
rect 8378 13082 8384 13084
rect 8440 13082 8464 13084
rect 8520 13082 8544 13084
rect 8600 13082 8624 13084
rect 8680 13082 8686 13084
rect 8440 13030 8442 13082
rect 8622 13030 8624 13082
rect 8378 13028 8384 13030
rect 8440 13028 8464 13030
rect 8520 13028 8544 13030
rect 8600 13028 8624 13030
rect 8680 13028 8686 13030
rect 8378 13019 8686 13028
rect 9232 12986 9260 13194
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9508 12850 9536 13194
rect 9588 13184 9640 13190
rect 9588 13126 9640 13132
rect 9600 12986 9628 13126
rect 9588 12980 9640 12986
rect 9588 12922 9640 12928
rect 9496 12844 9548 12850
rect 9496 12786 9548 12792
rect 8300 12776 8352 12782
rect 8300 12718 8352 12724
rect 9128 12708 9180 12714
rect 9128 12650 9180 12656
rect 7840 12640 7892 12646
rect 7840 12582 7892 12588
rect 7852 12238 7880 12582
rect 7840 12232 7892 12238
rect 7840 12174 7892 12180
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 7932 12164 7984 12170
rect 7932 12106 7984 12112
rect 7944 11898 7972 12106
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 7932 11892 7984 11898
rect 7932 11834 7984 11840
rect 7564 11756 7616 11762
rect 7564 11698 7616 11704
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 5448 11144 5500 11150
rect 5448 11086 5500 11092
rect 5552 10266 5580 11154
rect 5632 11144 5684 11150
rect 5632 11086 5684 11092
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5552 9518 5580 10202
rect 5644 9586 5672 11086
rect 5724 11076 5776 11082
rect 5724 11018 5776 11024
rect 5736 10742 5764 11018
rect 5724 10736 5776 10742
rect 5724 10678 5776 10684
rect 6840 9586 6868 11630
rect 7576 11354 7604 11698
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 7852 10742 7880 11698
rect 8024 11620 8076 11626
rect 8024 11562 8076 11568
rect 8036 11218 8064 11562
rect 8024 11212 8076 11218
rect 8024 11154 8076 11160
rect 8036 10742 8064 11154
rect 8128 10810 8156 12174
rect 8378 11996 8686 12005
rect 8378 11994 8384 11996
rect 8440 11994 8464 11996
rect 8520 11994 8544 11996
rect 8600 11994 8624 11996
rect 8680 11994 8686 11996
rect 8440 11942 8442 11994
rect 8622 11942 8624 11994
rect 8378 11940 8384 11942
rect 8440 11940 8464 11942
rect 8520 11940 8544 11942
rect 8600 11940 8624 11942
rect 8680 11940 8686 11942
rect 8378 11931 8686 11940
rect 8944 11756 8996 11762
rect 8944 11698 8996 11704
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 7840 10736 7892 10742
rect 7840 10678 7892 10684
rect 8024 10736 8076 10742
rect 8024 10678 8076 10684
rect 7656 9920 7708 9926
rect 7656 9862 7708 9868
rect 7668 9654 7696 9862
rect 7656 9648 7708 9654
rect 7656 9590 7708 9596
rect 5632 9580 5684 9586
rect 5632 9522 5684 9528
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 5540 9512 5592 9518
rect 5540 9454 5592 9460
rect 5644 8974 5672 9522
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 5080 6384 5132 6390
rect 5080 6326 5132 6332
rect 5276 6322 5304 7346
rect 5368 6866 5396 8434
rect 5448 8424 5500 8430
rect 5448 8366 5500 8372
rect 5460 7410 5488 8366
rect 5644 7478 5672 8910
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 5736 7954 5764 8230
rect 5724 7948 5776 7954
rect 5724 7890 5776 7896
rect 6092 7812 6144 7818
rect 6092 7754 6144 7760
rect 6104 7546 6132 7754
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 6656 7546 6684 7686
rect 6092 7540 6144 7546
rect 6092 7482 6144 7488
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 5632 7472 5684 7478
rect 5632 7414 5684 7420
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5356 6860 5408 6866
rect 5356 6802 5408 6808
rect 5460 6322 5488 7346
rect 6932 7002 6960 8298
rect 7852 7886 7880 10678
rect 8220 10130 8248 11154
rect 8378 10908 8686 10917
rect 8378 10906 8384 10908
rect 8440 10906 8464 10908
rect 8520 10906 8544 10908
rect 8600 10906 8624 10908
rect 8680 10906 8686 10908
rect 8440 10854 8442 10906
rect 8622 10854 8624 10906
rect 8378 10852 8384 10854
rect 8440 10852 8464 10854
rect 8520 10852 8544 10854
rect 8600 10852 8624 10854
rect 8680 10852 8686 10854
rect 8378 10843 8686 10852
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8300 9920 8352 9926
rect 8300 9862 8352 9868
rect 8312 9722 8340 9862
rect 8378 9820 8686 9829
rect 8378 9818 8384 9820
rect 8440 9818 8464 9820
rect 8520 9818 8544 9820
rect 8600 9818 8624 9820
rect 8680 9818 8686 9820
rect 8440 9766 8442 9818
rect 8622 9766 8624 9818
rect 8378 9764 8384 9766
rect 8440 9764 8464 9766
rect 8520 9764 8544 9766
rect 8600 9764 8624 9766
rect 8680 9764 8686 9766
rect 8378 9755 8686 9764
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 8392 9716 8444 9722
rect 8392 9658 8444 9664
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 8312 8974 8340 9522
rect 8404 9042 8432 9658
rect 8392 9036 8444 9042
rect 8392 8978 8444 8984
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8312 8634 8340 8910
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8378 8732 8686 8741
rect 8378 8730 8384 8732
rect 8440 8730 8464 8732
rect 8520 8730 8544 8732
rect 8600 8730 8624 8732
rect 8680 8730 8686 8732
rect 8440 8678 8442 8730
rect 8622 8678 8624 8730
rect 8378 8676 8384 8678
rect 8440 8676 8464 8678
rect 8520 8676 8544 8678
rect 8600 8676 8624 8678
rect 8680 8676 8686 8678
rect 8378 8667 8686 8676
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8312 8430 8340 8570
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 7748 7744 7800 7750
rect 7748 7686 7800 7692
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 7116 7410 7144 7686
rect 7760 7410 7788 7686
rect 8036 7478 8064 7686
rect 8378 7644 8686 7653
rect 8378 7642 8384 7644
rect 8440 7642 8464 7644
rect 8520 7642 8544 7644
rect 8600 7642 8624 7644
rect 8680 7642 8686 7644
rect 8440 7590 8442 7642
rect 8622 7590 8624 7642
rect 8378 7588 8384 7590
rect 8440 7588 8464 7590
rect 8520 7588 8544 7590
rect 8600 7588 8624 7590
rect 8680 7588 8686 7590
rect 8378 7579 8686 7588
rect 8772 7478 8800 8774
rect 8024 7472 8076 7478
rect 8024 7414 8076 7420
rect 8760 7472 8812 7478
rect 8760 7414 8812 7420
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 8956 6914 8984 11698
rect 9140 11218 9168 12650
rect 9496 11688 9548 11694
rect 9600 11676 9628 12922
rect 10416 12640 10468 12646
rect 10416 12582 10468 12588
rect 9680 11756 9732 11762
rect 9680 11698 9732 11704
rect 9548 11648 9628 11676
rect 9496 11630 9548 11636
rect 9128 11212 9180 11218
rect 9128 11154 9180 11160
rect 9220 10464 9272 10470
rect 9220 10406 9272 10412
rect 9232 9994 9260 10406
rect 9220 9988 9272 9994
rect 9220 9930 9272 9936
rect 9232 8566 9260 9930
rect 9588 9580 9640 9586
rect 9588 9522 9640 9528
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 9312 8968 9364 8974
rect 9312 8910 9364 8916
rect 9220 8560 9272 8566
rect 9220 8502 9272 8508
rect 9324 8498 9352 8910
rect 9508 8906 9536 9454
rect 9496 8900 9548 8906
rect 9496 8842 9548 8848
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 9324 7342 9352 7822
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 8864 6886 8984 6914
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 8760 6792 8812 6798
rect 8864 6780 8892 6886
rect 8812 6752 8892 6780
rect 8760 6734 8812 6740
rect 5908 6724 5960 6730
rect 5908 6666 5960 6672
rect 5920 6458 5948 6666
rect 7208 6458 7236 6734
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 8312 6322 8340 6598
rect 8378 6556 8686 6565
rect 8378 6554 8384 6556
rect 8440 6554 8464 6556
rect 8520 6554 8544 6556
rect 8600 6554 8624 6556
rect 8680 6554 8686 6556
rect 8440 6502 8442 6554
rect 8622 6502 8624 6554
rect 8378 6500 8384 6502
rect 8440 6500 8464 6502
rect 8520 6500 8544 6502
rect 8600 6500 8624 6502
rect 8680 6500 8686 6502
rect 8378 6491 8686 6500
rect 5264 6316 5316 6322
rect 5264 6258 5316 6264
rect 5448 6316 5500 6322
rect 5448 6258 5500 6264
rect 8300 6316 8352 6322
rect 8300 6258 8352 6264
rect 8772 6254 8800 6734
rect 9404 6724 9456 6730
rect 9404 6666 9456 6672
rect 9416 6458 9444 6666
rect 9404 6452 9456 6458
rect 9404 6394 9456 6400
rect 9508 6338 9536 8842
rect 9600 6914 9628 9522
rect 9692 9178 9720 11698
rect 10428 11558 10456 12582
rect 10704 11762 10732 14418
rect 11624 14414 11652 16050
rect 11716 14822 11744 18294
rect 12360 18154 12388 18770
rect 12912 18290 12940 19314
rect 13004 18970 13032 19314
rect 12992 18964 13044 18970
rect 12992 18906 13044 18912
rect 13832 18766 13860 21082
rect 14476 19242 14504 29038
rect 14924 28552 14976 28558
rect 14924 28494 14976 28500
rect 14936 28218 14964 28494
rect 15292 28416 15344 28422
rect 15292 28358 15344 28364
rect 15304 28218 15332 28358
rect 14924 28212 14976 28218
rect 14924 28154 14976 28160
rect 15292 28212 15344 28218
rect 15292 28154 15344 28160
rect 14648 27464 14700 27470
rect 14648 27406 14700 27412
rect 14660 27062 14688 27406
rect 14648 27056 14700 27062
rect 14648 26998 14700 27004
rect 14556 26444 14608 26450
rect 14556 26386 14608 26392
rect 14568 25906 14596 26386
rect 14556 25900 14608 25906
rect 14556 25842 14608 25848
rect 14556 25220 14608 25226
rect 14556 25162 14608 25168
rect 14568 21146 14596 25162
rect 14660 24818 14688 26998
rect 14936 26382 14964 28154
rect 15016 26784 15068 26790
rect 15016 26726 15068 26732
rect 15028 26450 15056 26726
rect 15016 26444 15068 26450
rect 15016 26386 15068 26392
rect 15200 26444 15252 26450
rect 15200 26386 15252 26392
rect 14924 26376 14976 26382
rect 14924 26318 14976 26324
rect 15108 25764 15160 25770
rect 15108 25706 15160 25712
rect 14648 24812 14700 24818
rect 14648 24754 14700 24760
rect 14660 23798 14688 24754
rect 15120 24750 15148 25706
rect 15016 24744 15068 24750
rect 15016 24686 15068 24692
rect 15108 24744 15160 24750
rect 15108 24686 15160 24692
rect 15028 24138 15056 24686
rect 15016 24132 15068 24138
rect 15016 24074 15068 24080
rect 14648 23792 14700 23798
rect 14648 23734 14700 23740
rect 14924 23656 14976 23662
rect 14924 23598 14976 23604
rect 14740 22976 14792 22982
rect 14740 22918 14792 22924
rect 14752 22710 14780 22918
rect 14740 22704 14792 22710
rect 14740 22646 14792 22652
rect 14740 22432 14792 22438
rect 14740 22374 14792 22380
rect 14556 21140 14608 21146
rect 14556 21082 14608 21088
rect 14752 20942 14780 22374
rect 14936 22098 14964 23598
rect 15016 22432 15068 22438
rect 15016 22374 15068 22380
rect 14924 22092 14976 22098
rect 14924 22034 14976 22040
rect 14936 21554 14964 22034
rect 15028 21962 15056 22374
rect 15212 22166 15240 26386
rect 15200 22160 15252 22166
rect 15200 22102 15252 22108
rect 15016 21956 15068 21962
rect 15016 21898 15068 21904
rect 14924 21548 14976 21554
rect 14924 21490 14976 21496
rect 14740 20936 14792 20942
rect 14740 20878 14792 20884
rect 14648 20460 14700 20466
rect 14648 20402 14700 20408
rect 14464 19236 14516 19242
rect 14464 19178 14516 19184
rect 14280 19168 14332 19174
rect 14280 19110 14332 19116
rect 13820 18760 13872 18766
rect 13820 18702 13872 18708
rect 14292 18698 14320 19110
rect 14372 18828 14424 18834
rect 14372 18770 14424 18776
rect 14280 18692 14332 18698
rect 14280 18634 14332 18640
rect 12900 18284 12952 18290
rect 12900 18226 12952 18232
rect 14280 18284 14332 18290
rect 14280 18226 14332 18232
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 11888 18148 11940 18154
rect 11888 18090 11940 18096
rect 12348 18148 12400 18154
rect 12348 18090 12400 18096
rect 11796 17196 11848 17202
rect 11796 17138 11848 17144
rect 11808 16794 11836 17138
rect 11900 16794 11928 18090
rect 11980 18080 12032 18086
rect 11980 18022 12032 18028
rect 11992 17746 12020 18022
rect 12092 17980 12400 17989
rect 12092 17978 12098 17980
rect 12154 17978 12178 17980
rect 12234 17978 12258 17980
rect 12314 17978 12338 17980
rect 12394 17978 12400 17980
rect 12154 17926 12156 17978
rect 12336 17926 12338 17978
rect 12092 17924 12098 17926
rect 12154 17924 12178 17926
rect 12234 17924 12258 17926
rect 12314 17924 12338 17926
rect 12394 17924 12400 17926
rect 12092 17915 12400 17924
rect 12452 17882 12480 18158
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 11980 17740 12032 17746
rect 11980 17682 12032 17688
rect 12912 17678 12940 18226
rect 14292 17882 14320 18226
rect 14280 17876 14332 17882
rect 14280 17818 14332 17824
rect 14384 17814 14412 18770
rect 14372 17808 14424 17814
rect 14372 17750 14424 17756
rect 12440 17672 12492 17678
rect 12440 17614 12492 17620
rect 12900 17672 12952 17678
rect 12900 17614 12952 17620
rect 12452 17270 12480 17614
rect 13820 17332 13872 17338
rect 13820 17274 13872 17280
rect 12440 17264 12492 17270
rect 12440 17206 12492 17212
rect 13084 17060 13136 17066
rect 13084 17002 13136 17008
rect 12092 16892 12400 16901
rect 12092 16890 12098 16892
rect 12154 16890 12178 16892
rect 12234 16890 12258 16892
rect 12314 16890 12338 16892
rect 12394 16890 12400 16892
rect 12154 16838 12156 16890
rect 12336 16838 12338 16890
rect 12092 16836 12098 16838
rect 12154 16836 12178 16838
rect 12234 16836 12258 16838
rect 12314 16836 12338 16838
rect 12394 16836 12400 16838
rect 12092 16827 12400 16836
rect 11796 16788 11848 16794
rect 11796 16730 11848 16736
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 12348 16788 12400 16794
rect 12348 16730 12400 16736
rect 12360 16658 12388 16730
rect 13096 16658 13124 17002
rect 13832 16658 13860 17274
rect 14004 17264 14056 17270
rect 14004 17206 14056 17212
rect 12348 16652 12400 16658
rect 12348 16594 12400 16600
rect 13084 16652 13136 16658
rect 13084 16594 13136 16600
rect 13820 16652 13872 16658
rect 13820 16594 13872 16600
rect 13544 16584 13596 16590
rect 13544 16526 13596 16532
rect 13556 16250 13584 16526
rect 13544 16244 13596 16250
rect 13544 16186 13596 16192
rect 11796 16040 11848 16046
rect 11796 15982 11848 15988
rect 11704 14816 11756 14822
rect 11704 14758 11756 14764
rect 11808 14498 11836 15982
rect 11888 15904 11940 15910
rect 11888 15846 11940 15852
rect 11900 15026 11928 15846
rect 12092 15804 12400 15813
rect 12092 15802 12098 15804
rect 12154 15802 12178 15804
rect 12234 15802 12258 15804
rect 12314 15802 12338 15804
rect 12394 15802 12400 15804
rect 12154 15750 12156 15802
rect 12336 15750 12338 15802
rect 12092 15748 12098 15750
rect 12154 15748 12178 15750
rect 12234 15748 12258 15750
rect 12314 15748 12338 15750
rect 12394 15748 12400 15750
rect 12092 15739 12400 15748
rect 12624 15632 12676 15638
rect 12624 15574 12676 15580
rect 11980 15428 12032 15434
rect 11980 15370 12032 15376
rect 11992 15162 12020 15370
rect 12440 15360 12492 15366
rect 12440 15302 12492 15308
rect 11980 15156 12032 15162
rect 11980 15098 12032 15104
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 11992 14498 12020 15098
rect 12092 14716 12400 14725
rect 12092 14714 12098 14716
rect 12154 14714 12178 14716
rect 12234 14714 12258 14716
rect 12314 14714 12338 14716
rect 12394 14714 12400 14716
rect 12154 14662 12156 14714
rect 12336 14662 12338 14714
rect 12092 14660 12098 14662
rect 12154 14660 12178 14662
rect 12234 14660 12258 14662
rect 12314 14660 12338 14662
rect 12394 14660 12400 14662
rect 12092 14651 12400 14660
rect 11808 14470 11928 14498
rect 11992 14470 12112 14498
rect 11612 14408 11664 14414
rect 11612 14350 11664 14356
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 11520 14272 11572 14278
rect 11520 14214 11572 14220
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 9876 10606 9904 11086
rect 10048 11008 10100 11014
rect 10048 10950 10100 10956
rect 9864 10600 9916 10606
rect 9864 10542 9916 10548
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9784 10130 9812 10406
rect 9876 10266 9904 10542
rect 9864 10260 9916 10266
rect 9864 10202 9916 10208
rect 10060 10130 10088 10950
rect 11532 10742 11560 14214
rect 11808 12238 11836 14350
rect 11900 13938 11928 14470
rect 12084 14346 12112 14470
rect 12452 14414 12480 15302
rect 12440 14408 12492 14414
rect 12440 14350 12492 14356
rect 12072 14340 12124 14346
rect 12072 14282 12124 14288
rect 12440 14272 12492 14278
rect 12440 14214 12492 14220
rect 11888 13932 11940 13938
rect 11888 13874 11940 13880
rect 11900 12782 11928 13874
rect 12092 13628 12400 13637
rect 12092 13626 12098 13628
rect 12154 13626 12178 13628
rect 12234 13626 12258 13628
rect 12314 13626 12338 13628
rect 12394 13626 12400 13628
rect 12154 13574 12156 13626
rect 12336 13574 12338 13626
rect 12092 13572 12098 13574
rect 12154 13572 12178 13574
rect 12234 13572 12258 13574
rect 12314 13572 12338 13574
rect 12394 13572 12400 13574
rect 12092 13563 12400 13572
rect 11888 12776 11940 12782
rect 11888 12718 11940 12724
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 11900 11218 11928 12718
rect 12092 12540 12400 12549
rect 12092 12538 12098 12540
rect 12154 12538 12178 12540
rect 12234 12538 12258 12540
rect 12314 12538 12338 12540
rect 12394 12538 12400 12540
rect 12154 12486 12156 12538
rect 12336 12486 12338 12538
rect 12092 12484 12098 12486
rect 12154 12484 12178 12486
rect 12234 12484 12258 12486
rect 12314 12484 12338 12486
rect 12394 12484 12400 12486
rect 12092 12475 12400 12484
rect 12452 12238 12480 14214
rect 12532 13932 12584 13938
rect 12532 13874 12584 13880
rect 12544 13530 12572 13874
rect 12532 13524 12584 13530
rect 12532 13466 12584 13472
rect 12440 12232 12492 12238
rect 12440 12174 12492 12180
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 11888 11212 11940 11218
rect 11888 11154 11940 11160
rect 11992 10742 12020 11494
rect 12092 11452 12400 11461
rect 12092 11450 12098 11452
rect 12154 11450 12178 11452
rect 12234 11450 12258 11452
rect 12314 11450 12338 11452
rect 12394 11450 12400 11452
rect 12154 11398 12156 11450
rect 12336 11398 12338 11450
rect 12092 11396 12098 11398
rect 12154 11396 12178 11398
rect 12234 11396 12258 11398
rect 12314 11396 12338 11398
rect 12394 11396 12400 11398
rect 12092 11387 12400 11396
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 11520 10736 11572 10742
rect 11520 10678 11572 10684
rect 11980 10736 12032 10742
rect 11980 10678 12032 10684
rect 11152 10668 11204 10674
rect 11152 10610 11204 10616
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 10048 10124 10100 10130
rect 10048 10066 10100 10072
rect 11164 10010 11192 10610
rect 12084 10554 12112 11290
rect 12452 10810 12480 12174
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12440 10804 12492 10810
rect 12440 10746 12492 10752
rect 12544 10690 12572 12038
rect 12636 11898 12664 15574
rect 12716 15564 12768 15570
rect 12716 15506 12768 15512
rect 12808 15564 12860 15570
rect 12808 15506 12860 15512
rect 12624 11892 12676 11898
rect 12624 11834 12676 11840
rect 12624 11552 12676 11558
rect 12624 11494 12676 11500
rect 12636 11150 12664 11494
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12544 10662 12664 10690
rect 11992 10526 12112 10554
rect 12532 10600 12584 10606
rect 12532 10542 12584 10548
rect 11336 10056 11388 10062
rect 11164 10004 11336 10010
rect 11164 9998 11388 10004
rect 11060 9988 11112 9994
rect 11060 9930 11112 9936
rect 11164 9982 11376 9998
rect 11072 9654 11100 9930
rect 11060 9648 11112 9654
rect 11060 9590 11112 9596
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 11164 8498 11192 9982
rect 11992 9518 12020 10526
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12092 10364 12400 10373
rect 12092 10362 12098 10364
rect 12154 10362 12178 10364
rect 12234 10362 12258 10364
rect 12314 10362 12338 10364
rect 12394 10362 12400 10364
rect 12154 10310 12156 10362
rect 12336 10310 12338 10362
rect 12092 10308 12098 10310
rect 12154 10308 12178 10310
rect 12234 10308 12258 10310
rect 12314 10308 12338 10310
rect 12394 10308 12400 10310
rect 12092 10299 12400 10308
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 12084 9586 12112 10202
rect 12072 9580 12124 9586
rect 12072 9522 12124 9528
rect 12452 9518 12480 10406
rect 12544 10266 12572 10542
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 12532 10056 12584 10062
rect 12532 9998 12584 10004
rect 11980 9512 12032 9518
rect 11980 9454 12032 9460
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 12092 9276 12400 9285
rect 12092 9274 12098 9276
rect 12154 9274 12178 9276
rect 12234 9274 12258 9276
rect 12314 9274 12338 9276
rect 12394 9274 12400 9276
rect 12154 9222 12156 9274
rect 12336 9222 12338 9274
rect 12092 9220 12098 9222
rect 12154 9220 12178 9222
rect 12234 9220 12258 9222
rect 12314 9220 12338 9222
rect 12394 9220 12400 9222
rect 12092 9211 12400 9220
rect 12256 8968 12308 8974
rect 12256 8910 12308 8916
rect 12268 8498 12296 8910
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 12256 8492 12308 8498
rect 12256 8434 12308 8440
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 11072 7954 11100 8230
rect 11060 7948 11112 7954
rect 11060 7890 11112 7896
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10796 7546 10824 7822
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 10784 7540 10836 7546
rect 10784 7482 10836 7488
rect 9600 6886 9720 6914
rect 9692 6780 9720 6886
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 9416 6322 9536 6338
rect 9600 6752 9720 6780
rect 9600 6322 9628 6752
rect 9968 6458 9996 6802
rect 10048 6724 10100 6730
rect 10048 6666 10100 6672
rect 10060 6458 10088 6666
rect 11072 6662 11100 7686
rect 11256 7410 11284 8434
rect 12092 8188 12400 8197
rect 12092 8186 12098 8188
rect 12154 8186 12178 8188
rect 12234 8186 12258 8188
rect 12314 8186 12338 8188
rect 12394 8186 12400 8188
rect 12154 8134 12156 8186
rect 12336 8134 12338 8186
rect 12092 8132 12098 8134
rect 12154 8132 12178 8134
rect 12234 8132 12258 8134
rect 12314 8132 12338 8134
rect 12394 8132 12400 8134
rect 12092 8123 12400 8132
rect 12544 8090 12572 9998
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 11704 7812 11756 7818
rect 11704 7754 11756 7760
rect 11716 7546 11744 7754
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 11244 7404 11296 7410
rect 11244 7346 11296 7352
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 12092 7100 12400 7109
rect 12092 7098 12098 7100
rect 12154 7098 12178 7100
rect 12234 7098 12258 7100
rect 12314 7098 12338 7100
rect 12394 7098 12400 7100
rect 12154 7046 12156 7098
rect 12336 7046 12338 7098
rect 12092 7044 12098 7046
rect 12154 7044 12178 7046
rect 12234 7044 12258 7046
rect 12314 7044 12338 7046
rect 12394 7044 12400 7046
rect 12092 7035 12400 7044
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 11980 6384 12032 6390
rect 11980 6326 12032 6332
rect 9404 6316 9536 6322
rect 9456 6310 9536 6316
rect 9588 6316 9640 6322
rect 9404 6258 9456 6264
rect 9588 6258 9640 6264
rect 8760 6248 8812 6254
rect 8760 6190 8812 6196
rect 4664 6012 4972 6021
rect 4664 6010 4670 6012
rect 4726 6010 4750 6012
rect 4806 6010 4830 6012
rect 4886 6010 4910 6012
rect 4966 6010 4972 6012
rect 4726 5958 4728 6010
rect 4908 5958 4910 6010
rect 4664 5956 4670 5958
rect 4726 5956 4750 5958
rect 4806 5956 4830 5958
rect 4886 5956 4910 5958
rect 4966 5956 4972 5958
rect 4664 5947 4972 5956
rect 9416 5710 9444 6258
rect 9600 5778 9628 6258
rect 11992 5778 12020 6326
rect 12092 6012 12400 6021
rect 12092 6010 12098 6012
rect 12154 6010 12178 6012
rect 12234 6010 12258 6012
rect 12314 6010 12338 6012
rect 12394 6010 12400 6012
rect 12154 5958 12156 6010
rect 12336 5958 12338 6010
rect 12092 5956 12098 5958
rect 12154 5956 12178 5958
rect 12234 5956 12258 5958
rect 12314 5956 12338 5958
rect 12394 5956 12400 5958
rect 12092 5947 12400 5956
rect 9588 5772 9640 5778
rect 9588 5714 9640 5720
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 12452 5710 12480 7278
rect 12636 6458 12664 10662
rect 12728 10606 12756 15506
rect 12820 12714 12848 15506
rect 13556 15502 13584 16186
rect 14016 15978 14044 17206
rect 14280 17128 14332 17134
rect 14280 17070 14332 17076
rect 14292 16998 14320 17070
rect 14280 16992 14332 16998
rect 14280 16934 14332 16940
rect 14292 16658 14320 16934
rect 14384 16794 14412 17750
rect 14660 17338 14688 20402
rect 14752 19922 14780 20878
rect 14936 20806 14964 21490
rect 14924 20800 14976 20806
rect 14924 20742 14976 20748
rect 14740 19916 14792 19922
rect 14740 19858 14792 19864
rect 14740 18352 14792 18358
rect 14740 18294 14792 18300
rect 14752 17746 14780 18294
rect 14740 17740 14792 17746
rect 14740 17682 14792 17688
rect 14648 17332 14700 17338
rect 14648 17274 14700 17280
rect 14372 16788 14424 16794
rect 14372 16730 14424 16736
rect 14280 16652 14332 16658
rect 14280 16594 14332 16600
rect 15028 16574 15056 21898
rect 15212 21146 15240 22102
rect 15200 21140 15252 21146
rect 15200 21082 15252 21088
rect 15292 20936 15344 20942
rect 15292 20878 15344 20884
rect 15200 20800 15252 20806
rect 15200 20742 15252 20748
rect 15212 20534 15240 20742
rect 15304 20602 15332 20878
rect 15292 20596 15344 20602
rect 15292 20538 15344 20544
rect 15200 20528 15252 20534
rect 15200 20470 15252 20476
rect 15212 19446 15240 20470
rect 15396 19446 15424 29174
rect 22020 29170 22048 31334
rect 25870 31334 26004 31362
rect 25870 31200 25926 31334
rect 23234 29404 23542 29413
rect 23234 29402 23240 29404
rect 23296 29402 23320 29404
rect 23376 29402 23400 29404
rect 23456 29402 23480 29404
rect 23536 29402 23542 29404
rect 23296 29350 23298 29402
rect 23478 29350 23480 29402
rect 23234 29348 23240 29350
rect 23296 29348 23320 29350
rect 23376 29348 23400 29350
rect 23456 29348 23480 29350
rect 23536 29348 23542 29350
rect 23234 29339 23542 29348
rect 25976 29170 26004 31334
rect 29826 31200 29882 32000
rect 22008 29164 22060 29170
rect 22008 29106 22060 29112
rect 25964 29164 26016 29170
rect 25964 29106 26016 29112
rect 29736 29164 29788 29170
rect 29840 29152 29868 31200
rect 31022 29744 31078 29753
rect 31022 29679 31078 29688
rect 30662 29404 30970 29413
rect 30662 29402 30668 29404
rect 30724 29402 30748 29404
rect 30804 29402 30828 29404
rect 30884 29402 30908 29404
rect 30964 29402 30970 29404
rect 30724 29350 30726 29402
rect 30906 29350 30908 29402
rect 30662 29348 30668 29350
rect 30724 29348 30748 29350
rect 30804 29348 30828 29350
rect 30884 29348 30908 29350
rect 30964 29348 30970 29350
rect 30662 29339 30970 29348
rect 31036 29238 31064 29679
rect 31024 29232 31076 29238
rect 31024 29174 31076 29180
rect 29788 29124 29868 29152
rect 29736 29106 29788 29112
rect 28540 29096 28592 29102
rect 28540 29038 28592 29044
rect 29000 29096 29052 29102
rect 29000 29038 29052 29044
rect 22192 29028 22244 29034
rect 22192 28970 22244 28976
rect 25688 29028 25740 29034
rect 25688 28970 25740 28976
rect 18144 28960 18196 28966
rect 18144 28902 18196 28908
rect 18156 28558 18184 28902
rect 19520 28860 19828 28869
rect 19520 28858 19526 28860
rect 19582 28858 19606 28860
rect 19662 28858 19686 28860
rect 19742 28858 19766 28860
rect 19822 28858 19828 28860
rect 19582 28806 19584 28858
rect 19764 28806 19766 28858
rect 19520 28804 19526 28806
rect 19582 28804 19606 28806
rect 19662 28804 19686 28806
rect 19742 28804 19766 28806
rect 19822 28804 19828 28806
rect 19520 28795 19828 28804
rect 18144 28552 18196 28558
rect 18144 28494 18196 28500
rect 20720 28552 20772 28558
rect 20720 28494 20772 28500
rect 21824 28552 21876 28558
rect 21824 28494 21876 28500
rect 16212 28416 16264 28422
rect 16212 28358 16264 28364
rect 15806 28316 16114 28325
rect 15806 28314 15812 28316
rect 15868 28314 15892 28316
rect 15948 28314 15972 28316
rect 16028 28314 16052 28316
rect 16108 28314 16114 28316
rect 15868 28262 15870 28314
rect 16050 28262 16052 28314
rect 15806 28260 15812 28262
rect 15868 28260 15892 28262
rect 15948 28260 15972 28262
rect 16028 28260 16052 28262
rect 16108 28260 16114 28262
rect 15806 28251 16114 28260
rect 15476 28144 15528 28150
rect 15476 28086 15528 28092
rect 15488 27538 15516 28086
rect 16224 28082 16252 28358
rect 16212 28076 16264 28082
rect 16212 28018 16264 28024
rect 15476 27532 15528 27538
rect 15476 27474 15528 27480
rect 15806 27228 16114 27237
rect 15806 27226 15812 27228
rect 15868 27226 15892 27228
rect 15948 27226 15972 27228
rect 16028 27226 16052 27228
rect 16108 27226 16114 27228
rect 15868 27174 15870 27226
rect 16050 27174 16052 27226
rect 15806 27172 15812 27174
rect 15868 27172 15892 27174
rect 15948 27172 15972 27174
rect 16028 27172 16052 27174
rect 16108 27172 16114 27174
rect 15806 27163 16114 27172
rect 16212 26988 16264 26994
rect 16212 26930 16264 26936
rect 16224 26586 16252 26930
rect 16580 26920 16632 26926
rect 16580 26862 16632 26868
rect 18052 26920 18104 26926
rect 18052 26862 18104 26868
rect 16212 26580 16264 26586
rect 16212 26522 16264 26528
rect 15660 26308 15712 26314
rect 15660 26250 15712 26256
rect 15672 24886 15700 26250
rect 15806 26140 16114 26149
rect 15806 26138 15812 26140
rect 15868 26138 15892 26140
rect 15948 26138 15972 26140
rect 16028 26138 16052 26140
rect 16108 26138 16114 26140
rect 15868 26086 15870 26138
rect 16050 26086 16052 26138
rect 15806 26084 15812 26086
rect 15868 26084 15892 26086
rect 15948 26084 15972 26086
rect 16028 26084 16052 26086
rect 16108 26084 16114 26086
rect 15806 26075 16114 26084
rect 15806 25052 16114 25061
rect 15806 25050 15812 25052
rect 15868 25050 15892 25052
rect 15948 25050 15972 25052
rect 16028 25050 16052 25052
rect 16108 25050 16114 25052
rect 15868 24998 15870 25050
rect 16050 24998 16052 25050
rect 15806 24996 15812 24998
rect 15868 24996 15892 24998
rect 15948 24996 15972 24998
rect 16028 24996 16052 24998
rect 16108 24996 16114 24998
rect 15806 24987 16114 24996
rect 15660 24880 15712 24886
rect 15660 24822 15712 24828
rect 15936 24812 15988 24818
rect 15936 24754 15988 24760
rect 15948 24410 15976 24754
rect 16592 24750 16620 26862
rect 17868 24812 17920 24818
rect 17868 24754 17920 24760
rect 16304 24744 16356 24750
rect 16304 24686 16356 24692
rect 16580 24744 16632 24750
rect 16580 24686 16632 24692
rect 15936 24404 15988 24410
rect 15936 24346 15988 24352
rect 15806 23964 16114 23973
rect 15806 23962 15812 23964
rect 15868 23962 15892 23964
rect 15948 23962 15972 23964
rect 16028 23962 16052 23964
rect 16108 23962 16114 23964
rect 15868 23910 15870 23962
rect 16050 23910 16052 23962
rect 15806 23908 15812 23910
rect 15868 23908 15892 23910
rect 15948 23908 15972 23910
rect 16028 23908 16052 23910
rect 16108 23908 16114 23910
rect 15806 23899 16114 23908
rect 16316 23866 16344 24686
rect 17880 24410 17908 24754
rect 17868 24404 17920 24410
rect 17868 24346 17920 24352
rect 16304 23860 16356 23866
rect 16304 23802 16356 23808
rect 15476 23724 15528 23730
rect 15476 23666 15528 23672
rect 15488 23322 15516 23666
rect 15476 23316 15528 23322
rect 15476 23258 15528 23264
rect 15660 23180 15712 23186
rect 15660 23122 15712 23128
rect 15476 22976 15528 22982
rect 15476 22918 15528 22924
rect 15200 19440 15252 19446
rect 15200 19382 15252 19388
rect 15384 19440 15436 19446
rect 15384 19382 15436 19388
rect 15292 19236 15344 19242
rect 15292 19178 15344 19184
rect 15304 18766 15332 19178
rect 15292 18760 15344 18766
rect 15292 18702 15344 18708
rect 15200 18624 15252 18630
rect 15200 18566 15252 18572
rect 15212 18290 15240 18566
rect 15304 18290 15332 18702
rect 15396 18442 15424 19382
rect 15488 18630 15516 22918
rect 15672 22778 15700 23122
rect 16316 23118 16344 23802
rect 16580 23180 16632 23186
rect 16580 23122 16632 23128
rect 16304 23112 16356 23118
rect 16304 23054 16356 23060
rect 15806 22876 16114 22885
rect 15806 22874 15812 22876
rect 15868 22874 15892 22876
rect 15948 22874 15972 22876
rect 16028 22874 16052 22876
rect 16108 22874 16114 22876
rect 15868 22822 15870 22874
rect 16050 22822 16052 22874
rect 15806 22820 15812 22822
rect 15868 22820 15892 22822
rect 15948 22820 15972 22822
rect 16028 22820 16052 22822
rect 16108 22820 16114 22822
rect 15806 22811 16114 22820
rect 15660 22772 15712 22778
rect 15660 22714 15712 22720
rect 15672 22234 15700 22714
rect 16592 22506 16620 23122
rect 16580 22500 16632 22506
rect 16580 22442 16632 22448
rect 17408 22500 17460 22506
rect 17408 22442 17460 22448
rect 16672 22432 16724 22438
rect 16672 22374 16724 22380
rect 15660 22228 15712 22234
rect 15660 22170 15712 22176
rect 16684 22030 16712 22374
rect 16672 22024 16724 22030
rect 16672 21966 16724 21972
rect 17224 21956 17276 21962
rect 17224 21898 17276 21904
rect 15806 21788 16114 21797
rect 15806 21786 15812 21788
rect 15868 21786 15892 21788
rect 15948 21786 15972 21788
rect 16028 21786 16052 21788
rect 16108 21786 16114 21788
rect 15868 21734 15870 21786
rect 16050 21734 16052 21786
rect 15806 21732 15812 21734
rect 15868 21732 15892 21734
rect 15948 21732 15972 21734
rect 16028 21732 16052 21734
rect 16108 21732 16114 21734
rect 15806 21723 16114 21732
rect 17236 21554 17264 21898
rect 17224 21548 17276 21554
rect 17224 21490 17276 21496
rect 16488 20868 16540 20874
rect 16488 20810 16540 20816
rect 15806 20700 16114 20709
rect 15806 20698 15812 20700
rect 15868 20698 15892 20700
rect 15948 20698 15972 20700
rect 16028 20698 16052 20700
rect 16108 20698 16114 20700
rect 15868 20646 15870 20698
rect 16050 20646 16052 20698
rect 15806 20644 15812 20646
rect 15868 20644 15892 20646
rect 15948 20644 15972 20646
rect 16028 20644 16052 20646
rect 16108 20644 16114 20646
rect 15806 20635 16114 20644
rect 15660 20596 15712 20602
rect 15660 20538 15712 20544
rect 15568 20460 15620 20466
rect 15568 20402 15620 20408
rect 15476 18624 15528 18630
rect 15476 18566 15528 18572
rect 15396 18426 15516 18442
rect 15396 18420 15528 18426
rect 15396 18414 15476 18420
rect 15200 18284 15252 18290
rect 15200 18226 15252 18232
rect 15292 18284 15344 18290
rect 15292 18226 15344 18232
rect 15396 18222 15424 18414
rect 15476 18362 15528 18368
rect 15384 18216 15436 18222
rect 15384 18158 15436 18164
rect 15200 17672 15252 17678
rect 15200 17614 15252 17620
rect 15108 17604 15160 17610
rect 15108 17546 15160 17552
rect 14752 16546 15056 16574
rect 13820 15972 13872 15978
rect 13820 15914 13872 15920
rect 14004 15972 14056 15978
rect 14004 15914 14056 15920
rect 13544 15496 13596 15502
rect 13544 15438 13596 15444
rect 13832 15434 13860 15914
rect 14096 15904 14148 15910
rect 14096 15846 14148 15852
rect 13452 15428 13504 15434
rect 13452 15370 13504 15376
rect 13820 15428 13872 15434
rect 13820 15370 13872 15376
rect 13176 15088 13228 15094
rect 13176 15030 13228 15036
rect 13188 14550 13216 15030
rect 13464 15026 13492 15370
rect 13452 15020 13504 15026
rect 13452 14962 13504 14968
rect 13820 14952 13872 14958
rect 13820 14894 13872 14900
rect 13832 14550 13860 14894
rect 13176 14544 13228 14550
rect 13176 14486 13228 14492
rect 13820 14544 13872 14550
rect 13820 14486 13872 14492
rect 14108 13938 14136 15846
rect 14752 15094 14780 16546
rect 15120 16130 15148 17546
rect 15212 17202 15240 17614
rect 15396 17270 15424 18158
rect 15476 17604 15528 17610
rect 15476 17546 15528 17552
rect 15292 17264 15344 17270
rect 15292 17206 15344 17212
rect 15384 17264 15436 17270
rect 15384 17206 15436 17212
rect 15200 17196 15252 17202
rect 15200 17138 15252 17144
rect 15212 16658 15240 17138
rect 15200 16652 15252 16658
rect 15200 16594 15252 16600
rect 15304 16454 15332 17206
rect 15488 17202 15516 17546
rect 15476 17196 15528 17202
rect 15476 17138 15528 17144
rect 15384 17060 15436 17066
rect 15384 17002 15436 17008
rect 15292 16448 15344 16454
rect 15292 16390 15344 16396
rect 15028 16102 15148 16130
rect 15396 16114 15424 17002
rect 15488 16590 15516 17138
rect 15580 17066 15608 20402
rect 15672 20262 15700 20538
rect 16500 20466 16528 20810
rect 16488 20460 16540 20466
rect 16488 20402 16540 20408
rect 15660 20256 15712 20262
rect 15660 20198 15712 20204
rect 17236 19786 17264 21490
rect 17420 21486 17448 22442
rect 17960 21548 18012 21554
rect 17960 21490 18012 21496
rect 17408 21480 17460 21486
rect 17408 21422 17460 21428
rect 17420 20466 17448 21422
rect 17500 20936 17552 20942
rect 17500 20878 17552 20884
rect 17408 20460 17460 20466
rect 17408 20402 17460 20408
rect 17512 20398 17540 20878
rect 17868 20868 17920 20874
rect 17868 20810 17920 20816
rect 17500 20392 17552 20398
rect 17500 20334 17552 20340
rect 17684 20392 17736 20398
rect 17684 20334 17736 20340
rect 17224 19780 17276 19786
rect 17224 19722 17276 19728
rect 17592 19780 17644 19786
rect 17592 19722 17644 19728
rect 15806 19612 16114 19621
rect 15806 19610 15812 19612
rect 15868 19610 15892 19612
rect 15948 19610 15972 19612
rect 16028 19610 16052 19612
rect 16108 19610 16114 19612
rect 15868 19558 15870 19610
rect 16050 19558 16052 19610
rect 15806 19556 15812 19558
rect 15868 19556 15892 19558
rect 15948 19556 15972 19558
rect 16028 19556 16052 19558
rect 16108 19556 16114 19558
rect 15806 19547 16114 19556
rect 15660 19372 15712 19378
rect 15660 19314 15712 19320
rect 15672 18358 15700 19314
rect 16212 19304 16264 19310
rect 16212 19246 16264 19252
rect 15806 18524 16114 18533
rect 15806 18522 15812 18524
rect 15868 18522 15892 18524
rect 15948 18522 15972 18524
rect 16028 18522 16052 18524
rect 16108 18522 16114 18524
rect 15868 18470 15870 18522
rect 16050 18470 16052 18522
rect 15806 18468 15812 18470
rect 15868 18468 15892 18470
rect 15948 18468 15972 18470
rect 16028 18468 16052 18470
rect 16108 18468 16114 18470
rect 15806 18459 16114 18468
rect 15660 18352 15712 18358
rect 15660 18294 15712 18300
rect 16224 18290 16252 19246
rect 17132 18828 17184 18834
rect 17132 18770 17184 18776
rect 16304 18760 16356 18766
rect 16304 18702 16356 18708
rect 16212 18284 16264 18290
rect 16212 18226 16264 18232
rect 16316 18086 16344 18702
rect 16396 18624 16448 18630
rect 16396 18566 16448 18572
rect 16304 18080 16356 18086
rect 16304 18022 16356 18028
rect 16316 17746 16344 18022
rect 16304 17740 16356 17746
rect 16304 17682 16356 17688
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 15568 17060 15620 17066
rect 15568 17002 15620 17008
rect 15568 16720 15620 16726
rect 15568 16662 15620 16668
rect 15476 16584 15528 16590
rect 15476 16526 15528 16532
rect 15580 16250 15608 16662
rect 15568 16244 15620 16250
rect 15568 16186 15620 16192
rect 15580 16114 15608 16186
rect 15672 16182 15700 17614
rect 15806 17436 16114 17445
rect 15806 17434 15812 17436
rect 15868 17434 15892 17436
rect 15948 17434 15972 17436
rect 16028 17434 16052 17436
rect 16108 17434 16114 17436
rect 15868 17382 15870 17434
rect 16050 17382 16052 17434
rect 15806 17380 15812 17382
rect 15868 17380 15892 17382
rect 15948 17380 15972 17382
rect 16028 17380 16052 17382
rect 16108 17380 16114 17382
rect 15806 17371 16114 17380
rect 16212 17264 16264 17270
rect 16212 17206 16264 17212
rect 16120 17196 16172 17202
rect 16120 17138 16172 17144
rect 15752 17128 15804 17134
rect 15752 17070 15804 17076
rect 15764 16998 15792 17070
rect 15752 16992 15804 16998
rect 15752 16934 15804 16940
rect 16132 16454 16160 17138
rect 16224 16522 16252 17206
rect 16316 17134 16344 17682
rect 16408 17678 16436 18566
rect 17144 18426 17172 18770
rect 17132 18420 17184 18426
rect 17132 18362 17184 18368
rect 16488 18216 16540 18222
rect 16488 18158 16540 18164
rect 16396 17672 16448 17678
rect 16396 17614 16448 17620
rect 16304 17128 16356 17134
rect 16304 17070 16356 17076
rect 16500 16726 16528 18158
rect 16764 17332 16816 17338
rect 16764 17274 16816 17280
rect 16776 17202 16804 17274
rect 16764 17196 16816 17202
rect 16764 17138 16816 17144
rect 16580 17128 16632 17134
rect 16580 17070 16632 17076
rect 16488 16720 16540 16726
rect 16488 16662 16540 16668
rect 16212 16516 16264 16522
rect 16212 16458 16264 16464
rect 16488 16516 16540 16522
rect 16488 16458 16540 16464
rect 16120 16448 16172 16454
rect 16120 16390 16172 16396
rect 15806 16348 16114 16357
rect 15806 16346 15812 16348
rect 15868 16346 15892 16348
rect 15948 16346 15972 16348
rect 16028 16346 16052 16348
rect 16108 16346 16114 16348
rect 15868 16294 15870 16346
rect 16050 16294 16052 16346
rect 15806 16292 15812 16294
rect 15868 16292 15892 16294
rect 15948 16292 15972 16294
rect 16028 16292 16052 16294
rect 16108 16292 16114 16294
rect 15806 16283 16114 16292
rect 15660 16176 15712 16182
rect 15660 16118 15712 16124
rect 16224 16114 16252 16458
rect 15384 16108 15436 16114
rect 14740 15088 14792 15094
rect 14740 15030 14792 15036
rect 14648 14816 14700 14822
rect 14648 14758 14700 14764
rect 14924 14816 14976 14822
rect 14924 14758 14976 14764
rect 14188 14408 14240 14414
rect 14188 14350 14240 14356
rect 14200 14074 14228 14350
rect 14188 14068 14240 14074
rect 14188 14010 14240 14016
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 13176 13728 13228 13734
rect 13176 13670 13228 13676
rect 13188 13394 13216 13670
rect 13176 13388 13228 13394
rect 13176 13330 13228 13336
rect 13268 13388 13320 13394
rect 13268 13330 13320 13336
rect 12808 12708 12860 12714
rect 12808 12650 12860 12656
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 12716 10600 12768 10606
rect 12716 10542 12768 10548
rect 12820 9926 12848 11834
rect 13084 11688 13136 11694
rect 13084 11630 13136 11636
rect 13096 11354 13124 11630
rect 13084 11348 13136 11354
rect 13084 11290 13136 11296
rect 13188 11098 13216 13330
rect 13280 11694 13308 13330
rect 13360 13252 13412 13258
rect 13360 13194 13412 13200
rect 13268 11688 13320 11694
rect 13268 11630 13320 11636
rect 13004 11070 13216 11098
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12912 8634 12940 10610
rect 13004 8906 13032 11070
rect 12992 8900 13044 8906
rect 12992 8842 13044 8848
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 13004 8498 13032 8842
rect 13084 8832 13136 8838
rect 13084 8774 13136 8780
rect 13096 8498 13124 8774
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 13084 8492 13136 8498
rect 13084 8434 13136 8440
rect 13372 7546 13400 13194
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 14292 10266 14320 10610
rect 14556 10464 14608 10470
rect 14556 10406 14608 10412
rect 14280 10260 14332 10266
rect 14280 10202 14332 10208
rect 14568 10130 14596 10406
rect 14556 10124 14608 10130
rect 14556 10066 14608 10072
rect 14660 10062 14688 14758
rect 14936 14482 14964 14758
rect 14924 14476 14976 14482
rect 14924 14418 14976 14424
rect 15028 14328 15056 16102
rect 15384 16050 15436 16056
rect 15568 16108 15620 16114
rect 15568 16050 15620 16056
rect 16212 16108 16264 16114
rect 16212 16050 16264 16056
rect 16500 16046 16528 16458
rect 15108 16040 15160 16046
rect 15108 15982 15160 15988
rect 16488 16040 16540 16046
rect 16488 15982 16540 15988
rect 14936 14300 15056 14328
rect 14936 13938 14964 14300
rect 14924 13932 14976 13938
rect 14924 13874 14976 13880
rect 14936 12850 14964 13874
rect 15120 13394 15148 15982
rect 15384 15632 15436 15638
rect 15384 15574 15436 15580
rect 15200 14952 15252 14958
rect 15200 14894 15252 14900
rect 15108 13388 15160 13394
rect 15108 13330 15160 13336
rect 14924 12844 14976 12850
rect 14924 12786 14976 12792
rect 14936 11082 14964 12786
rect 15120 12714 15148 13330
rect 15108 12708 15160 12714
rect 15108 12650 15160 12656
rect 14924 11076 14976 11082
rect 14924 11018 14976 11024
rect 15120 10130 15148 12650
rect 15108 10124 15160 10130
rect 15108 10066 15160 10072
rect 14648 10056 14700 10062
rect 14648 9998 14700 10004
rect 14660 9722 14688 9998
rect 14648 9716 14700 9722
rect 14648 9658 14700 9664
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14476 9178 14504 9454
rect 14832 9376 14884 9382
rect 14832 9318 14884 9324
rect 14464 9172 14516 9178
rect 14464 9114 14516 9120
rect 14476 8498 14504 9114
rect 14844 8974 14872 9318
rect 14832 8968 14884 8974
rect 14832 8910 14884 8916
rect 13452 8492 13504 8498
rect 13452 8434 13504 8440
rect 13912 8492 13964 8498
rect 13912 8434 13964 8440
rect 14464 8492 14516 8498
rect 14464 8434 14516 8440
rect 13464 8090 13492 8434
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 13924 7818 13952 8434
rect 14476 7886 14504 8434
rect 15212 7886 15240 14894
rect 15396 9518 15424 15574
rect 16500 15502 16528 15982
rect 16592 15638 16620 17070
rect 16776 16658 16804 17138
rect 17040 16720 17092 16726
rect 17040 16662 17092 16668
rect 16764 16652 16816 16658
rect 16764 16594 16816 16600
rect 16580 15632 16632 15638
rect 16580 15574 16632 15580
rect 16212 15496 16264 15502
rect 16212 15438 16264 15444
rect 16488 15496 16540 15502
rect 16488 15438 16540 15444
rect 15806 15260 16114 15269
rect 15806 15258 15812 15260
rect 15868 15258 15892 15260
rect 15948 15258 15972 15260
rect 16028 15258 16052 15260
rect 16108 15258 16114 15260
rect 15868 15206 15870 15258
rect 16050 15206 16052 15258
rect 15806 15204 15812 15206
rect 15868 15204 15892 15206
rect 15948 15204 15972 15206
rect 16028 15204 16052 15206
rect 16108 15204 16114 15206
rect 15806 15195 16114 15204
rect 16224 14822 16252 15438
rect 16856 15428 16908 15434
rect 16856 15370 16908 15376
rect 16868 15162 16896 15370
rect 16856 15156 16908 15162
rect 16856 15098 16908 15104
rect 17052 14958 17080 16662
rect 17132 15088 17184 15094
rect 17132 15030 17184 15036
rect 17040 14952 17092 14958
rect 17040 14894 17092 14900
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 15568 14340 15620 14346
rect 15568 14282 15620 14288
rect 15580 14074 15608 14282
rect 15806 14172 16114 14181
rect 15806 14170 15812 14172
rect 15868 14170 15892 14172
rect 15948 14170 15972 14172
rect 16028 14170 16052 14172
rect 16108 14170 16114 14172
rect 15868 14118 15870 14170
rect 16050 14118 16052 14170
rect 15806 14116 15812 14118
rect 15868 14116 15892 14118
rect 15948 14116 15972 14118
rect 16028 14116 16052 14118
rect 16108 14116 16114 14118
rect 15806 14107 16114 14116
rect 15568 14068 15620 14074
rect 15568 14010 15620 14016
rect 16224 13326 16252 14758
rect 17144 14482 17172 15030
rect 17236 15026 17264 19722
rect 17604 19446 17632 19722
rect 17592 19440 17644 19446
rect 17592 19382 17644 19388
rect 17408 18692 17460 18698
rect 17408 18634 17460 18640
rect 17500 18692 17552 18698
rect 17500 18634 17552 18640
rect 17420 18358 17448 18634
rect 17408 18352 17460 18358
rect 17408 18294 17460 18300
rect 17512 17202 17540 18634
rect 17696 18358 17724 20334
rect 17776 20324 17828 20330
rect 17776 20266 17828 20272
rect 17684 18352 17736 18358
rect 17684 18294 17736 18300
rect 17788 17338 17816 20266
rect 17880 17610 17908 20810
rect 17972 20806 18000 21490
rect 18064 21146 18092 26862
rect 18156 22030 18184 28494
rect 18604 28416 18656 28422
rect 18604 28358 18656 28364
rect 18616 26994 18644 28358
rect 18788 28212 18840 28218
rect 18788 28154 18840 28160
rect 18604 26988 18656 26994
rect 18604 26930 18656 26936
rect 18800 26382 18828 28154
rect 18880 28144 18932 28150
rect 18880 28086 18932 28092
rect 18892 27538 18920 28086
rect 19892 28008 19944 28014
rect 19892 27950 19944 27956
rect 19520 27772 19828 27781
rect 19520 27770 19526 27772
rect 19582 27770 19606 27772
rect 19662 27770 19686 27772
rect 19742 27770 19766 27772
rect 19822 27770 19828 27772
rect 19582 27718 19584 27770
rect 19764 27718 19766 27770
rect 19520 27716 19526 27718
rect 19582 27716 19606 27718
rect 19662 27716 19686 27718
rect 19742 27716 19766 27718
rect 19822 27716 19828 27718
rect 19520 27707 19828 27716
rect 19904 27674 19932 27950
rect 19892 27668 19944 27674
rect 19892 27610 19944 27616
rect 18880 27532 18932 27538
rect 18880 27474 18932 27480
rect 20732 27334 20760 28494
rect 20904 28416 20956 28422
rect 20904 28358 20956 28364
rect 20812 28076 20864 28082
rect 20812 28018 20864 28024
rect 20824 27606 20852 28018
rect 20916 27674 20944 28358
rect 21836 28082 21864 28494
rect 21088 28076 21140 28082
rect 21088 28018 21140 28024
rect 21824 28076 21876 28082
rect 21824 28018 21876 28024
rect 20904 27668 20956 27674
rect 20904 27610 20956 27616
rect 20812 27600 20864 27606
rect 20812 27542 20864 27548
rect 20824 27334 20852 27542
rect 21100 27538 21128 28018
rect 21364 28008 21416 28014
rect 21364 27950 21416 27956
rect 21088 27532 21140 27538
rect 21088 27474 21140 27480
rect 20720 27328 20772 27334
rect 20720 27270 20772 27276
rect 20812 27328 20864 27334
rect 20812 27270 20864 27276
rect 20076 26988 20128 26994
rect 20076 26930 20128 26936
rect 19520 26684 19828 26693
rect 19520 26682 19526 26684
rect 19582 26682 19606 26684
rect 19662 26682 19686 26684
rect 19742 26682 19766 26684
rect 19822 26682 19828 26684
rect 19582 26630 19584 26682
rect 19764 26630 19766 26682
rect 19520 26628 19526 26630
rect 19582 26628 19606 26630
rect 19662 26628 19686 26630
rect 19742 26628 19766 26630
rect 19822 26628 19828 26630
rect 19520 26619 19828 26628
rect 18788 26376 18840 26382
rect 18788 26318 18840 26324
rect 18420 26240 18472 26246
rect 18420 26182 18472 26188
rect 18432 25906 18460 26182
rect 18420 25900 18472 25906
rect 18420 25842 18472 25848
rect 18800 25294 18828 26318
rect 19432 26240 19484 26246
rect 19432 26182 19484 26188
rect 19444 25974 19472 26182
rect 19432 25968 19484 25974
rect 19432 25910 19484 25916
rect 19520 25596 19828 25605
rect 19520 25594 19526 25596
rect 19582 25594 19606 25596
rect 19662 25594 19686 25596
rect 19742 25594 19766 25596
rect 19822 25594 19828 25596
rect 19582 25542 19584 25594
rect 19764 25542 19766 25594
rect 19520 25540 19526 25542
rect 19582 25540 19606 25542
rect 19662 25540 19686 25542
rect 19742 25540 19766 25542
rect 19822 25540 19828 25542
rect 19520 25531 19828 25540
rect 19524 25356 19576 25362
rect 19524 25298 19576 25304
rect 18788 25288 18840 25294
rect 18788 25230 18840 25236
rect 18236 24948 18288 24954
rect 18236 24890 18288 24896
rect 18248 24206 18276 24890
rect 19536 24682 19564 25298
rect 19892 24744 19944 24750
rect 19892 24686 19944 24692
rect 19340 24676 19392 24682
rect 19340 24618 19392 24624
rect 19524 24676 19576 24682
rect 19524 24618 19576 24624
rect 18512 24608 18564 24614
rect 18512 24550 18564 24556
rect 18420 24268 18472 24274
rect 18420 24210 18472 24216
rect 18236 24200 18288 24206
rect 18236 24142 18288 24148
rect 18432 23526 18460 24210
rect 18524 23730 18552 24550
rect 19352 24206 19380 24618
rect 19520 24508 19828 24517
rect 19520 24506 19526 24508
rect 19582 24506 19606 24508
rect 19662 24506 19686 24508
rect 19742 24506 19766 24508
rect 19822 24506 19828 24508
rect 19582 24454 19584 24506
rect 19764 24454 19766 24506
rect 19520 24452 19526 24454
rect 19582 24452 19606 24454
rect 19662 24452 19686 24454
rect 19742 24452 19766 24454
rect 19822 24452 19828 24454
rect 19520 24443 19828 24452
rect 19904 24274 19932 24686
rect 19892 24268 19944 24274
rect 19892 24210 19944 24216
rect 19984 24268 20036 24274
rect 19984 24210 20036 24216
rect 19340 24200 19392 24206
rect 19340 24142 19392 24148
rect 19432 24064 19484 24070
rect 19432 24006 19484 24012
rect 19444 23798 19472 24006
rect 19904 23866 19932 24210
rect 19892 23860 19944 23866
rect 19892 23802 19944 23808
rect 19432 23792 19484 23798
rect 19432 23734 19484 23740
rect 18512 23724 18564 23730
rect 18512 23666 18564 23672
rect 18420 23520 18472 23526
rect 18420 23462 18472 23468
rect 18144 22024 18196 22030
rect 18144 21966 18196 21972
rect 18432 21622 18460 23462
rect 18524 22642 18552 23666
rect 19996 23526 20024 24210
rect 19984 23520 20036 23526
rect 19984 23462 20036 23468
rect 19520 23420 19828 23429
rect 19520 23418 19526 23420
rect 19582 23418 19606 23420
rect 19662 23418 19686 23420
rect 19742 23418 19766 23420
rect 19822 23418 19828 23420
rect 19582 23366 19584 23418
rect 19764 23366 19766 23418
rect 19520 23364 19526 23366
rect 19582 23364 19606 23366
rect 19662 23364 19686 23366
rect 19742 23364 19766 23366
rect 19822 23364 19828 23366
rect 19520 23355 19828 23364
rect 19996 23186 20024 23462
rect 19984 23180 20036 23186
rect 19984 23122 20036 23128
rect 20088 22982 20116 26930
rect 20444 25832 20496 25838
rect 20444 25774 20496 25780
rect 20456 24818 20484 25774
rect 20444 24812 20496 24818
rect 20444 24754 20496 24760
rect 20352 24608 20404 24614
rect 20352 24550 20404 24556
rect 20168 24064 20220 24070
rect 20168 24006 20220 24012
rect 19432 22976 19484 22982
rect 19432 22918 19484 22924
rect 20076 22976 20128 22982
rect 20076 22918 20128 22924
rect 19444 22710 19472 22918
rect 20180 22778 20208 24006
rect 20364 23594 20392 24550
rect 20732 23730 20760 27270
rect 20824 26450 20852 27270
rect 20812 26444 20864 26450
rect 20812 26386 20864 26392
rect 20720 23724 20772 23730
rect 20720 23666 20772 23672
rect 20352 23588 20404 23594
rect 20352 23530 20404 23536
rect 20168 22772 20220 22778
rect 20168 22714 20220 22720
rect 19432 22704 19484 22710
rect 19432 22646 19484 22652
rect 18512 22636 18564 22642
rect 18512 22578 18564 22584
rect 18524 22098 18552 22578
rect 20352 22500 20404 22506
rect 20352 22442 20404 22448
rect 19520 22332 19828 22341
rect 19520 22330 19526 22332
rect 19582 22330 19606 22332
rect 19662 22330 19686 22332
rect 19742 22330 19766 22332
rect 19822 22330 19828 22332
rect 19582 22278 19584 22330
rect 19764 22278 19766 22330
rect 19520 22276 19526 22278
rect 19582 22276 19606 22278
rect 19662 22276 19686 22278
rect 19742 22276 19766 22278
rect 19822 22276 19828 22278
rect 19520 22267 19828 22276
rect 18512 22092 18564 22098
rect 18512 22034 18564 22040
rect 18420 21616 18472 21622
rect 18420 21558 18472 21564
rect 18328 21548 18380 21554
rect 18328 21490 18380 21496
rect 18052 21140 18104 21146
rect 18052 21082 18104 21088
rect 17960 20800 18012 20806
rect 17960 20742 18012 20748
rect 17868 17604 17920 17610
rect 17868 17546 17920 17552
rect 17776 17332 17828 17338
rect 17776 17274 17828 17280
rect 17500 17196 17552 17202
rect 17500 17138 17552 17144
rect 17880 16590 17908 17546
rect 17972 17542 18000 20742
rect 18340 20262 18368 21490
rect 18524 21434 18552 22034
rect 18432 21406 18552 21434
rect 18432 20534 18460 21406
rect 20168 21344 20220 21350
rect 20168 21286 20220 21292
rect 19520 21244 19828 21253
rect 19520 21242 19526 21244
rect 19582 21242 19606 21244
rect 19662 21242 19686 21244
rect 19742 21242 19766 21244
rect 19822 21242 19828 21244
rect 19582 21190 19584 21242
rect 19764 21190 19766 21242
rect 19520 21188 19526 21190
rect 19582 21188 19606 21190
rect 19662 21188 19686 21190
rect 19742 21188 19766 21190
rect 19822 21188 19828 21190
rect 19520 21179 19828 21188
rect 20180 21078 20208 21286
rect 20168 21072 20220 21078
rect 20168 21014 20220 21020
rect 18788 20936 18840 20942
rect 18788 20878 18840 20884
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19984 20936 20036 20942
rect 19984 20878 20036 20884
rect 18800 20602 18828 20878
rect 18788 20596 18840 20602
rect 18788 20538 18840 20544
rect 18420 20528 18472 20534
rect 18420 20470 18472 20476
rect 18328 20256 18380 20262
rect 18328 20198 18380 20204
rect 18340 19854 18368 20198
rect 18512 20052 18564 20058
rect 18512 19994 18564 20000
rect 18328 19848 18380 19854
rect 18328 19790 18380 19796
rect 18052 18692 18104 18698
rect 18052 18634 18104 18640
rect 18064 18426 18092 18634
rect 18340 18630 18368 19790
rect 18420 19780 18472 19786
rect 18420 19722 18472 19728
rect 18432 19514 18460 19722
rect 18420 19508 18472 19514
rect 18420 19450 18472 19456
rect 18524 19378 18552 19994
rect 18972 19916 19024 19922
rect 18972 19858 19024 19864
rect 18512 19372 18564 19378
rect 18512 19314 18564 19320
rect 18420 18760 18472 18766
rect 18420 18702 18472 18708
rect 18328 18624 18380 18630
rect 18328 18566 18380 18572
rect 18052 18420 18104 18426
rect 18052 18362 18104 18368
rect 18328 18352 18380 18358
rect 18328 18294 18380 18300
rect 18236 18216 18288 18222
rect 18236 18158 18288 18164
rect 18144 17604 18196 17610
rect 18144 17546 18196 17552
rect 17960 17536 18012 17542
rect 17960 17478 18012 17484
rect 17972 16726 18000 17478
rect 18156 17270 18184 17546
rect 18144 17264 18196 17270
rect 18144 17206 18196 17212
rect 18248 17202 18276 18158
rect 18340 17202 18368 18294
rect 18432 17678 18460 18702
rect 18984 18290 19012 19858
rect 19444 19854 19472 20878
rect 19996 20466 20024 20878
rect 19984 20460 20036 20466
rect 19984 20402 20036 20408
rect 19892 20392 19944 20398
rect 19892 20334 19944 20340
rect 19520 20156 19828 20165
rect 19520 20154 19526 20156
rect 19582 20154 19606 20156
rect 19662 20154 19686 20156
rect 19742 20154 19766 20156
rect 19822 20154 19828 20156
rect 19582 20102 19584 20154
rect 19764 20102 19766 20154
rect 19520 20100 19526 20102
rect 19582 20100 19606 20102
rect 19662 20100 19686 20102
rect 19742 20100 19766 20102
rect 19822 20100 19828 20102
rect 19520 20091 19828 20100
rect 19432 19848 19484 19854
rect 19432 19790 19484 19796
rect 19520 19068 19828 19077
rect 19520 19066 19526 19068
rect 19582 19066 19606 19068
rect 19662 19066 19686 19068
rect 19742 19066 19766 19068
rect 19822 19066 19828 19068
rect 19582 19014 19584 19066
rect 19764 19014 19766 19066
rect 19520 19012 19526 19014
rect 19582 19012 19606 19014
rect 19662 19012 19686 19014
rect 19742 19012 19766 19014
rect 19822 19012 19828 19014
rect 19520 19003 19828 19012
rect 19904 18766 19932 20334
rect 20364 19922 20392 22442
rect 20824 22098 20852 26386
rect 21100 26382 21128 27474
rect 21376 27402 21404 27950
rect 21364 27396 21416 27402
rect 21364 27338 21416 27344
rect 21088 26376 21140 26382
rect 21088 26318 21140 26324
rect 21824 26376 21876 26382
rect 21824 26318 21876 26324
rect 20904 23656 20956 23662
rect 20904 23598 20956 23604
rect 20916 23118 20944 23598
rect 21100 23322 21128 26318
rect 21836 24750 21864 26318
rect 22204 26246 22232 28970
rect 22836 28552 22888 28558
rect 22836 28494 22888 28500
rect 22376 28416 22428 28422
rect 22376 28358 22428 28364
rect 22388 27538 22416 28358
rect 22744 28008 22796 28014
rect 22744 27950 22796 27956
rect 22756 27674 22784 27950
rect 22744 27668 22796 27674
rect 22744 27610 22796 27616
rect 22376 27532 22428 27538
rect 22376 27474 22428 27480
rect 22284 26308 22336 26314
rect 22284 26250 22336 26256
rect 22008 26240 22060 26246
rect 22008 26182 22060 26188
rect 22192 26240 22244 26246
rect 22192 26182 22244 26188
rect 22020 25906 22048 26182
rect 22008 25900 22060 25906
rect 22008 25842 22060 25848
rect 22204 24954 22232 26182
rect 22296 26042 22324 26250
rect 22284 26036 22336 26042
rect 22284 25978 22336 25984
rect 22652 25764 22704 25770
rect 22652 25706 22704 25712
rect 22664 25362 22692 25706
rect 22652 25356 22704 25362
rect 22652 25298 22704 25304
rect 22192 24948 22244 24954
rect 22192 24890 22244 24896
rect 22192 24812 22244 24818
rect 22192 24754 22244 24760
rect 21364 24744 21416 24750
rect 21364 24686 21416 24692
rect 21824 24744 21876 24750
rect 21824 24686 21876 24692
rect 21376 24274 21404 24686
rect 21364 24268 21416 24274
rect 21364 24210 21416 24216
rect 22008 24132 22060 24138
rect 22008 24074 22060 24080
rect 22020 23866 22048 24074
rect 22008 23860 22060 23866
rect 22008 23802 22060 23808
rect 21088 23316 21140 23322
rect 21088 23258 21140 23264
rect 20904 23112 20956 23118
rect 20904 23054 20956 23060
rect 20916 22778 20944 23054
rect 20904 22772 20956 22778
rect 20904 22714 20956 22720
rect 20812 22092 20864 22098
rect 20812 22034 20864 22040
rect 20824 20466 20852 22034
rect 20904 20936 20956 20942
rect 20904 20878 20956 20884
rect 20916 20602 20944 20878
rect 20904 20596 20956 20602
rect 20904 20538 20956 20544
rect 21100 20466 21128 23258
rect 21456 23044 21508 23050
rect 21456 22986 21508 22992
rect 21272 22976 21324 22982
rect 21272 22918 21324 22924
rect 21180 22024 21232 22030
rect 21180 21966 21232 21972
rect 20812 20460 20864 20466
rect 20812 20402 20864 20408
rect 21088 20460 21140 20466
rect 21088 20402 21140 20408
rect 20352 19916 20404 19922
rect 20352 19858 20404 19864
rect 19432 18760 19484 18766
rect 19432 18702 19484 18708
rect 19892 18760 19944 18766
rect 19892 18702 19944 18708
rect 20996 18760 21048 18766
rect 20996 18702 21048 18708
rect 18972 18284 19024 18290
rect 18972 18226 19024 18232
rect 18420 17672 18472 17678
rect 18420 17614 18472 17620
rect 19444 17338 19472 18702
rect 20628 18624 20680 18630
rect 20628 18566 20680 18572
rect 20640 18358 20668 18566
rect 20628 18352 20680 18358
rect 20628 18294 20680 18300
rect 21008 18086 21036 18702
rect 20076 18080 20128 18086
rect 20076 18022 20128 18028
rect 20996 18080 21048 18086
rect 20996 18022 21048 18028
rect 19520 17980 19828 17989
rect 19520 17978 19526 17980
rect 19582 17978 19606 17980
rect 19662 17978 19686 17980
rect 19742 17978 19766 17980
rect 19822 17978 19828 17980
rect 19582 17926 19584 17978
rect 19764 17926 19766 17978
rect 19520 17924 19526 17926
rect 19582 17924 19606 17926
rect 19662 17924 19686 17926
rect 19742 17924 19766 17926
rect 19822 17924 19828 17926
rect 19520 17915 19828 17924
rect 20088 17746 20116 18022
rect 20076 17740 20128 17746
rect 20076 17682 20128 17688
rect 19432 17332 19484 17338
rect 19432 17274 19484 17280
rect 18236 17196 18288 17202
rect 18236 17138 18288 17144
rect 18328 17196 18380 17202
rect 18328 17138 18380 17144
rect 21008 17134 21036 18022
rect 19432 17128 19484 17134
rect 19432 17070 19484 17076
rect 20996 17128 21048 17134
rect 20996 17070 21048 17076
rect 18420 17060 18472 17066
rect 18420 17002 18472 17008
rect 18052 16992 18104 16998
rect 18052 16934 18104 16940
rect 17960 16720 18012 16726
rect 17960 16662 18012 16668
rect 17868 16584 17920 16590
rect 17868 16526 17920 16532
rect 18064 16454 18092 16934
rect 18432 16794 18460 17002
rect 18420 16788 18472 16794
rect 18420 16730 18472 16736
rect 19444 16658 19472 17070
rect 19520 16892 19828 16901
rect 19520 16890 19526 16892
rect 19582 16890 19606 16892
rect 19662 16890 19686 16892
rect 19742 16890 19766 16892
rect 19822 16890 19828 16892
rect 19582 16838 19584 16890
rect 19764 16838 19766 16890
rect 19520 16836 19526 16838
rect 19582 16836 19606 16838
rect 19662 16836 19686 16838
rect 19742 16836 19766 16838
rect 19822 16836 19828 16838
rect 19520 16827 19828 16836
rect 19432 16652 19484 16658
rect 19432 16594 19484 16600
rect 19984 16652 20036 16658
rect 19984 16594 20036 16600
rect 18052 16448 18104 16454
rect 18052 16390 18104 16396
rect 19432 16448 19484 16454
rect 19432 16390 19484 16396
rect 19524 16448 19576 16454
rect 19524 16390 19576 16396
rect 19892 16448 19944 16454
rect 19892 16390 19944 16396
rect 19444 16182 19472 16390
rect 19432 16176 19484 16182
rect 19432 16118 19484 16124
rect 19536 15994 19564 16390
rect 19444 15966 19564 15994
rect 18604 15496 18656 15502
rect 18604 15438 18656 15444
rect 18616 15366 18644 15438
rect 18788 15428 18840 15434
rect 18788 15370 18840 15376
rect 18604 15360 18656 15366
rect 18604 15302 18656 15308
rect 18616 15094 18644 15302
rect 18604 15088 18656 15094
rect 18604 15030 18656 15036
rect 18800 15026 18828 15370
rect 17224 15020 17276 15026
rect 17224 14962 17276 14968
rect 17500 15020 17552 15026
rect 17500 14962 17552 14968
rect 18788 15020 18840 15026
rect 18788 14962 18840 14968
rect 17408 14952 17460 14958
rect 17408 14894 17460 14900
rect 17224 14816 17276 14822
rect 17224 14758 17276 14764
rect 17132 14476 17184 14482
rect 17132 14418 17184 14424
rect 16764 14340 16816 14346
rect 16764 14282 16816 14288
rect 16304 14272 16356 14278
rect 16304 14214 16356 14220
rect 16488 14272 16540 14278
rect 16488 14214 16540 14220
rect 16316 14074 16344 14214
rect 16304 14068 16356 14074
rect 16304 14010 16356 14016
rect 16396 14068 16448 14074
rect 16396 14010 16448 14016
rect 16212 13320 16264 13326
rect 16212 13262 16264 13268
rect 15806 13084 16114 13093
rect 15806 13082 15812 13084
rect 15868 13082 15892 13084
rect 15948 13082 15972 13084
rect 16028 13082 16052 13084
rect 16108 13082 16114 13084
rect 15868 13030 15870 13082
rect 16050 13030 16052 13082
rect 15806 13028 15812 13030
rect 15868 13028 15892 13030
rect 15948 13028 15972 13030
rect 16028 13028 16052 13030
rect 16108 13028 16114 13030
rect 15806 13019 16114 13028
rect 16224 12170 16252 13262
rect 16408 12238 16436 14010
rect 16500 13938 16528 14214
rect 16488 13932 16540 13938
rect 16488 13874 16540 13880
rect 16396 12232 16448 12238
rect 16396 12174 16448 12180
rect 16212 12164 16264 12170
rect 16212 12106 16264 12112
rect 15806 11996 16114 12005
rect 15806 11994 15812 11996
rect 15868 11994 15892 11996
rect 15948 11994 15972 11996
rect 16028 11994 16052 11996
rect 16108 11994 16114 11996
rect 15868 11942 15870 11994
rect 16050 11942 16052 11994
rect 15806 11940 15812 11942
rect 15868 11940 15892 11942
rect 15948 11940 15972 11942
rect 16028 11940 16052 11942
rect 16108 11940 16114 11942
rect 15806 11931 16114 11940
rect 15806 10908 16114 10917
rect 15806 10906 15812 10908
rect 15868 10906 15892 10908
rect 15948 10906 15972 10908
rect 16028 10906 16052 10908
rect 16108 10906 16114 10908
rect 15868 10854 15870 10906
rect 16050 10854 16052 10906
rect 15806 10852 15812 10854
rect 15868 10852 15892 10854
rect 15948 10852 15972 10854
rect 16028 10852 16052 10854
rect 16108 10852 16114 10854
rect 15806 10843 16114 10852
rect 15806 9820 16114 9829
rect 15806 9818 15812 9820
rect 15868 9818 15892 9820
rect 15948 9818 15972 9820
rect 16028 9818 16052 9820
rect 16108 9818 16114 9820
rect 15868 9766 15870 9818
rect 16050 9766 16052 9818
rect 15806 9764 15812 9766
rect 15868 9764 15892 9766
rect 15948 9764 15972 9766
rect 16028 9764 16052 9766
rect 16108 9764 16114 9766
rect 15806 9755 16114 9764
rect 15384 9512 15436 9518
rect 15384 9454 15436 9460
rect 16224 8974 16252 12106
rect 16304 11008 16356 11014
rect 16304 10950 16356 10956
rect 16316 10674 16344 10950
rect 16776 10674 16804 14282
rect 17236 14074 17264 14758
rect 17224 14068 17276 14074
rect 17224 14010 17276 14016
rect 17420 13870 17448 14894
rect 17512 13938 17540 14962
rect 18604 14952 18656 14958
rect 18604 14894 18656 14900
rect 18512 14612 18564 14618
rect 18512 14554 18564 14560
rect 17500 13932 17552 13938
rect 17500 13874 17552 13880
rect 17316 13864 17368 13870
rect 17316 13806 17368 13812
rect 17408 13864 17460 13870
rect 17408 13806 17460 13812
rect 17328 13394 17356 13806
rect 17316 13388 17368 13394
rect 17316 13330 17368 13336
rect 16856 13252 16908 13258
rect 16856 13194 16908 13200
rect 16868 12986 16896 13194
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 17328 12442 17356 13330
rect 17420 12782 17448 13806
rect 17512 13190 17540 13874
rect 18236 13320 18288 13326
rect 18236 13262 18288 13268
rect 17500 13184 17552 13190
rect 17500 13126 17552 13132
rect 17592 13184 17644 13190
rect 17592 13126 17644 13132
rect 17604 12850 17632 13126
rect 17592 12844 17644 12850
rect 17592 12786 17644 12792
rect 17408 12776 17460 12782
rect 17408 12718 17460 12724
rect 17776 12708 17828 12714
rect 17776 12650 17828 12656
rect 17316 12436 17368 12442
rect 17316 12378 17368 12384
rect 17316 12096 17368 12102
rect 17316 12038 17368 12044
rect 17328 11218 17356 12038
rect 17788 11762 17816 12650
rect 18248 12238 18276 13262
rect 18236 12232 18288 12238
rect 18236 12174 18288 12180
rect 18248 11830 18276 12174
rect 18236 11824 18288 11830
rect 18236 11766 18288 11772
rect 17776 11756 17828 11762
rect 17776 11698 17828 11704
rect 17868 11688 17920 11694
rect 17868 11630 17920 11636
rect 17316 11212 17368 11218
rect 17316 11154 17368 11160
rect 16304 10668 16356 10674
rect 16304 10610 16356 10616
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 16396 9580 16448 9586
rect 16396 9522 16448 9528
rect 16580 9580 16632 9586
rect 16580 9522 16632 9528
rect 16212 8968 16264 8974
rect 16212 8910 16264 8916
rect 15806 8732 16114 8741
rect 15806 8730 15812 8732
rect 15868 8730 15892 8732
rect 15948 8730 15972 8732
rect 16028 8730 16052 8732
rect 16108 8730 16114 8732
rect 15868 8678 15870 8730
rect 16050 8678 16052 8730
rect 15806 8676 15812 8678
rect 15868 8676 15892 8678
rect 15948 8676 15972 8678
rect 16028 8676 16052 8678
rect 16108 8676 16114 8678
rect 15806 8667 16114 8676
rect 14464 7880 14516 7886
rect 14464 7822 14516 7828
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 13912 7812 13964 7818
rect 13912 7754 13964 7760
rect 15806 7644 16114 7653
rect 15806 7642 15812 7644
rect 15868 7642 15892 7644
rect 15948 7642 15972 7644
rect 16028 7642 16052 7644
rect 16108 7642 16114 7644
rect 15868 7590 15870 7642
rect 16050 7590 16052 7642
rect 15806 7588 15812 7590
rect 15868 7588 15892 7590
rect 15948 7588 15972 7590
rect 16028 7588 16052 7590
rect 16108 7588 16114 7590
rect 15806 7579 16114 7588
rect 13360 7540 13412 7546
rect 13360 7482 13412 7488
rect 16224 7342 16252 8910
rect 16408 7546 16436 9522
rect 16592 8514 16620 9522
rect 16500 8486 16620 8514
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16212 7336 16264 7342
rect 16212 7278 16264 7284
rect 14648 6792 14700 6798
rect 14648 6734 14700 6740
rect 13544 6656 13596 6662
rect 13544 6598 13596 6604
rect 14372 6656 14424 6662
rect 14372 6598 14424 6604
rect 12624 6452 12676 6458
rect 12624 6394 12676 6400
rect 13556 6322 13584 6598
rect 13544 6316 13596 6322
rect 13544 6258 13596 6264
rect 9404 5704 9456 5710
rect 9404 5646 9456 5652
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 8378 5468 8686 5477
rect 8378 5466 8384 5468
rect 8440 5466 8464 5468
rect 8520 5466 8544 5468
rect 8600 5466 8624 5468
rect 8680 5466 8686 5468
rect 8440 5414 8442 5466
rect 8622 5414 8624 5466
rect 8378 5412 8384 5414
rect 8440 5412 8464 5414
rect 8520 5412 8544 5414
rect 8600 5412 8624 5414
rect 8680 5412 8686 5414
rect 8378 5403 8686 5412
rect 14384 5166 14412 6598
rect 14660 5914 14688 6734
rect 16500 6730 16528 8486
rect 16672 8288 16724 8294
rect 16672 8230 16724 8236
rect 16684 8090 16712 8230
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 16776 7410 16804 10610
rect 17880 10606 17908 11630
rect 18248 11354 18276 11766
rect 18524 11762 18552 14554
rect 18512 11756 18564 11762
rect 18512 11698 18564 11704
rect 18236 11348 18288 11354
rect 18236 11290 18288 11296
rect 17960 11076 18012 11082
rect 17960 11018 18012 11024
rect 17868 10600 17920 10606
rect 17868 10542 17920 10548
rect 17880 10266 17908 10542
rect 17868 10260 17920 10266
rect 17868 10202 17920 10208
rect 17972 10130 18000 11018
rect 18616 11014 18644 14894
rect 19444 12714 19472 15966
rect 19904 15910 19932 16390
rect 19892 15904 19944 15910
rect 19892 15846 19944 15852
rect 19520 15804 19828 15813
rect 19520 15802 19526 15804
rect 19582 15802 19606 15804
rect 19662 15802 19686 15804
rect 19742 15802 19766 15804
rect 19822 15802 19828 15804
rect 19582 15750 19584 15802
rect 19764 15750 19766 15802
rect 19520 15748 19526 15750
rect 19582 15748 19606 15750
rect 19662 15748 19686 15750
rect 19742 15748 19766 15750
rect 19822 15748 19828 15750
rect 19520 15739 19828 15748
rect 19904 14958 19932 15846
rect 19996 15638 20024 16594
rect 21192 16574 21220 21966
rect 21284 20874 21312 22918
rect 21468 22778 21496 22986
rect 21456 22772 21508 22778
rect 21456 22714 21508 22720
rect 22100 22432 22152 22438
rect 22100 22374 22152 22380
rect 22112 21622 22140 22374
rect 22100 21616 22152 21622
rect 22100 21558 22152 21564
rect 22204 21146 22232 24754
rect 22376 24064 22428 24070
rect 22376 24006 22428 24012
rect 22388 23730 22416 24006
rect 22376 23724 22428 23730
rect 22428 23684 22508 23712
rect 22376 23666 22428 23672
rect 22376 22976 22428 22982
rect 22376 22918 22428 22924
rect 22388 22778 22416 22918
rect 22376 22772 22428 22778
rect 22376 22714 22428 22720
rect 22284 22704 22336 22710
rect 22284 22646 22336 22652
rect 22296 22574 22324 22646
rect 22284 22568 22336 22574
rect 22284 22510 22336 22516
rect 22192 21140 22244 21146
rect 22192 21082 22244 21088
rect 21272 20868 21324 20874
rect 21272 20810 21324 20816
rect 22192 20868 22244 20874
rect 22192 20810 22244 20816
rect 21364 20392 21416 20398
rect 21364 20334 21416 20340
rect 21376 19786 21404 20334
rect 22100 20256 22152 20262
rect 22100 20198 22152 20204
rect 22112 19922 22140 20198
rect 22100 19916 22152 19922
rect 22100 19858 22152 19864
rect 21364 19780 21416 19786
rect 21364 19722 21416 19728
rect 22008 19780 22060 19786
rect 22008 19722 22060 19728
rect 22020 19446 22048 19722
rect 22008 19440 22060 19446
rect 22008 19382 22060 19388
rect 22204 18426 22232 20810
rect 22376 20800 22428 20806
rect 22376 20742 22428 20748
rect 22388 20466 22416 20742
rect 22376 20460 22428 20466
rect 22376 20402 22428 20408
rect 22388 19990 22416 20402
rect 22376 19984 22428 19990
rect 22376 19926 22428 19932
rect 22480 18630 22508 23684
rect 22664 23662 22692 25298
rect 22744 25288 22796 25294
rect 22744 25230 22796 25236
rect 22756 24410 22784 25230
rect 22744 24404 22796 24410
rect 22744 24346 22796 24352
rect 22756 24138 22784 24346
rect 22744 24132 22796 24138
rect 22744 24074 22796 24080
rect 22756 23866 22784 24074
rect 22744 23860 22796 23866
rect 22744 23802 22796 23808
rect 22652 23656 22704 23662
rect 22652 23598 22704 23604
rect 22664 21350 22692 23598
rect 22848 22030 22876 28494
rect 23572 28484 23624 28490
rect 23572 28426 23624 28432
rect 23234 28316 23542 28325
rect 23234 28314 23240 28316
rect 23296 28314 23320 28316
rect 23376 28314 23400 28316
rect 23456 28314 23480 28316
rect 23536 28314 23542 28316
rect 23296 28262 23298 28314
rect 23478 28262 23480 28314
rect 23234 28260 23240 28262
rect 23296 28260 23320 28262
rect 23376 28260 23400 28262
rect 23456 28260 23480 28262
rect 23536 28260 23542 28262
rect 23234 28251 23542 28260
rect 23584 28218 23612 28426
rect 23756 28416 23808 28422
rect 23756 28358 23808 28364
rect 23572 28212 23624 28218
rect 23572 28154 23624 28160
rect 23480 27872 23532 27878
rect 23480 27814 23532 27820
rect 23492 27606 23520 27814
rect 23480 27600 23532 27606
rect 23480 27542 23532 27548
rect 23584 27470 23612 28154
rect 23768 28150 23796 28358
rect 23756 28144 23808 28150
rect 23756 28086 23808 28092
rect 23664 27600 23716 27606
rect 23664 27542 23716 27548
rect 23572 27464 23624 27470
rect 23572 27406 23624 27412
rect 22928 27396 22980 27402
rect 22928 27338 22980 27344
rect 22940 25294 22968 27338
rect 23234 27228 23542 27237
rect 23234 27226 23240 27228
rect 23296 27226 23320 27228
rect 23376 27226 23400 27228
rect 23456 27226 23480 27228
rect 23536 27226 23542 27228
rect 23296 27174 23298 27226
rect 23478 27174 23480 27226
rect 23234 27172 23240 27174
rect 23296 27172 23320 27174
rect 23376 27172 23400 27174
rect 23456 27172 23480 27174
rect 23536 27172 23542 27174
rect 23234 27163 23542 27172
rect 23584 27062 23612 27406
rect 23676 27130 23704 27542
rect 23664 27124 23716 27130
rect 23664 27066 23716 27072
rect 23572 27056 23624 27062
rect 23572 26998 23624 27004
rect 24952 26988 25004 26994
rect 24952 26930 25004 26936
rect 23112 26920 23164 26926
rect 23112 26862 23164 26868
rect 24584 26920 24636 26926
rect 24584 26862 24636 26868
rect 23124 26518 23152 26862
rect 23112 26512 23164 26518
rect 23112 26454 23164 26460
rect 23124 26042 23152 26454
rect 23234 26140 23542 26149
rect 23234 26138 23240 26140
rect 23296 26138 23320 26140
rect 23376 26138 23400 26140
rect 23456 26138 23480 26140
rect 23536 26138 23542 26140
rect 23296 26086 23298 26138
rect 23478 26086 23480 26138
rect 23234 26084 23240 26086
rect 23296 26084 23320 26086
rect 23376 26084 23400 26086
rect 23456 26084 23480 26086
rect 23536 26084 23542 26086
rect 23234 26075 23542 26084
rect 23112 26036 23164 26042
rect 23112 25978 23164 25984
rect 24596 25838 24624 26862
rect 24964 26586 24992 26930
rect 24952 26580 25004 26586
rect 24952 26522 25004 26528
rect 25412 26444 25464 26450
rect 25412 26386 25464 26392
rect 24676 25900 24728 25906
rect 24676 25842 24728 25848
rect 24860 25900 24912 25906
rect 24860 25842 24912 25848
rect 24584 25832 24636 25838
rect 24584 25774 24636 25780
rect 22928 25288 22980 25294
rect 22928 25230 22980 25236
rect 22940 24206 22968 25230
rect 23664 25152 23716 25158
rect 23664 25094 23716 25100
rect 23234 25052 23542 25061
rect 23234 25050 23240 25052
rect 23296 25050 23320 25052
rect 23376 25050 23400 25052
rect 23456 25050 23480 25052
rect 23536 25050 23542 25052
rect 23296 24998 23298 25050
rect 23478 24998 23480 25050
rect 23234 24996 23240 24998
rect 23296 24996 23320 24998
rect 23376 24996 23400 24998
rect 23456 24996 23480 24998
rect 23536 24996 23542 24998
rect 23234 24987 23542 24996
rect 23112 24608 23164 24614
rect 23112 24550 23164 24556
rect 22928 24200 22980 24206
rect 22928 24142 22980 24148
rect 23124 23798 23152 24550
rect 23572 24064 23624 24070
rect 23572 24006 23624 24012
rect 23234 23964 23542 23973
rect 23234 23962 23240 23964
rect 23296 23962 23320 23964
rect 23376 23962 23400 23964
rect 23456 23962 23480 23964
rect 23536 23962 23542 23964
rect 23296 23910 23298 23962
rect 23478 23910 23480 23962
rect 23234 23908 23240 23910
rect 23296 23908 23320 23910
rect 23376 23908 23400 23910
rect 23456 23908 23480 23910
rect 23536 23908 23542 23910
rect 23234 23899 23542 23908
rect 23112 23792 23164 23798
rect 23112 23734 23164 23740
rect 23020 23520 23072 23526
rect 23020 23462 23072 23468
rect 23032 23118 23060 23462
rect 23124 23254 23152 23734
rect 23584 23254 23612 24006
rect 23112 23248 23164 23254
rect 23112 23190 23164 23196
rect 23572 23248 23624 23254
rect 23572 23190 23624 23196
rect 23676 23118 23704 25094
rect 24596 24750 24624 25774
rect 24584 24744 24636 24750
rect 24584 24686 24636 24692
rect 24596 23186 24624 24686
rect 24688 24138 24716 25842
rect 24872 25498 24900 25842
rect 24860 25492 24912 25498
rect 24860 25434 24912 25440
rect 25424 25362 25452 26386
rect 25504 26308 25556 26314
rect 25504 26250 25556 26256
rect 25412 25356 25464 25362
rect 25412 25298 25464 25304
rect 25044 25152 25096 25158
rect 25044 25094 25096 25100
rect 24952 24200 25004 24206
rect 24952 24142 25004 24148
rect 24676 24132 24728 24138
rect 24676 24074 24728 24080
rect 24584 23180 24636 23186
rect 24584 23122 24636 23128
rect 23020 23112 23072 23118
rect 23020 23054 23072 23060
rect 23112 23112 23164 23118
rect 23112 23054 23164 23060
rect 23664 23112 23716 23118
rect 23664 23054 23716 23060
rect 23124 22778 23152 23054
rect 23234 22876 23542 22885
rect 23234 22874 23240 22876
rect 23296 22874 23320 22876
rect 23376 22874 23400 22876
rect 23456 22874 23480 22876
rect 23536 22874 23542 22876
rect 23296 22822 23298 22874
rect 23478 22822 23480 22874
rect 23234 22820 23240 22822
rect 23296 22820 23320 22822
rect 23376 22820 23400 22822
rect 23456 22820 23480 22822
rect 23536 22820 23542 22822
rect 23234 22811 23542 22820
rect 23112 22772 23164 22778
rect 23112 22714 23164 22720
rect 23020 22704 23072 22710
rect 23020 22646 23072 22652
rect 22836 22024 22888 22030
rect 22836 21966 22888 21972
rect 23032 21690 23060 22646
rect 23112 22636 23164 22642
rect 23112 22578 23164 22584
rect 24584 22636 24636 22642
rect 24584 22578 24636 22584
rect 23020 21684 23072 21690
rect 23020 21626 23072 21632
rect 22652 21344 22704 21350
rect 22652 21286 22704 21292
rect 23124 20806 23152 22578
rect 23572 21956 23624 21962
rect 23572 21898 23624 21904
rect 23234 21788 23542 21797
rect 23234 21786 23240 21788
rect 23296 21786 23320 21788
rect 23376 21786 23400 21788
rect 23456 21786 23480 21788
rect 23536 21786 23542 21788
rect 23296 21734 23298 21786
rect 23478 21734 23480 21786
rect 23234 21732 23240 21734
rect 23296 21732 23320 21734
rect 23376 21732 23400 21734
rect 23456 21732 23480 21734
rect 23536 21732 23542 21734
rect 23234 21723 23542 21732
rect 23584 21554 23612 21898
rect 24596 21554 24624 22578
rect 24688 22114 24716 24074
rect 24860 24064 24912 24070
rect 24860 24006 24912 24012
rect 24872 23118 24900 24006
rect 24964 23322 24992 24142
rect 24952 23316 25004 23322
rect 24952 23258 25004 23264
rect 24860 23112 24912 23118
rect 24860 23054 24912 23060
rect 25056 22982 25084 25094
rect 25136 24268 25188 24274
rect 25136 24210 25188 24216
rect 25044 22976 25096 22982
rect 25044 22918 25096 22924
rect 24768 22636 24820 22642
rect 24768 22578 24820 22584
rect 24780 22234 24808 22578
rect 25148 22438 25176 24210
rect 25136 22432 25188 22438
rect 25136 22374 25188 22380
rect 24768 22228 24820 22234
rect 24768 22170 24820 22176
rect 24688 22086 24808 22114
rect 25148 22098 25176 22374
rect 23572 21548 23624 21554
rect 23572 21490 23624 21496
rect 24584 21548 24636 21554
rect 24584 21490 24636 21496
rect 24596 20942 24624 21490
rect 24676 21344 24728 21350
rect 24676 21286 24728 21292
rect 24688 20942 24716 21286
rect 24584 20936 24636 20942
rect 24584 20878 24636 20884
rect 24676 20936 24728 20942
rect 24676 20878 24728 20884
rect 23112 20800 23164 20806
rect 23112 20742 23164 20748
rect 23234 20700 23542 20709
rect 23234 20698 23240 20700
rect 23296 20698 23320 20700
rect 23376 20698 23400 20700
rect 23456 20698 23480 20700
rect 23536 20698 23542 20700
rect 23296 20646 23298 20698
rect 23478 20646 23480 20698
rect 23234 20644 23240 20646
rect 23296 20644 23320 20646
rect 23376 20644 23400 20646
rect 23456 20644 23480 20646
rect 23536 20644 23542 20646
rect 23234 20635 23542 20644
rect 23572 20528 23624 20534
rect 23572 20470 23624 20476
rect 23234 19612 23542 19621
rect 23234 19610 23240 19612
rect 23296 19610 23320 19612
rect 23376 19610 23400 19612
rect 23456 19610 23480 19612
rect 23536 19610 23542 19612
rect 23296 19558 23298 19610
rect 23478 19558 23480 19610
rect 23234 19556 23240 19558
rect 23296 19556 23320 19558
rect 23376 19556 23400 19558
rect 23456 19556 23480 19558
rect 23536 19556 23542 19558
rect 23234 19547 23542 19556
rect 23584 19378 23612 20470
rect 24596 20466 24624 20878
rect 24584 20460 24636 20466
rect 24584 20402 24636 20408
rect 23572 19372 23624 19378
rect 23572 19314 23624 19320
rect 23664 19372 23716 19378
rect 23664 19314 23716 19320
rect 23676 18834 23704 19314
rect 24596 18834 24624 20402
rect 24676 19712 24728 19718
rect 24676 19654 24728 19660
rect 24688 19446 24716 19654
rect 24676 19440 24728 19446
rect 24676 19382 24728 19388
rect 22928 18828 22980 18834
rect 22928 18770 22980 18776
rect 23664 18828 23716 18834
rect 23664 18770 23716 18776
rect 24584 18828 24636 18834
rect 24584 18770 24636 18776
rect 22468 18624 22520 18630
rect 22468 18566 22520 18572
rect 22192 18420 22244 18426
rect 22192 18362 22244 18368
rect 22940 18222 22968 18770
rect 23234 18524 23542 18533
rect 23234 18522 23240 18524
rect 23296 18522 23320 18524
rect 23376 18522 23400 18524
rect 23456 18522 23480 18524
rect 23536 18522 23542 18524
rect 23296 18470 23298 18522
rect 23478 18470 23480 18522
rect 23234 18468 23240 18470
rect 23296 18468 23320 18470
rect 23376 18468 23400 18470
rect 23456 18468 23480 18470
rect 23536 18468 23542 18470
rect 23234 18459 23542 18468
rect 21456 18216 21508 18222
rect 21456 18158 21508 18164
rect 22928 18216 22980 18222
rect 22928 18158 22980 18164
rect 21468 17882 21496 18158
rect 22008 18080 22060 18086
rect 22008 18022 22060 18028
rect 21456 17876 21508 17882
rect 21456 17818 21508 17824
rect 21272 16992 21324 16998
rect 21272 16934 21324 16940
rect 20916 16546 21220 16574
rect 19984 15632 20036 15638
rect 19984 15574 20036 15580
rect 19892 14952 19944 14958
rect 19892 14894 19944 14900
rect 19520 14716 19828 14725
rect 19520 14714 19526 14716
rect 19582 14714 19606 14716
rect 19662 14714 19686 14716
rect 19742 14714 19766 14716
rect 19822 14714 19828 14716
rect 19582 14662 19584 14714
rect 19764 14662 19766 14714
rect 19520 14660 19526 14662
rect 19582 14660 19606 14662
rect 19662 14660 19686 14662
rect 19742 14660 19766 14662
rect 19822 14660 19828 14662
rect 19520 14651 19828 14660
rect 19996 14498 20024 15574
rect 20720 15360 20772 15366
rect 20720 15302 20772 15308
rect 20732 15094 20760 15302
rect 20720 15088 20772 15094
rect 20720 15030 20772 15036
rect 20916 14618 20944 16546
rect 21088 15360 21140 15366
rect 21088 15302 21140 15308
rect 21180 15360 21232 15366
rect 21180 15302 21232 15308
rect 21100 15094 21128 15302
rect 21088 15088 21140 15094
rect 21088 15030 21140 15036
rect 21192 15026 21220 15302
rect 21180 15020 21232 15026
rect 21180 14962 21232 14968
rect 20996 14884 21048 14890
rect 20996 14826 21048 14832
rect 20904 14612 20956 14618
rect 20904 14554 20956 14560
rect 21008 14550 21036 14826
rect 21284 14618 21312 16934
rect 21468 15502 21496 17818
rect 22020 17678 22048 18022
rect 22008 17672 22060 17678
rect 22008 17614 22060 17620
rect 22744 17672 22796 17678
rect 22744 17614 22796 17620
rect 22468 17604 22520 17610
rect 22468 17546 22520 17552
rect 22480 17338 22508 17546
rect 22468 17332 22520 17338
rect 22468 17274 22520 17280
rect 22756 17202 22784 17614
rect 22744 17196 22796 17202
rect 22744 17138 22796 17144
rect 22008 16584 22060 16590
rect 22008 16526 22060 16532
rect 21456 15496 21508 15502
rect 21456 15438 21508 15444
rect 22020 15162 22048 16526
rect 22756 15502 22784 17138
rect 22940 17134 22968 18158
rect 23676 17610 23704 18770
rect 23664 17604 23716 17610
rect 23664 17546 23716 17552
rect 23572 17536 23624 17542
rect 23572 17478 23624 17484
rect 23234 17436 23542 17445
rect 23234 17434 23240 17436
rect 23296 17434 23320 17436
rect 23376 17434 23400 17436
rect 23456 17434 23480 17436
rect 23536 17434 23542 17436
rect 23296 17382 23298 17434
rect 23478 17382 23480 17434
rect 23234 17380 23240 17382
rect 23296 17380 23320 17382
rect 23376 17380 23400 17382
rect 23456 17380 23480 17382
rect 23536 17380 23542 17382
rect 23234 17371 23542 17380
rect 23584 17202 23612 17478
rect 23572 17196 23624 17202
rect 23572 17138 23624 17144
rect 22928 17128 22980 17134
rect 22928 17070 22980 17076
rect 23112 16516 23164 16522
rect 23112 16458 23164 16464
rect 22744 15496 22796 15502
rect 22744 15438 22796 15444
rect 22008 15156 22060 15162
rect 22008 15098 22060 15104
rect 21916 15020 21968 15026
rect 21916 14962 21968 14968
rect 21928 14618 21956 14962
rect 21272 14612 21324 14618
rect 21272 14554 21324 14560
rect 21916 14612 21968 14618
rect 21916 14554 21968 14560
rect 20996 14544 21048 14550
rect 19996 14470 20116 14498
rect 20996 14486 21048 14492
rect 19984 14340 20036 14346
rect 19984 14282 20036 14288
rect 19996 14074 20024 14282
rect 19984 14068 20036 14074
rect 19984 14010 20036 14016
rect 20088 13802 20116 14470
rect 20904 14476 20956 14482
rect 20904 14418 20956 14424
rect 20916 14278 20944 14418
rect 21732 14408 21784 14414
rect 21732 14350 21784 14356
rect 21456 14340 21508 14346
rect 21456 14282 21508 14288
rect 21548 14340 21600 14346
rect 21548 14282 21600 14288
rect 20904 14272 20956 14278
rect 20904 14214 20956 14220
rect 20996 14272 21048 14278
rect 20996 14214 21048 14220
rect 21008 14074 21036 14214
rect 20996 14068 21048 14074
rect 20996 14010 21048 14016
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 20076 13796 20128 13802
rect 20076 13738 20128 13744
rect 19520 13628 19828 13637
rect 19520 13626 19526 13628
rect 19582 13626 19606 13628
rect 19662 13626 19686 13628
rect 19742 13626 19766 13628
rect 19822 13626 19828 13628
rect 19582 13574 19584 13626
rect 19764 13574 19766 13626
rect 19520 13572 19526 13574
rect 19582 13572 19606 13574
rect 19662 13572 19686 13574
rect 19742 13572 19766 13574
rect 19822 13572 19828 13574
rect 19520 13563 19828 13572
rect 20456 13530 20484 13874
rect 20444 13524 20496 13530
rect 20444 13466 20496 13472
rect 21008 13394 21036 14010
rect 20996 13388 21048 13394
rect 20996 13330 21048 13336
rect 19892 12844 19944 12850
rect 19892 12786 19944 12792
rect 19432 12708 19484 12714
rect 19432 12650 19484 12656
rect 19520 12540 19828 12549
rect 19520 12538 19526 12540
rect 19582 12538 19606 12540
rect 19662 12538 19686 12540
rect 19742 12538 19766 12540
rect 19822 12538 19828 12540
rect 19582 12486 19584 12538
rect 19764 12486 19766 12538
rect 19520 12484 19526 12486
rect 19582 12484 19606 12486
rect 19662 12484 19686 12486
rect 19742 12484 19766 12486
rect 19822 12484 19828 12486
rect 19520 12475 19828 12484
rect 19904 11762 19932 12786
rect 21468 12782 21496 14282
rect 21560 13530 21588 14282
rect 21744 13938 21772 14350
rect 21732 13932 21784 13938
rect 21732 13874 21784 13880
rect 21548 13524 21600 13530
rect 21548 13466 21600 13472
rect 21456 12776 21508 12782
rect 21456 12718 21508 12724
rect 19892 11756 19944 11762
rect 19892 11698 19944 11704
rect 20444 11756 20496 11762
rect 20444 11698 20496 11704
rect 19432 11552 19484 11558
rect 19432 11494 19484 11500
rect 19892 11552 19944 11558
rect 19892 11494 19944 11500
rect 19444 11218 19472 11494
rect 19520 11452 19828 11461
rect 19520 11450 19526 11452
rect 19582 11450 19606 11452
rect 19662 11450 19686 11452
rect 19742 11450 19766 11452
rect 19822 11450 19828 11452
rect 19582 11398 19584 11450
rect 19764 11398 19766 11450
rect 19520 11396 19526 11398
rect 19582 11396 19606 11398
rect 19662 11396 19686 11398
rect 19742 11396 19766 11398
rect 19822 11396 19828 11398
rect 19520 11387 19828 11396
rect 19904 11234 19932 11494
rect 20456 11354 20484 11698
rect 22020 11642 22048 15098
rect 22468 14952 22520 14958
rect 22468 14894 22520 14900
rect 22480 14074 22508 14894
rect 22756 14822 22784 15438
rect 22744 14816 22796 14822
rect 22744 14758 22796 14764
rect 22468 14068 22520 14074
rect 22468 14010 22520 14016
rect 23124 14006 23152 16458
rect 23234 16348 23542 16357
rect 23234 16346 23240 16348
rect 23296 16346 23320 16348
rect 23376 16346 23400 16348
rect 23456 16346 23480 16348
rect 23536 16346 23542 16348
rect 23296 16294 23298 16346
rect 23478 16294 23480 16346
rect 23234 16292 23240 16294
rect 23296 16292 23320 16294
rect 23376 16292 23400 16294
rect 23456 16292 23480 16294
rect 23536 16292 23542 16294
rect 23234 16283 23542 16292
rect 24780 16114 24808 22086
rect 25136 22092 25188 22098
rect 25136 22034 25188 22040
rect 25148 21486 25176 22034
rect 25228 21684 25280 21690
rect 25228 21626 25280 21632
rect 25136 21480 25188 21486
rect 25136 21422 25188 21428
rect 25240 21434 25268 21626
rect 25516 21554 25544 26250
rect 25700 23730 25728 28970
rect 26948 28860 27256 28869
rect 26948 28858 26954 28860
rect 27010 28858 27034 28860
rect 27090 28858 27114 28860
rect 27170 28858 27194 28860
rect 27250 28858 27256 28860
rect 27010 28806 27012 28858
rect 27192 28806 27194 28858
rect 26948 28804 26954 28806
rect 27010 28804 27034 28806
rect 27090 28804 27114 28806
rect 27170 28804 27194 28806
rect 27250 28804 27256 28806
rect 26948 28795 27256 28804
rect 26424 28552 26476 28558
rect 26424 28494 26476 28500
rect 27896 28552 27948 28558
rect 27896 28494 27948 28500
rect 25872 27532 25924 27538
rect 25872 27474 25924 27480
rect 26056 27532 26108 27538
rect 26056 27474 26108 27480
rect 25884 26858 25912 27474
rect 25872 26852 25924 26858
rect 25872 26794 25924 26800
rect 25884 26518 25912 26794
rect 25964 26784 26016 26790
rect 25964 26726 26016 26732
rect 25872 26512 25924 26518
rect 25872 26454 25924 26460
rect 25976 26450 26004 26726
rect 26068 26586 26096 27474
rect 26436 27470 26464 28494
rect 27620 28484 27672 28490
rect 27620 28426 27672 28432
rect 27436 28416 27488 28422
rect 27436 28358 27488 28364
rect 27448 28150 27476 28358
rect 27436 28144 27488 28150
rect 27436 28086 27488 28092
rect 26608 28008 26660 28014
rect 26608 27950 26660 27956
rect 26620 27674 26648 27950
rect 26948 27772 27256 27781
rect 26948 27770 26954 27772
rect 27010 27770 27034 27772
rect 27090 27770 27114 27772
rect 27170 27770 27194 27772
rect 27250 27770 27256 27772
rect 27010 27718 27012 27770
rect 27192 27718 27194 27770
rect 26948 27716 26954 27718
rect 27010 27716 27034 27718
rect 27090 27716 27114 27718
rect 27170 27716 27194 27718
rect 27250 27716 27256 27718
rect 26948 27707 27256 27716
rect 26608 27668 26660 27674
rect 26608 27610 26660 27616
rect 27632 27470 27660 28426
rect 27908 27470 27936 28494
rect 28172 28144 28224 28150
rect 28172 28086 28224 28092
rect 28184 27538 28212 28086
rect 28172 27532 28224 27538
rect 28172 27474 28224 27480
rect 26424 27464 26476 27470
rect 26424 27406 26476 27412
rect 26608 27464 26660 27470
rect 26608 27406 26660 27412
rect 27620 27464 27672 27470
rect 27620 27406 27672 27412
rect 27896 27464 27948 27470
rect 27896 27406 27948 27412
rect 26148 27396 26200 27402
rect 26148 27338 26200 27344
rect 26160 26790 26188 27338
rect 26148 26784 26200 26790
rect 26148 26726 26200 26732
rect 26056 26580 26108 26586
rect 26056 26522 26108 26528
rect 26148 26580 26200 26586
rect 26148 26522 26200 26528
rect 25964 26444 26016 26450
rect 25964 26386 26016 26392
rect 26056 26308 26108 26314
rect 26056 26250 26108 26256
rect 25964 25696 26016 25702
rect 25964 25638 26016 25644
rect 25976 25362 26004 25638
rect 25964 25356 26016 25362
rect 25964 25298 26016 25304
rect 26068 24750 26096 26250
rect 25780 24744 25832 24750
rect 25780 24686 25832 24692
rect 26056 24744 26108 24750
rect 26056 24686 26108 24692
rect 25792 24070 25820 24686
rect 26160 24274 26188 26522
rect 26332 26376 26384 26382
rect 26332 26318 26384 26324
rect 26344 25430 26372 26318
rect 26620 26314 26648 27406
rect 27632 27334 27660 27406
rect 27620 27328 27672 27334
rect 27620 27270 27672 27276
rect 26948 26684 27256 26693
rect 26948 26682 26954 26684
rect 27010 26682 27034 26684
rect 27090 26682 27114 26684
rect 27170 26682 27194 26684
rect 27250 26682 27256 26684
rect 27010 26630 27012 26682
rect 27192 26630 27194 26682
rect 26948 26628 26954 26630
rect 27010 26628 27034 26630
rect 27090 26628 27114 26630
rect 27170 26628 27194 26630
rect 27250 26628 27256 26630
rect 26948 26619 27256 26628
rect 27632 26450 27660 27270
rect 27620 26444 27672 26450
rect 27620 26386 27672 26392
rect 26608 26308 26660 26314
rect 26608 26250 26660 26256
rect 26332 25424 26384 25430
rect 26332 25366 26384 25372
rect 26424 25356 26476 25362
rect 26424 25298 26476 25304
rect 26148 24268 26200 24274
rect 26148 24210 26200 24216
rect 26332 24200 26384 24206
rect 26332 24142 26384 24148
rect 25780 24064 25832 24070
rect 25780 24006 25832 24012
rect 26148 24064 26200 24070
rect 26148 24006 26200 24012
rect 25688 23724 25740 23730
rect 25688 23666 25740 23672
rect 25700 21962 25728 23666
rect 25792 23322 25820 24006
rect 25964 23724 26016 23730
rect 25964 23666 26016 23672
rect 25780 23316 25832 23322
rect 25780 23258 25832 23264
rect 25872 23180 25924 23186
rect 25872 23122 25924 23128
rect 25884 22778 25912 23122
rect 25872 22772 25924 22778
rect 25872 22714 25924 22720
rect 25884 22030 25912 22714
rect 25976 22098 26004 23666
rect 25964 22092 26016 22098
rect 25964 22034 26016 22040
rect 25872 22024 25924 22030
rect 25872 21966 25924 21972
rect 25688 21956 25740 21962
rect 25688 21898 25740 21904
rect 25504 21548 25556 21554
rect 25504 21490 25556 21496
rect 25320 21480 25372 21486
rect 25240 21428 25320 21434
rect 25240 21422 25372 21428
rect 24860 21412 24912 21418
rect 24860 21354 24912 21360
rect 25240 21406 25360 21422
rect 26160 21418 26188 24006
rect 26344 23866 26372 24142
rect 26332 23860 26384 23866
rect 26332 23802 26384 23808
rect 26436 23662 26464 25298
rect 26620 25294 26648 26250
rect 26948 25596 27256 25605
rect 26948 25594 26954 25596
rect 27010 25594 27034 25596
rect 27090 25594 27114 25596
rect 27170 25594 27194 25596
rect 27250 25594 27256 25596
rect 27010 25542 27012 25594
rect 27192 25542 27194 25594
rect 26948 25540 26954 25542
rect 27010 25540 27034 25542
rect 27090 25540 27114 25542
rect 27170 25540 27194 25542
rect 27250 25540 27256 25542
rect 26948 25531 27256 25540
rect 26608 25288 26660 25294
rect 26608 25230 26660 25236
rect 26948 24508 27256 24517
rect 26948 24506 26954 24508
rect 27010 24506 27034 24508
rect 27090 24506 27114 24508
rect 27170 24506 27194 24508
rect 27250 24506 27256 24508
rect 27010 24454 27012 24506
rect 27192 24454 27194 24506
rect 26948 24452 26954 24454
rect 27010 24452 27034 24454
rect 27090 24452 27114 24454
rect 27170 24452 27194 24454
rect 27250 24452 27256 24454
rect 26948 24443 27256 24452
rect 27632 24274 27660 26386
rect 27908 26382 27936 27406
rect 27896 26376 27948 26382
rect 27896 26318 27948 26324
rect 27804 25288 27856 25294
rect 27804 25230 27856 25236
rect 27816 24818 27844 25230
rect 27804 24812 27856 24818
rect 27804 24754 27856 24760
rect 27620 24268 27672 24274
rect 27620 24210 27672 24216
rect 27908 24206 27936 26318
rect 27988 25832 28040 25838
rect 27988 25774 28040 25780
rect 28000 25498 28028 25774
rect 27988 25492 28040 25498
rect 27988 25434 28040 25440
rect 28448 25152 28500 25158
rect 28448 25094 28500 25100
rect 28460 24886 28488 25094
rect 28448 24880 28500 24886
rect 28448 24822 28500 24828
rect 28264 24608 28316 24614
rect 28264 24550 28316 24556
rect 27896 24200 27948 24206
rect 27896 24142 27948 24148
rect 28172 24200 28224 24206
rect 28172 24142 28224 24148
rect 28184 23798 28212 24142
rect 28276 23866 28304 24550
rect 28448 24200 28500 24206
rect 28448 24142 28500 24148
rect 28264 23860 28316 23866
rect 28264 23802 28316 23808
rect 28172 23792 28224 23798
rect 28172 23734 28224 23740
rect 26516 23724 26568 23730
rect 26516 23666 26568 23672
rect 26424 23656 26476 23662
rect 26424 23598 26476 23604
rect 26528 23322 26556 23666
rect 26948 23420 27256 23429
rect 26948 23418 26954 23420
rect 27010 23418 27034 23420
rect 27090 23418 27114 23420
rect 27170 23418 27194 23420
rect 27250 23418 27256 23420
rect 27010 23366 27012 23418
rect 27192 23366 27194 23418
rect 26948 23364 26954 23366
rect 27010 23364 27034 23366
rect 27090 23364 27114 23366
rect 27170 23364 27194 23366
rect 27250 23364 27256 23366
rect 26948 23355 27256 23364
rect 26516 23316 26568 23322
rect 26516 23258 26568 23264
rect 26948 22332 27256 22341
rect 26948 22330 26954 22332
rect 27010 22330 27034 22332
rect 27090 22330 27114 22332
rect 27170 22330 27194 22332
rect 27250 22330 27256 22332
rect 27010 22278 27012 22330
rect 27192 22278 27194 22330
rect 26948 22276 26954 22278
rect 27010 22276 27034 22278
rect 27090 22276 27114 22278
rect 27170 22276 27194 22278
rect 27250 22276 27256 22278
rect 26948 22267 27256 22276
rect 26240 22092 26292 22098
rect 26240 22034 26292 22040
rect 26252 21622 26280 22034
rect 28184 22030 28212 23734
rect 28356 22976 28408 22982
rect 28356 22918 28408 22924
rect 28368 22642 28396 22918
rect 28356 22636 28408 22642
rect 28356 22578 28408 22584
rect 28460 22030 28488 24142
rect 28552 24138 28580 29038
rect 28908 27872 28960 27878
rect 28908 27814 28960 27820
rect 28920 27470 28948 27814
rect 29012 27606 29040 29038
rect 29184 28416 29236 28422
rect 29184 28358 29236 28364
rect 29000 27600 29052 27606
rect 29000 27542 29052 27548
rect 28908 27464 28960 27470
rect 28908 27406 28960 27412
rect 29196 27062 29224 28358
rect 30662 28316 30970 28325
rect 30662 28314 30668 28316
rect 30724 28314 30748 28316
rect 30804 28314 30828 28316
rect 30884 28314 30908 28316
rect 30964 28314 30970 28316
rect 30724 28262 30726 28314
rect 30906 28262 30908 28314
rect 30662 28260 30668 28262
rect 30724 28260 30748 28262
rect 30804 28260 30828 28262
rect 30884 28260 30908 28262
rect 30964 28260 30970 28262
rect 30662 28251 30970 28260
rect 29460 28076 29512 28082
rect 29460 28018 29512 28024
rect 29184 27056 29236 27062
rect 29184 26998 29236 27004
rect 29472 26790 29500 28018
rect 29920 27872 29972 27878
rect 29920 27814 29972 27820
rect 29932 27062 29960 27814
rect 30196 27328 30248 27334
rect 30196 27270 30248 27276
rect 29920 27056 29972 27062
rect 29920 26998 29972 27004
rect 30208 26994 30236 27270
rect 30662 27228 30970 27237
rect 30662 27226 30668 27228
rect 30724 27226 30748 27228
rect 30804 27226 30828 27228
rect 30884 27226 30908 27228
rect 30964 27226 30970 27228
rect 30724 27174 30726 27226
rect 30906 27174 30908 27226
rect 30662 27172 30668 27174
rect 30724 27172 30748 27174
rect 30804 27172 30828 27174
rect 30884 27172 30908 27174
rect 30964 27172 30970 27174
rect 30662 27163 30970 27172
rect 30196 26988 30248 26994
rect 30196 26930 30248 26936
rect 29460 26784 29512 26790
rect 29460 26726 29512 26732
rect 29920 26376 29972 26382
rect 29920 26318 29972 26324
rect 29184 26240 29236 26246
rect 29184 26182 29236 26188
rect 29828 26240 29880 26246
rect 29828 26182 29880 26188
rect 29196 25974 29224 26182
rect 29184 25968 29236 25974
rect 29184 25910 29236 25916
rect 29840 25838 29868 26182
rect 29932 26042 29960 26318
rect 30662 26140 30970 26149
rect 30662 26138 30668 26140
rect 30724 26138 30748 26140
rect 30804 26138 30828 26140
rect 30884 26138 30908 26140
rect 30964 26138 30970 26140
rect 30724 26086 30726 26138
rect 30906 26086 30908 26138
rect 30662 26084 30668 26086
rect 30724 26084 30748 26086
rect 30804 26084 30828 26086
rect 30884 26084 30908 26086
rect 30964 26084 30970 26086
rect 30662 26075 30970 26084
rect 29920 26036 29972 26042
rect 29920 25978 29972 25984
rect 29828 25832 29880 25838
rect 29828 25774 29880 25780
rect 31022 25800 31078 25809
rect 31022 25735 31078 25744
rect 31036 25362 31064 25735
rect 31024 25356 31076 25362
rect 31024 25298 31076 25304
rect 28908 25288 28960 25294
rect 28908 25230 28960 25236
rect 29828 25288 29880 25294
rect 29828 25230 29880 25236
rect 28920 24750 28948 25230
rect 29552 24812 29604 24818
rect 29552 24754 29604 24760
rect 28908 24744 28960 24750
rect 28908 24686 28960 24692
rect 29564 24274 29592 24754
rect 29552 24268 29604 24274
rect 29552 24210 29604 24216
rect 28540 24132 28592 24138
rect 28540 24074 28592 24080
rect 28908 23724 28960 23730
rect 28908 23666 28960 23672
rect 28920 23118 28948 23666
rect 28540 23112 28592 23118
rect 28540 23054 28592 23060
rect 28908 23112 28960 23118
rect 28908 23054 28960 23060
rect 27620 22024 27672 22030
rect 27620 21966 27672 21972
rect 28172 22024 28224 22030
rect 28172 21966 28224 21972
rect 28448 22024 28500 22030
rect 28448 21966 28500 21972
rect 27632 21690 27660 21966
rect 27896 21888 27948 21894
rect 27896 21830 27948 21836
rect 27620 21684 27672 21690
rect 27620 21626 27672 21632
rect 27908 21622 27936 21830
rect 26240 21616 26292 21622
rect 26240 21558 26292 21564
rect 27896 21616 27948 21622
rect 27896 21558 27948 21564
rect 26148 21412 26200 21418
rect 24872 21146 24900 21354
rect 24860 21140 24912 21146
rect 24860 21082 24912 21088
rect 24860 18692 24912 18698
rect 24860 18634 24912 18640
rect 24872 18426 24900 18634
rect 24860 18420 24912 18426
rect 24860 18362 24912 18368
rect 25240 18290 25268 21406
rect 26148 21354 26200 21360
rect 26252 21146 26280 21558
rect 27620 21480 27672 21486
rect 27620 21422 27672 21428
rect 26700 21412 26752 21418
rect 26700 21354 26752 21360
rect 26240 21140 26292 21146
rect 26240 21082 26292 21088
rect 25320 20256 25372 20262
rect 25320 20198 25372 20204
rect 25332 18698 25360 20198
rect 26712 19922 26740 21354
rect 26948 21244 27256 21253
rect 26948 21242 26954 21244
rect 27010 21242 27034 21244
rect 27090 21242 27114 21244
rect 27170 21242 27194 21244
rect 27250 21242 27256 21244
rect 27010 21190 27012 21242
rect 27192 21190 27194 21242
rect 26948 21188 26954 21190
rect 27010 21188 27034 21190
rect 27090 21188 27114 21190
rect 27170 21188 27194 21190
rect 27250 21188 27256 21190
rect 26948 21179 27256 21188
rect 27632 21146 27660 21422
rect 27620 21140 27672 21146
rect 27620 21082 27672 21088
rect 28184 21010 28212 21966
rect 28172 21004 28224 21010
rect 28172 20946 28224 20952
rect 28460 20942 28488 21966
rect 28552 21690 28580 23054
rect 28632 22976 28684 22982
rect 28632 22918 28684 22924
rect 28644 22710 28672 22918
rect 28920 22778 28948 23054
rect 28908 22772 28960 22778
rect 28908 22714 28960 22720
rect 28632 22704 28684 22710
rect 28632 22646 28684 22652
rect 29184 22704 29236 22710
rect 29184 22646 29236 22652
rect 29196 22098 29224 22646
rect 29184 22092 29236 22098
rect 29184 22034 29236 22040
rect 29368 22024 29420 22030
rect 29368 21966 29420 21972
rect 28540 21684 28592 21690
rect 28540 21626 28592 21632
rect 29000 21548 29052 21554
rect 29000 21490 29052 21496
rect 29012 21010 29040 21490
rect 29000 21004 29052 21010
rect 29000 20946 29052 20952
rect 28448 20936 28500 20942
rect 28448 20878 28500 20884
rect 26948 20156 27256 20165
rect 26948 20154 26954 20156
rect 27010 20154 27034 20156
rect 27090 20154 27114 20156
rect 27170 20154 27194 20156
rect 27250 20154 27256 20156
rect 27010 20102 27012 20154
rect 27192 20102 27194 20154
rect 26948 20100 26954 20102
rect 27010 20100 27034 20102
rect 27090 20100 27114 20102
rect 27170 20100 27194 20102
rect 27250 20100 27256 20102
rect 26948 20091 27256 20100
rect 27988 20052 28040 20058
rect 27988 19994 28040 20000
rect 25412 19916 25464 19922
rect 25412 19858 25464 19864
rect 26700 19916 26752 19922
rect 26700 19858 26752 19864
rect 25424 18970 25452 19858
rect 25872 19712 25924 19718
rect 25872 19654 25924 19660
rect 25884 19514 25912 19654
rect 25872 19508 25924 19514
rect 25872 19450 25924 19456
rect 27436 19508 27488 19514
rect 27436 19450 27488 19456
rect 26948 19068 27256 19077
rect 26948 19066 26954 19068
rect 27010 19066 27034 19068
rect 27090 19066 27114 19068
rect 27170 19066 27194 19068
rect 27250 19066 27256 19068
rect 27010 19014 27012 19066
rect 27192 19014 27194 19066
rect 26948 19012 26954 19014
rect 27010 19012 27034 19014
rect 27090 19012 27114 19014
rect 27170 19012 27194 19014
rect 27250 19012 27256 19014
rect 26948 19003 27256 19012
rect 25412 18964 25464 18970
rect 25412 18906 25464 18912
rect 25320 18692 25372 18698
rect 25320 18634 25372 18640
rect 25228 18284 25280 18290
rect 25228 18226 25280 18232
rect 25240 17678 25268 18226
rect 25424 18222 25452 18906
rect 27448 18766 27476 19450
rect 28000 19446 28028 19994
rect 28448 19780 28500 19786
rect 28448 19722 28500 19728
rect 27988 19440 28040 19446
rect 27988 19382 28040 19388
rect 27712 19236 27764 19242
rect 27712 19178 27764 19184
rect 27436 18760 27488 18766
rect 27436 18702 27488 18708
rect 27724 18698 27752 19178
rect 28000 18902 28028 19382
rect 28460 18970 28488 19722
rect 28632 19712 28684 19718
rect 28632 19654 28684 19660
rect 28644 19514 28672 19654
rect 28632 19508 28684 19514
rect 28632 19450 28684 19456
rect 28448 18964 28500 18970
rect 28448 18906 28500 18912
rect 27988 18896 28040 18902
rect 27988 18838 28040 18844
rect 28644 18766 28672 19450
rect 29000 19372 29052 19378
rect 29000 19314 29052 19320
rect 29184 19372 29236 19378
rect 29184 19314 29236 19320
rect 29012 18970 29040 19314
rect 29196 19174 29224 19314
rect 29380 19310 29408 21966
rect 29840 21078 29868 25230
rect 30662 25052 30970 25061
rect 30662 25050 30668 25052
rect 30724 25050 30748 25052
rect 30804 25050 30828 25052
rect 30884 25050 30908 25052
rect 30964 25050 30970 25052
rect 30724 24998 30726 25050
rect 30906 24998 30908 25050
rect 30662 24996 30668 24998
rect 30724 24996 30748 24998
rect 30804 24996 30828 24998
rect 30884 24996 30908 24998
rect 30964 24996 30970 24998
rect 30662 24987 30970 24996
rect 30662 23964 30970 23973
rect 30662 23962 30668 23964
rect 30724 23962 30748 23964
rect 30804 23962 30828 23964
rect 30884 23962 30908 23964
rect 30964 23962 30970 23964
rect 30724 23910 30726 23962
rect 30906 23910 30908 23962
rect 30662 23908 30668 23910
rect 30724 23908 30748 23910
rect 30804 23908 30828 23910
rect 30884 23908 30908 23910
rect 30964 23908 30970 23910
rect 30662 23899 30970 23908
rect 30662 22876 30970 22885
rect 30662 22874 30668 22876
rect 30724 22874 30748 22876
rect 30804 22874 30828 22876
rect 30884 22874 30908 22876
rect 30964 22874 30970 22876
rect 30724 22822 30726 22874
rect 30906 22822 30908 22874
rect 30662 22820 30668 22822
rect 30724 22820 30748 22822
rect 30804 22820 30828 22822
rect 30884 22820 30908 22822
rect 30964 22820 30970 22822
rect 30662 22811 30970 22820
rect 31022 21992 31078 22001
rect 31022 21927 31024 21936
rect 31076 21927 31078 21936
rect 31024 21898 31076 21904
rect 30662 21788 30970 21797
rect 30662 21786 30668 21788
rect 30724 21786 30748 21788
rect 30804 21786 30828 21788
rect 30884 21786 30908 21788
rect 30964 21786 30970 21788
rect 30724 21734 30726 21786
rect 30906 21734 30908 21786
rect 30662 21732 30668 21734
rect 30724 21732 30748 21734
rect 30804 21732 30828 21734
rect 30884 21732 30908 21734
rect 30964 21732 30970 21734
rect 30662 21723 30970 21732
rect 29828 21072 29880 21078
rect 29828 21014 29880 21020
rect 30662 20700 30970 20709
rect 30662 20698 30668 20700
rect 30724 20698 30748 20700
rect 30804 20698 30828 20700
rect 30884 20698 30908 20700
rect 30964 20698 30970 20700
rect 30724 20646 30726 20698
rect 30906 20646 30908 20698
rect 30662 20644 30668 20646
rect 30724 20644 30748 20646
rect 30804 20644 30828 20646
rect 30884 20644 30908 20646
rect 30964 20644 30970 20646
rect 30662 20635 30970 20644
rect 30662 19612 30970 19621
rect 30662 19610 30668 19612
rect 30724 19610 30748 19612
rect 30804 19610 30828 19612
rect 30884 19610 30908 19612
rect 30964 19610 30970 19612
rect 30724 19558 30726 19610
rect 30906 19558 30908 19610
rect 30662 19556 30668 19558
rect 30724 19556 30748 19558
rect 30804 19556 30828 19558
rect 30884 19556 30908 19558
rect 30964 19556 30970 19558
rect 30662 19547 30970 19556
rect 29920 19440 29972 19446
rect 29920 19382 29972 19388
rect 29368 19304 29420 19310
rect 29368 19246 29420 19252
rect 29184 19168 29236 19174
rect 29184 19110 29236 19116
rect 29000 18964 29052 18970
rect 29000 18906 29052 18912
rect 29196 18766 29224 19110
rect 29932 18834 29960 19382
rect 29828 18828 29880 18834
rect 29828 18770 29880 18776
rect 29920 18828 29972 18834
rect 29920 18770 29972 18776
rect 28632 18760 28684 18766
rect 28632 18702 28684 18708
rect 29184 18760 29236 18766
rect 29184 18702 29236 18708
rect 27712 18692 27764 18698
rect 27712 18634 27764 18640
rect 26332 18624 26384 18630
rect 26332 18566 26384 18572
rect 26344 18426 26372 18566
rect 26332 18420 26384 18426
rect 26332 18362 26384 18368
rect 29840 18290 29868 18770
rect 29828 18284 29880 18290
rect 29828 18226 29880 18232
rect 25412 18216 25464 18222
rect 25412 18158 25464 18164
rect 25228 17672 25280 17678
rect 25228 17614 25280 17620
rect 24952 16992 25004 16998
rect 24952 16934 25004 16940
rect 23756 16108 23808 16114
rect 23756 16050 23808 16056
rect 24400 16108 24452 16114
rect 24400 16050 24452 16056
rect 24768 16108 24820 16114
rect 24768 16050 24820 16056
rect 23664 16040 23716 16046
rect 23664 15982 23716 15988
rect 23572 15360 23624 15366
rect 23572 15302 23624 15308
rect 23234 15260 23542 15269
rect 23234 15258 23240 15260
rect 23296 15258 23320 15260
rect 23376 15258 23400 15260
rect 23456 15258 23480 15260
rect 23536 15258 23542 15260
rect 23296 15206 23298 15258
rect 23478 15206 23480 15258
rect 23234 15204 23240 15206
rect 23296 15204 23320 15206
rect 23376 15204 23400 15206
rect 23456 15204 23480 15206
rect 23536 15204 23542 15206
rect 23234 15195 23542 15204
rect 23584 15094 23612 15302
rect 23676 15094 23704 15982
rect 23768 15502 23796 16050
rect 24308 16040 24360 16046
rect 24308 15982 24360 15988
rect 24320 15638 24348 15982
rect 24308 15632 24360 15638
rect 24308 15574 24360 15580
rect 23756 15496 23808 15502
rect 23756 15438 23808 15444
rect 23572 15088 23624 15094
rect 23572 15030 23624 15036
rect 23664 15088 23716 15094
rect 23664 15030 23716 15036
rect 23234 14172 23542 14181
rect 23234 14170 23240 14172
rect 23296 14170 23320 14172
rect 23376 14170 23400 14172
rect 23456 14170 23480 14172
rect 23536 14170 23542 14172
rect 23296 14118 23298 14170
rect 23478 14118 23480 14170
rect 23234 14116 23240 14118
rect 23296 14116 23320 14118
rect 23376 14116 23400 14118
rect 23456 14116 23480 14118
rect 23536 14116 23542 14118
rect 23234 14107 23542 14116
rect 23112 14000 23164 14006
rect 23112 13942 23164 13948
rect 23020 13932 23072 13938
rect 23020 13874 23072 13880
rect 23032 13818 23060 13874
rect 23032 13790 23152 13818
rect 22928 13320 22980 13326
rect 22928 13262 22980 13268
rect 22940 12850 22968 13262
rect 23124 12850 23152 13790
rect 23234 13084 23542 13093
rect 23234 13082 23240 13084
rect 23296 13082 23320 13084
rect 23376 13082 23400 13084
rect 23456 13082 23480 13084
rect 23536 13082 23542 13084
rect 23296 13030 23298 13082
rect 23478 13030 23480 13082
rect 23234 13028 23240 13030
rect 23296 13028 23320 13030
rect 23376 13028 23400 13030
rect 23456 13028 23480 13030
rect 23536 13028 23542 13030
rect 23234 13019 23542 13028
rect 22928 12844 22980 12850
rect 22928 12786 22980 12792
rect 23112 12844 23164 12850
rect 23112 12786 23164 12792
rect 22468 12640 22520 12646
rect 22468 12582 22520 12588
rect 22480 12306 22508 12582
rect 22468 12300 22520 12306
rect 22468 12242 22520 12248
rect 22928 12300 22980 12306
rect 22928 12242 22980 12248
rect 22940 11762 22968 12242
rect 22928 11756 22980 11762
rect 22928 11698 22980 11704
rect 23020 11756 23072 11762
rect 23020 11698 23072 11704
rect 21928 11614 22048 11642
rect 21732 11552 21784 11558
rect 21732 11494 21784 11500
rect 20444 11348 20496 11354
rect 20444 11290 20496 11296
rect 19812 11218 19932 11234
rect 21744 11218 21772 11494
rect 19432 11212 19484 11218
rect 19432 11154 19484 11160
rect 19800 11212 19932 11218
rect 19852 11206 19932 11212
rect 21732 11212 21784 11218
rect 19800 11154 19852 11160
rect 21732 11154 21784 11160
rect 20720 11076 20772 11082
rect 20720 11018 20772 11024
rect 18604 11008 18656 11014
rect 18604 10950 18656 10956
rect 18616 10810 18644 10950
rect 18604 10804 18656 10810
rect 18604 10746 18656 10752
rect 20732 10742 20760 11018
rect 18144 10736 18196 10742
rect 18144 10678 18196 10684
rect 20720 10736 20772 10742
rect 20720 10678 20772 10684
rect 17960 10124 18012 10130
rect 17960 10066 18012 10072
rect 17592 10056 17644 10062
rect 17592 9998 17644 10004
rect 17604 9586 17632 9998
rect 17592 9580 17644 9586
rect 17592 9522 17644 9528
rect 18156 9518 18184 10678
rect 19984 10668 20036 10674
rect 19984 10610 20036 10616
rect 19520 10364 19828 10373
rect 19520 10362 19526 10364
rect 19582 10362 19606 10364
rect 19662 10362 19686 10364
rect 19742 10362 19766 10364
rect 19822 10362 19828 10364
rect 19582 10310 19584 10362
rect 19764 10310 19766 10362
rect 19520 10308 19526 10310
rect 19582 10308 19606 10310
rect 19662 10308 19686 10310
rect 19742 10308 19766 10310
rect 19822 10308 19828 10310
rect 19520 10299 19828 10308
rect 19996 10266 20024 10610
rect 19984 10260 20036 10266
rect 19984 10202 20036 10208
rect 21928 9586 21956 11614
rect 22008 11552 22060 11558
rect 22008 11494 22060 11500
rect 22020 11218 22048 11494
rect 22008 11212 22060 11218
rect 22008 11154 22060 11160
rect 22940 10606 22968 11698
rect 23032 10674 23060 11698
rect 23124 11626 23152 12786
rect 23480 12640 23532 12646
rect 23480 12582 23532 12588
rect 23492 12442 23520 12582
rect 23480 12436 23532 12442
rect 23480 12378 23532 12384
rect 23234 11996 23542 12005
rect 23234 11994 23240 11996
rect 23296 11994 23320 11996
rect 23376 11994 23400 11996
rect 23456 11994 23480 11996
rect 23536 11994 23542 11996
rect 23296 11942 23298 11994
rect 23478 11942 23480 11994
rect 23234 11940 23240 11942
rect 23296 11940 23320 11942
rect 23376 11940 23400 11942
rect 23456 11940 23480 11942
rect 23536 11940 23542 11942
rect 23234 11931 23542 11940
rect 23112 11620 23164 11626
rect 23112 11562 23164 11568
rect 23124 11354 23152 11562
rect 23112 11348 23164 11354
rect 23112 11290 23164 11296
rect 23676 11218 23704 15030
rect 23768 14278 23796 15438
rect 24412 14482 24440 16050
rect 24860 15904 24912 15910
rect 24860 15846 24912 15852
rect 24872 15502 24900 15846
rect 24860 15496 24912 15502
rect 24860 15438 24912 15444
rect 24584 15360 24636 15366
rect 24584 15302 24636 15308
rect 24596 15162 24624 15302
rect 24584 15156 24636 15162
rect 24584 15098 24636 15104
rect 24596 14482 24624 15098
rect 24400 14476 24452 14482
rect 24400 14418 24452 14424
rect 24584 14476 24636 14482
rect 24584 14418 24636 14424
rect 24768 14408 24820 14414
rect 24768 14350 24820 14356
rect 23756 14272 23808 14278
rect 23756 14214 23808 14220
rect 24780 13802 24808 14350
rect 24768 13796 24820 13802
rect 24768 13738 24820 13744
rect 24584 13728 24636 13734
rect 24584 13670 24636 13676
rect 24596 13258 24624 13670
rect 24780 13326 24808 13738
rect 24964 13734 24992 16934
rect 24952 13728 25004 13734
rect 24952 13670 25004 13676
rect 24768 13320 24820 13326
rect 24768 13262 24820 13268
rect 24584 13252 24636 13258
rect 24584 13194 24636 13200
rect 23940 12776 23992 12782
rect 23940 12718 23992 12724
rect 23952 12442 23980 12718
rect 23940 12436 23992 12442
rect 23940 12378 23992 12384
rect 23756 12164 23808 12170
rect 23756 12106 23808 12112
rect 23768 11830 23796 12106
rect 23756 11824 23808 11830
rect 23756 11766 23808 11772
rect 23664 11212 23716 11218
rect 23664 11154 23716 11160
rect 23112 11144 23164 11150
rect 23112 11086 23164 11092
rect 23124 10742 23152 11086
rect 23234 10908 23542 10917
rect 23234 10906 23240 10908
rect 23296 10906 23320 10908
rect 23376 10906 23400 10908
rect 23456 10906 23480 10908
rect 23536 10906 23542 10908
rect 23296 10854 23298 10906
rect 23478 10854 23480 10906
rect 23234 10852 23240 10854
rect 23296 10852 23320 10854
rect 23376 10852 23400 10854
rect 23456 10852 23480 10854
rect 23536 10852 23542 10854
rect 23234 10843 23542 10852
rect 23112 10736 23164 10742
rect 23112 10678 23164 10684
rect 23020 10668 23072 10674
rect 23020 10610 23072 10616
rect 22928 10600 22980 10606
rect 22928 10542 22980 10548
rect 23032 10266 23060 10610
rect 23020 10260 23072 10266
rect 23020 10202 23072 10208
rect 24596 10062 24624 13194
rect 25044 13184 25096 13190
rect 25044 13126 25096 13132
rect 25056 12918 25084 13126
rect 25044 12912 25096 12918
rect 25044 12854 25096 12860
rect 25044 12640 25096 12646
rect 25044 12582 25096 12588
rect 24768 11212 24820 11218
rect 24768 11154 24820 11160
rect 24676 11144 24728 11150
rect 24676 11086 24728 11092
rect 24584 10056 24636 10062
rect 24584 9998 24636 10004
rect 23234 9820 23542 9829
rect 23234 9818 23240 9820
rect 23296 9818 23320 9820
rect 23376 9818 23400 9820
rect 23456 9818 23480 9820
rect 23536 9818 23542 9820
rect 23296 9766 23298 9818
rect 23478 9766 23480 9818
rect 23234 9764 23240 9766
rect 23296 9764 23320 9766
rect 23376 9764 23400 9766
rect 23456 9764 23480 9766
rect 23536 9764 23542 9766
rect 23234 9755 23542 9764
rect 21916 9580 21968 9586
rect 21916 9522 21968 9528
rect 22836 9580 22888 9586
rect 22836 9522 22888 9528
rect 18144 9512 18196 9518
rect 18144 9454 18196 9460
rect 19520 9276 19828 9285
rect 19520 9274 19526 9276
rect 19582 9274 19606 9276
rect 19662 9274 19686 9276
rect 19742 9274 19766 9276
rect 19822 9274 19828 9276
rect 19582 9222 19584 9274
rect 19764 9222 19766 9274
rect 19520 9220 19526 9222
rect 19582 9220 19606 9222
rect 19662 9220 19686 9222
rect 19742 9220 19766 9222
rect 19822 9220 19828 9222
rect 19520 9211 19828 9220
rect 22848 9178 22876 9522
rect 23848 9376 23900 9382
rect 23848 9318 23900 9324
rect 22836 9172 22888 9178
rect 22836 9114 22888 9120
rect 23860 8974 23888 9318
rect 24688 8974 24716 11086
rect 24780 10674 24808 11154
rect 24860 11008 24912 11014
rect 24860 10950 24912 10956
rect 24872 10810 24900 10950
rect 24860 10804 24912 10810
rect 24860 10746 24912 10752
rect 24768 10668 24820 10674
rect 24768 10610 24820 10616
rect 24780 9722 24808 10610
rect 25056 10062 25084 12582
rect 25424 11218 25452 18158
rect 26948 17980 27256 17989
rect 26948 17978 26954 17980
rect 27010 17978 27034 17980
rect 27090 17978 27114 17980
rect 27170 17978 27194 17980
rect 27250 17978 27256 17980
rect 27010 17926 27012 17978
rect 27192 17926 27194 17978
rect 26948 17924 26954 17926
rect 27010 17924 27034 17926
rect 27090 17924 27114 17926
rect 27170 17924 27194 17926
rect 27250 17924 27256 17926
rect 26948 17915 27256 17924
rect 27620 17672 27672 17678
rect 27620 17614 27672 17620
rect 26424 17536 26476 17542
rect 26424 17478 26476 17484
rect 26148 16992 26200 16998
rect 26148 16934 26200 16940
rect 26160 16658 26188 16934
rect 26436 16658 26464 17478
rect 27632 17338 27660 17614
rect 27620 17332 27672 17338
rect 27620 17274 27672 17280
rect 27436 17264 27488 17270
rect 27436 17206 27488 17212
rect 26948 16892 27256 16901
rect 26948 16890 26954 16892
rect 27010 16890 27034 16892
rect 27090 16890 27114 16892
rect 27170 16890 27194 16892
rect 27250 16890 27256 16892
rect 27010 16838 27012 16890
rect 27192 16838 27194 16890
rect 26948 16836 26954 16838
rect 27010 16836 27034 16838
rect 27090 16836 27114 16838
rect 27170 16836 27194 16838
rect 27250 16836 27256 16838
rect 26948 16827 27256 16836
rect 26148 16652 26200 16658
rect 26148 16594 26200 16600
rect 26424 16652 26476 16658
rect 26424 16594 26476 16600
rect 27448 16522 27476 17206
rect 27632 16794 27660 17274
rect 28356 17196 28408 17202
rect 28356 17138 28408 17144
rect 27896 17128 27948 17134
rect 27896 17070 27948 17076
rect 27988 17128 28040 17134
rect 27988 17070 28040 17076
rect 27620 16788 27672 16794
rect 27620 16730 27672 16736
rect 27908 16590 27936 17070
rect 27896 16584 27948 16590
rect 27896 16526 27948 16532
rect 27436 16516 27488 16522
rect 27436 16458 27488 16464
rect 25964 16040 26016 16046
rect 25964 15982 26016 15988
rect 25976 15706 26004 15982
rect 26948 15804 27256 15813
rect 26948 15802 26954 15804
rect 27010 15802 27034 15804
rect 27090 15802 27114 15804
rect 27170 15802 27194 15804
rect 27250 15802 27256 15804
rect 27010 15750 27012 15802
rect 27192 15750 27194 15802
rect 26948 15748 26954 15750
rect 27010 15748 27034 15750
rect 27090 15748 27114 15750
rect 27170 15748 27194 15750
rect 27250 15748 27256 15750
rect 26948 15739 27256 15748
rect 25964 15700 26016 15706
rect 25964 15642 26016 15648
rect 25976 14958 26004 15642
rect 28000 15502 28028 17070
rect 28264 16584 28316 16590
rect 28264 16526 28316 16532
rect 28276 16250 28304 16526
rect 28264 16244 28316 16250
rect 28264 16186 28316 16192
rect 28368 15502 28396 17138
rect 29736 17128 29788 17134
rect 29736 17070 29788 17076
rect 29644 16584 29696 16590
rect 29644 16526 29696 16532
rect 28724 16448 28776 16454
rect 28724 16390 28776 16396
rect 28736 16046 28764 16390
rect 28724 16040 28776 16046
rect 28724 15982 28776 15988
rect 29656 15570 29684 16526
rect 29748 16182 29776 17070
rect 29736 16176 29788 16182
rect 29736 16118 29788 16124
rect 29644 15564 29696 15570
rect 29644 15506 29696 15512
rect 27988 15496 28040 15502
rect 27988 15438 28040 15444
rect 28356 15496 28408 15502
rect 28356 15438 28408 15444
rect 27804 15020 27856 15026
rect 27804 14962 27856 14968
rect 25964 14952 26016 14958
rect 25964 14894 26016 14900
rect 25872 14816 25924 14822
rect 25872 14758 25924 14764
rect 25596 14476 25648 14482
rect 25596 14418 25648 14424
rect 25608 14006 25636 14418
rect 25688 14340 25740 14346
rect 25688 14282 25740 14288
rect 25596 14000 25648 14006
rect 25596 13942 25648 13948
rect 25412 11212 25464 11218
rect 25412 11154 25464 11160
rect 25320 11008 25372 11014
rect 25320 10950 25372 10956
rect 25332 10742 25360 10950
rect 25320 10736 25372 10742
rect 25320 10678 25372 10684
rect 25424 10130 25452 11154
rect 25700 11150 25728 14282
rect 25884 13938 25912 14758
rect 26948 14716 27256 14725
rect 26948 14714 26954 14716
rect 27010 14714 27034 14716
rect 27090 14714 27114 14716
rect 27170 14714 27194 14716
rect 27250 14714 27256 14716
rect 27010 14662 27012 14714
rect 27192 14662 27194 14714
rect 26948 14660 26954 14662
rect 27010 14660 27034 14662
rect 27090 14660 27114 14662
rect 27170 14660 27194 14662
rect 27250 14660 27256 14662
rect 26948 14651 27256 14660
rect 27816 14414 27844 14962
rect 27896 14952 27948 14958
rect 27896 14894 27948 14900
rect 27908 14618 27936 14894
rect 27896 14612 27948 14618
rect 27896 14554 27948 14560
rect 27804 14408 27856 14414
rect 27804 14350 27856 14356
rect 27528 14272 27580 14278
rect 27528 14214 27580 14220
rect 25872 13932 25924 13938
rect 25872 13874 25924 13880
rect 26516 13932 26568 13938
rect 26516 13874 26568 13880
rect 26056 13184 26108 13190
rect 26056 13126 26108 13132
rect 26068 12986 26096 13126
rect 26056 12980 26108 12986
rect 26056 12922 26108 12928
rect 26068 12238 26096 12922
rect 26148 12844 26200 12850
rect 26148 12786 26200 12792
rect 26160 12306 26188 12786
rect 26528 12782 26556 13874
rect 27344 13728 27396 13734
rect 27344 13670 27396 13676
rect 26948 13628 27256 13637
rect 26948 13626 26954 13628
rect 27010 13626 27034 13628
rect 27090 13626 27114 13628
rect 27170 13626 27194 13628
rect 27250 13626 27256 13628
rect 27010 13574 27012 13626
rect 27192 13574 27194 13626
rect 26948 13572 26954 13574
rect 27010 13572 27034 13574
rect 27090 13572 27114 13574
rect 27170 13572 27194 13574
rect 27250 13572 27256 13574
rect 26948 13563 27256 13572
rect 27356 13394 27384 13670
rect 27344 13388 27396 13394
rect 27344 13330 27396 13336
rect 27540 13258 27568 14214
rect 27528 13252 27580 13258
rect 27528 13194 27580 13200
rect 27436 12844 27488 12850
rect 27436 12786 27488 12792
rect 26516 12776 26568 12782
rect 26516 12718 26568 12724
rect 26948 12540 27256 12549
rect 26948 12538 26954 12540
rect 27010 12538 27034 12540
rect 27090 12538 27114 12540
rect 27170 12538 27194 12540
rect 27250 12538 27256 12540
rect 27010 12486 27012 12538
rect 27192 12486 27194 12538
rect 26948 12484 26954 12486
rect 27010 12484 27034 12486
rect 27090 12484 27114 12486
rect 27170 12484 27194 12486
rect 27250 12484 27256 12486
rect 26948 12475 27256 12484
rect 27448 12374 27476 12786
rect 28000 12782 28028 15438
rect 28172 15360 28224 15366
rect 28172 15302 28224 15308
rect 28184 15094 28212 15302
rect 28172 15088 28224 15094
rect 28172 15030 28224 15036
rect 28264 13252 28316 13258
rect 28264 13194 28316 13200
rect 28276 12918 28304 13194
rect 28264 12912 28316 12918
rect 28264 12854 28316 12860
rect 28368 12850 28396 15438
rect 29184 15428 29236 15434
rect 29184 15370 29236 15376
rect 29196 15094 29224 15370
rect 29656 15162 29684 15506
rect 29644 15156 29696 15162
rect 29644 15098 29696 15104
rect 29184 15088 29236 15094
rect 29184 15030 29236 15036
rect 28724 14408 28776 14414
rect 28724 14350 28776 14356
rect 28632 14272 28684 14278
rect 28632 14214 28684 14220
rect 28644 14006 28672 14214
rect 28632 14000 28684 14006
rect 28632 13942 28684 13948
rect 28632 13864 28684 13870
rect 28632 13806 28684 13812
rect 28644 13530 28672 13806
rect 28632 13524 28684 13530
rect 28632 13466 28684 13472
rect 28736 13462 28764 14350
rect 29644 14340 29696 14346
rect 29644 14282 29696 14288
rect 29656 14074 29684 14282
rect 29644 14068 29696 14074
rect 29644 14010 29696 14016
rect 28724 13456 28776 13462
rect 28724 13398 28776 13404
rect 29656 13326 29684 14010
rect 29736 13932 29788 13938
rect 29736 13874 29788 13880
rect 29644 13320 29696 13326
rect 29644 13262 29696 13268
rect 29748 12918 29776 13874
rect 29736 12912 29788 12918
rect 29736 12854 29788 12860
rect 28356 12844 28408 12850
rect 28356 12786 28408 12792
rect 27988 12776 28040 12782
rect 27988 12718 28040 12724
rect 27436 12368 27488 12374
rect 27436 12310 27488 12316
rect 26148 12300 26200 12306
rect 26148 12242 26200 12248
rect 26056 12232 26108 12238
rect 26056 12174 26108 12180
rect 26948 11452 27256 11461
rect 26948 11450 26954 11452
rect 27010 11450 27034 11452
rect 27090 11450 27114 11452
rect 27170 11450 27194 11452
rect 27250 11450 27256 11452
rect 27010 11398 27012 11450
rect 27192 11398 27194 11450
rect 26948 11396 26954 11398
rect 27010 11396 27034 11398
rect 27090 11396 27114 11398
rect 27170 11396 27194 11398
rect 27250 11396 27256 11398
rect 26948 11387 27256 11396
rect 29000 11280 29052 11286
rect 29000 11222 29052 11228
rect 25688 11144 25740 11150
rect 25688 11086 25740 11092
rect 26516 11076 26568 11082
rect 26516 11018 26568 11024
rect 28724 11076 28776 11082
rect 28724 11018 28776 11024
rect 26528 10606 26556 11018
rect 27436 10736 27488 10742
rect 27436 10678 27488 10684
rect 27988 10736 28040 10742
rect 27988 10678 28040 10684
rect 26516 10600 26568 10606
rect 26516 10542 26568 10548
rect 26948 10364 27256 10373
rect 26948 10362 26954 10364
rect 27010 10362 27034 10364
rect 27090 10362 27114 10364
rect 27170 10362 27194 10364
rect 27250 10362 27256 10364
rect 27010 10310 27012 10362
rect 27192 10310 27194 10362
rect 26948 10308 26954 10310
rect 27010 10308 27034 10310
rect 27090 10308 27114 10310
rect 27170 10308 27194 10310
rect 27250 10308 27256 10310
rect 26948 10299 27256 10308
rect 25412 10124 25464 10130
rect 25412 10066 25464 10072
rect 25044 10056 25096 10062
rect 25044 9998 25096 10004
rect 27448 9926 27476 10678
rect 27712 10600 27764 10606
rect 27712 10542 27764 10548
rect 27724 9994 27752 10542
rect 28000 10062 28028 10678
rect 28736 10674 28764 11018
rect 29012 10742 29040 11222
rect 29828 11212 29880 11218
rect 29828 11154 29880 11160
rect 29840 10810 29868 11154
rect 29828 10804 29880 10810
rect 29828 10746 29880 10752
rect 29932 10742 29960 18770
rect 30662 18524 30970 18533
rect 30662 18522 30668 18524
rect 30724 18522 30748 18524
rect 30804 18522 30828 18524
rect 30884 18522 30908 18524
rect 30964 18522 30970 18524
rect 30724 18470 30726 18522
rect 30906 18470 30908 18522
rect 30662 18468 30668 18470
rect 30724 18468 30748 18470
rect 30804 18468 30828 18470
rect 30884 18468 30908 18470
rect 30964 18468 30970 18470
rect 30662 18459 30970 18468
rect 31024 18216 31076 18222
rect 31024 18158 31076 18164
rect 31036 17921 31064 18158
rect 31022 17912 31078 17921
rect 31022 17847 31078 17856
rect 30662 17436 30970 17445
rect 30662 17434 30668 17436
rect 30724 17434 30748 17436
rect 30804 17434 30828 17436
rect 30884 17434 30908 17436
rect 30964 17434 30970 17436
rect 30724 17382 30726 17434
rect 30906 17382 30908 17434
rect 30662 17380 30668 17382
rect 30724 17380 30748 17382
rect 30804 17380 30828 17382
rect 30884 17380 30908 17382
rect 30964 17380 30970 17382
rect 30662 17371 30970 17380
rect 30012 16448 30064 16454
rect 30012 16390 30064 16396
rect 30024 16114 30052 16390
rect 30662 16348 30970 16357
rect 30662 16346 30668 16348
rect 30724 16346 30748 16348
rect 30804 16346 30828 16348
rect 30884 16346 30908 16348
rect 30964 16346 30970 16348
rect 30724 16294 30726 16346
rect 30906 16294 30908 16346
rect 30662 16292 30668 16294
rect 30724 16292 30748 16294
rect 30804 16292 30828 16294
rect 30884 16292 30908 16294
rect 30964 16292 30970 16294
rect 30662 16283 30970 16292
rect 30012 16108 30064 16114
rect 30012 16050 30064 16056
rect 30662 15260 30970 15269
rect 30662 15258 30668 15260
rect 30724 15258 30748 15260
rect 30804 15258 30828 15260
rect 30884 15258 30908 15260
rect 30964 15258 30970 15260
rect 30724 15206 30726 15258
rect 30906 15206 30908 15258
rect 30662 15204 30668 15206
rect 30724 15204 30748 15206
rect 30804 15204 30828 15206
rect 30884 15204 30908 15206
rect 30964 15204 30970 15206
rect 30662 15195 30970 15204
rect 30288 14408 30340 14414
rect 30288 14350 30340 14356
rect 30300 11286 30328 14350
rect 31024 14340 31076 14346
rect 31024 14282 31076 14288
rect 30662 14172 30970 14181
rect 30662 14170 30668 14172
rect 30724 14170 30748 14172
rect 30804 14170 30828 14172
rect 30884 14170 30908 14172
rect 30964 14170 30970 14172
rect 30724 14118 30726 14170
rect 30906 14118 30908 14170
rect 30662 14116 30668 14118
rect 30724 14116 30748 14118
rect 30804 14116 30828 14118
rect 30884 14116 30908 14118
rect 30964 14116 30970 14118
rect 30662 14107 30970 14116
rect 31036 13977 31064 14282
rect 31022 13968 31078 13977
rect 31022 13903 31078 13912
rect 30662 13084 30970 13093
rect 30662 13082 30668 13084
rect 30724 13082 30748 13084
rect 30804 13082 30828 13084
rect 30884 13082 30908 13084
rect 30964 13082 30970 13084
rect 30724 13030 30726 13082
rect 30906 13030 30908 13082
rect 30662 13028 30668 13030
rect 30724 13028 30748 13030
rect 30804 13028 30828 13030
rect 30884 13028 30908 13030
rect 30964 13028 30970 13030
rect 30662 13019 30970 13028
rect 30662 11996 30970 12005
rect 30662 11994 30668 11996
rect 30724 11994 30748 11996
rect 30804 11994 30828 11996
rect 30884 11994 30908 11996
rect 30964 11994 30970 11996
rect 30724 11942 30726 11994
rect 30906 11942 30908 11994
rect 30662 11940 30668 11942
rect 30724 11940 30748 11942
rect 30804 11940 30828 11942
rect 30884 11940 30908 11942
rect 30964 11940 30970 11942
rect 30662 11931 30970 11940
rect 30288 11280 30340 11286
rect 30288 11222 30340 11228
rect 30662 10908 30970 10917
rect 30662 10906 30668 10908
rect 30724 10906 30748 10908
rect 30804 10906 30828 10908
rect 30884 10906 30908 10908
rect 30964 10906 30970 10908
rect 30724 10854 30726 10906
rect 30906 10854 30908 10906
rect 30662 10852 30668 10854
rect 30724 10852 30748 10854
rect 30804 10852 30828 10854
rect 30884 10852 30908 10854
rect 30964 10852 30970 10854
rect 30662 10843 30970 10852
rect 29000 10736 29052 10742
rect 29000 10678 29052 10684
rect 29920 10736 29972 10742
rect 29920 10678 29972 10684
rect 28172 10668 28224 10674
rect 28172 10610 28224 10616
rect 28724 10668 28776 10674
rect 28724 10610 28776 10616
rect 28908 10668 28960 10674
rect 28908 10610 28960 10616
rect 28184 10062 28212 10610
rect 28736 10266 28764 10610
rect 28724 10260 28776 10266
rect 28724 10202 28776 10208
rect 27988 10056 28040 10062
rect 27908 10004 27988 10010
rect 27908 9998 28040 10004
rect 28172 10056 28224 10062
rect 28172 9998 28224 10004
rect 27712 9988 27764 9994
rect 27712 9930 27764 9936
rect 27908 9982 28028 9998
rect 24860 9920 24912 9926
rect 24860 9862 24912 9868
rect 26056 9920 26108 9926
rect 26056 9862 26108 9868
rect 27436 9920 27488 9926
rect 27436 9862 27488 9868
rect 24768 9716 24820 9722
rect 24768 9658 24820 9664
rect 24780 8974 24808 9658
rect 24872 9654 24900 9862
rect 26068 9722 26096 9862
rect 26056 9716 26108 9722
rect 26056 9658 26108 9664
rect 24860 9648 24912 9654
rect 24860 9590 24912 9596
rect 25044 9648 25096 9654
rect 25044 9590 25096 9596
rect 25056 9178 25084 9590
rect 26948 9276 27256 9285
rect 26948 9274 26954 9276
rect 27010 9274 27034 9276
rect 27090 9274 27114 9276
rect 27170 9274 27194 9276
rect 27250 9274 27256 9276
rect 27010 9222 27012 9274
rect 27192 9222 27194 9274
rect 26948 9220 26954 9222
rect 27010 9220 27034 9222
rect 27090 9220 27114 9222
rect 27170 9220 27194 9222
rect 27250 9220 27256 9222
rect 26948 9211 27256 9220
rect 25044 9172 25096 9178
rect 25044 9114 25096 9120
rect 19892 8968 19944 8974
rect 19892 8910 19944 8916
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 23848 8968 23900 8974
rect 23848 8910 23900 8916
rect 24676 8968 24728 8974
rect 24676 8910 24728 8916
rect 24768 8968 24820 8974
rect 24768 8910 24820 8916
rect 19064 8628 19116 8634
rect 19064 8570 19116 8576
rect 19432 8628 19484 8634
rect 19432 8570 19484 8576
rect 19076 8514 19104 8570
rect 19076 8498 19196 8514
rect 19076 8492 19208 8498
rect 19076 8486 19156 8492
rect 19156 8434 19208 8440
rect 17132 8424 17184 8430
rect 17132 8366 17184 8372
rect 18972 8424 19024 8430
rect 18972 8366 19024 8372
rect 17144 8090 17172 8366
rect 18604 8288 18656 8294
rect 18604 8230 18656 8236
rect 17132 8084 17184 8090
rect 17132 8026 17184 8032
rect 18616 7954 18644 8230
rect 18984 7954 19012 8366
rect 19444 8090 19472 8570
rect 19520 8188 19828 8197
rect 19520 8186 19526 8188
rect 19582 8186 19606 8188
rect 19662 8186 19686 8188
rect 19742 8186 19766 8188
rect 19822 8186 19828 8188
rect 19582 8134 19584 8186
rect 19764 8134 19766 8186
rect 19520 8132 19526 8134
rect 19582 8132 19606 8134
rect 19662 8132 19686 8134
rect 19742 8132 19766 8134
rect 19822 8132 19828 8134
rect 19520 8123 19828 8132
rect 19432 8084 19484 8090
rect 19432 8026 19484 8032
rect 18604 7948 18656 7954
rect 18604 7890 18656 7896
rect 18972 7948 19024 7954
rect 18972 7890 19024 7896
rect 18512 7880 18564 7886
rect 18512 7822 18564 7828
rect 17408 7812 17460 7818
rect 17408 7754 17460 7760
rect 16672 7404 16724 7410
rect 16672 7346 16724 7352
rect 16764 7404 16816 7410
rect 16764 7346 16816 7352
rect 16684 6798 16712 7346
rect 16776 6914 16804 7346
rect 17132 7336 17184 7342
rect 17132 7278 17184 7284
rect 16776 6886 16896 6914
rect 16672 6792 16724 6798
rect 16672 6734 16724 6740
rect 16488 6724 16540 6730
rect 16488 6666 16540 6672
rect 16868 6662 16896 6886
rect 17144 6866 17172 7278
rect 17420 6866 17448 7754
rect 17684 7744 17736 7750
rect 17684 7686 17736 7692
rect 17500 7336 17552 7342
rect 17500 7278 17552 7284
rect 17132 6860 17184 6866
rect 17132 6802 17184 6808
rect 17408 6860 17460 6866
rect 17408 6802 17460 6808
rect 17512 6798 17540 7278
rect 17696 7206 17724 7686
rect 18524 7546 18552 7822
rect 18512 7540 18564 7546
rect 18512 7482 18564 7488
rect 17684 7200 17736 7206
rect 17684 7142 17736 7148
rect 17696 6798 17724 7142
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 17684 6792 17736 6798
rect 17684 6734 17736 6740
rect 16856 6656 16908 6662
rect 16856 6598 16908 6604
rect 15806 6556 16114 6565
rect 15806 6554 15812 6556
rect 15868 6554 15892 6556
rect 15948 6554 15972 6556
rect 16028 6554 16052 6556
rect 16108 6554 16114 6556
rect 15868 6502 15870 6554
rect 16050 6502 16052 6554
rect 15806 6500 15812 6502
rect 15868 6500 15892 6502
rect 15948 6500 15972 6502
rect 16028 6500 16052 6502
rect 16108 6500 16114 6502
rect 15806 6491 16114 6500
rect 14648 5908 14700 5914
rect 14648 5850 14700 5856
rect 16868 5778 16896 6598
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 17960 5568 18012 5574
rect 17960 5510 18012 5516
rect 15806 5468 16114 5477
rect 15806 5466 15812 5468
rect 15868 5466 15892 5468
rect 15948 5466 15972 5468
rect 16028 5466 16052 5468
rect 16108 5466 16114 5468
rect 15868 5414 15870 5466
rect 16050 5414 16052 5466
rect 15806 5412 15812 5414
rect 15868 5412 15892 5414
rect 15948 5412 15972 5414
rect 16028 5412 16052 5414
rect 16108 5412 16114 5414
rect 15806 5403 16114 5412
rect 14556 5228 14608 5234
rect 14556 5170 14608 5176
rect 17224 5228 17276 5234
rect 17224 5170 17276 5176
rect 14372 5160 14424 5166
rect 14372 5102 14424 5108
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 4664 4924 4972 4933
rect 4664 4922 4670 4924
rect 4726 4922 4750 4924
rect 4806 4922 4830 4924
rect 4886 4922 4910 4924
rect 4966 4922 4972 4924
rect 4726 4870 4728 4922
rect 4908 4870 4910 4922
rect 4664 4868 4670 4870
rect 4726 4868 4750 4870
rect 4806 4868 4830 4870
rect 4886 4868 4910 4870
rect 4966 4868 4972 4870
rect 4664 4859 4972 4868
rect 12092 4924 12400 4933
rect 12092 4922 12098 4924
rect 12154 4922 12178 4924
rect 12234 4922 12258 4924
rect 12314 4922 12338 4924
rect 12394 4922 12400 4924
rect 12154 4870 12156 4922
rect 12336 4870 12338 4922
rect 12092 4868 12098 4870
rect 12154 4868 12178 4870
rect 12234 4868 12258 4870
rect 12314 4868 12338 4870
rect 12394 4868 12400 4870
rect 12092 4859 12400 4868
rect 8378 4380 8686 4389
rect 8378 4378 8384 4380
rect 8440 4378 8464 4380
rect 8520 4378 8544 4380
rect 8600 4378 8624 4380
rect 8680 4378 8686 4380
rect 8440 4326 8442 4378
rect 8622 4326 8624 4378
rect 8378 4324 8384 4326
rect 8440 4324 8464 4326
rect 8520 4324 8544 4326
rect 8600 4324 8624 4326
rect 8680 4324 8686 4326
rect 8378 4315 8686 4324
rect 14016 4146 14044 4966
rect 14384 4758 14412 5102
rect 14372 4752 14424 4758
rect 14372 4694 14424 4700
rect 14384 4214 14412 4694
rect 14568 4622 14596 5170
rect 17236 4826 17264 5170
rect 17224 4820 17276 4826
rect 17224 4762 17276 4768
rect 14648 4684 14700 4690
rect 14648 4626 14700 4632
rect 14556 4616 14608 4622
rect 14556 4558 14608 4564
rect 14660 4282 14688 4626
rect 17972 4622 18000 5510
rect 18616 5234 18644 7890
rect 19904 7886 19932 8910
rect 19984 8832 20036 8838
rect 19984 8774 20036 8780
rect 19996 8566 20024 8774
rect 19984 8560 20036 8566
rect 19984 8502 20036 8508
rect 21468 8498 21496 8910
rect 22284 8900 22336 8906
rect 22284 8842 22336 8848
rect 22296 8498 22324 8842
rect 23234 8732 23542 8741
rect 23234 8730 23240 8732
rect 23296 8730 23320 8732
rect 23376 8730 23400 8732
rect 23456 8730 23480 8732
rect 23536 8730 23542 8732
rect 23296 8678 23298 8730
rect 23478 8678 23480 8730
rect 23234 8676 23240 8678
rect 23296 8676 23320 8678
rect 23376 8676 23400 8678
rect 23456 8676 23480 8678
rect 23536 8676 23542 8678
rect 23234 8667 23542 8676
rect 23860 8498 23888 8910
rect 24780 8566 24808 8910
rect 27448 8634 27476 9862
rect 27528 8968 27580 8974
rect 27528 8910 27580 8916
rect 27436 8628 27488 8634
rect 27436 8570 27488 8576
rect 27540 8566 27568 8910
rect 27724 8906 27752 9930
rect 27908 9654 27936 9982
rect 28184 9722 28212 9998
rect 28172 9716 28224 9722
rect 28172 9658 28224 9664
rect 27896 9648 27948 9654
rect 27896 9590 27948 9596
rect 27712 8900 27764 8906
rect 27712 8842 27764 8848
rect 27804 8900 27856 8906
rect 27804 8842 27856 8848
rect 24768 8560 24820 8566
rect 24768 8502 24820 8508
rect 27528 8560 27580 8566
rect 27528 8502 27580 8508
rect 21456 8492 21508 8498
rect 21456 8434 21508 8440
rect 22284 8492 22336 8498
rect 22284 8434 22336 8440
rect 23848 8492 23900 8498
rect 23848 8434 23900 8440
rect 20812 8288 20864 8294
rect 20812 8230 20864 8236
rect 20824 7954 20852 8230
rect 20812 7948 20864 7954
rect 20812 7890 20864 7896
rect 19616 7880 19668 7886
rect 19616 7822 19668 7828
rect 19892 7880 19944 7886
rect 19892 7822 19944 7828
rect 20444 7880 20496 7886
rect 20444 7822 20496 7828
rect 19628 7342 19656 7822
rect 19616 7336 19668 7342
rect 19616 7278 19668 7284
rect 19520 7100 19828 7109
rect 19520 7098 19526 7100
rect 19582 7098 19606 7100
rect 19662 7098 19686 7100
rect 19742 7098 19766 7100
rect 19822 7098 19828 7100
rect 19582 7046 19584 7098
rect 19764 7046 19766 7098
rect 19520 7044 19526 7046
rect 19582 7044 19606 7046
rect 19662 7044 19686 7046
rect 19742 7044 19766 7046
rect 19822 7044 19828 7046
rect 19520 7035 19828 7044
rect 20456 6866 20484 7822
rect 21468 7410 21496 8434
rect 22100 8288 22152 8294
rect 22100 8230 22152 8236
rect 22112 7818 22140 8230
rect 22100 7812 22152 7818
rect 22100 7754 22152 7760
rect 22192 7744 22244 7750
rect 22192 7686 22244 7692
rect 21456 7404 21508 7410
rect 21456 7346 21508 7352
rect 21364 7200 21416 7206
rect 21364 7142 21416 7148
rect 20444 6860 20496 6866
rect 20444 6802 20496 6808
rect 19520 6012 19828 6021
rect 19520 6010 19526 6012
rect 19582 6010 19606 6012
rect 19662 6010 19686 6012
rect 19742 6010 19766 6012
rect 19822 6010 19828 6012
rect 19582 5958 19584 6010
rect 19764 5958 19766 6010
rect 19520 5956 19526 5958
rect 19582 5956 19606 5958
rect 19662 5956 19686 5958
rect 19742 5956 19766 5958
rect 19822 5956 19828 5958
rect 19520 5947 19828 5956
rect 20456 5778 20484 6802
rect 21376 6730 21404 7142
rect 22204 6866 22232 7686
rect 22296 7478 22324 8434
rect 23860 7886 23888 8434
rect 26948 8188 27256 8197
rect 26948 8186 26954 8188
rect 27010 8186 27034 8188
rect 27090 8186 27114 8188
rect 27170 8186 27194 8188
rect 27250 8186 27256 8188
rect 27010 8134 27012 8186
rect 27192 8134 27194 8186
rect 26948 8132 26954 8134
rect 27010 8132 27034 8134
rect 27090 8132 27114 8134
rect 27170 8132 27194 8134
rect 27250 8132 27256 8134
rect 26948 8123 27256 8132
rect 27540 8090 27568 8502
rect 27724 8498 27752 8842
rect 27712 8492 27764 8498
rect 27712 8434 27764 8440
rect 27528 8084 27580 8090
rect 27528 8026 27580 8032
rect 23848 7880 23900 7886
rect 23848 7822 23900 7828
rect 24308 7880 24360 7886
rect 24308 7822 24360 7828
rect 23234 7644 23542 7653
rect 23234 7642 23240 7644
rect 23296 7642 23320 7644
rect 23376 7642 23400 7644
rect 23456 7642 23480 7644
rect 23536 7642 23542 7644
rect 23296 7590 23298 7642
rect 23478 7590 23480 7642
rect 23234 7588 23240 7590
rect 23296 7588 23320 7590
rect 23376 7588 23400 7590
rect 23456 7588 23480 7590
rect 23536 7588 23542 7590
rect 23234 7579 23542 7588
rect 22284 7472 22336 7478
rect 22284 7414 22336 7420
rect 22652 7200 22704 7206
rect 22652 7142 22704 7148
rect 22836 7200 22888 7206
rect 22836 7142 22888 7148
rect 22664 6914 22692 7142
rect 22664 6886 22784 6914
rect 22192 6860 22244 6866
rect 22192 6802 22244 6808
rect 21364 6724 21416 6730
rect 21364 6666 21416 6672
rect 22376 6656 22428 6662
rect 22376 6598 22428 6604
rect 22388 6322 22416 6598
rect 22756 6390 22784 6886
rect 22744 6384 22796 6390
rect 22744 6326 22796 6332
rect 22376 6316 22428 6322
rect 22376 6258 22428 6264
rect 21456 6248 21508 6254
rect 21456 6190 21508 6196
rect 21468 5778 21496 6190
rect 21732 6112 21784 6118
rect 21732 6054 21784 6060
rect 21744 5778 21772 6054
rect 19708 5772 19760 5778
rect 19708 5714 19760 5720
rect 19984 5772 20036 5778
rect 19984 5714 20036 5720
rect 20444 5772 20496 5778
rect 20444 5714 20496 5720
rect 20812 5772 20864 5778
rect 20812 5714 20864 5720
rect 21456 5772 21508 5778
rect 21456 5714 21508 5720
rect 21732 5772 21784 5778
rect 21732 5714 21784 5720
rect 19432 5636 19484 5642
rect 19432 5578 19484 5584
rect 18604 5228 18656 5234
rect 18604 5170 18656 5176
rect 19444 4826 19472 5578
rect 19720 5370 19748 5714
rect 19708 5364 19760 5370
rect 19708 5306 19760 5312
rect 19520 4924 19828 4933
rect 19520 4922 19526 4924
rect 19582 4922 19606 4924
rect 19662 4922 19686 4924
rect 19742 4922 19766 4924
rect 19822 4922 19828 4924
rect 19582 4870 19584 4922
rect 19764 4870 19766 4922
rect 19520 4868 19526 4870
rect 19582 4868 19606 4870
rect 19662 4868 19686 4870
rect 19742 4868 19766 4870
rect 19822 4868 19828 4870
rect 19520 4859 19828 4868
rect 19432 4820 19484 4826
rect 19432 4762 19484 4768
rect 19996 4622 20024 5714
rect 20824 4690 20852 5714
rect 22848 5710 22876 7142
rect 23234 6556 23542 6565
rect 23234 6554 23240 6556
rect 23296 6554 23320 6556
rect 23376 6554 23400 6556
rect 23456 6554 23480 6556
rect 23536 6554 23542 6556
rect 23296 6502 23298 6554
rect 23478 6502 23480 6554
rect 23234 6500 23240 6502
rect 23296 6500 23320 6502
rect 23376 6500 23400 6502
rect 23456 6500 23480 6502
rect 23536 6500 23542 6502
rect 23234 6491 23542 6500
rect 24320 6322 24348 7822
rect 25964 7404 26016 7410
rect 25964 7346 26016 7352
rect 27620 7404 27672 7410
rect 27620 7346 27672 7352
rect 25320 7200 25372 7206
rect 25320 7142 25372 7148
rect 25332 6798 25360 7142
rect 25976 7002 26004 7346
rect 26948 7100 27256 7109
rect 26948 7098 26954 7100
rect 27010 7098 27034 7100
rect 27090 7098 27114 7100
rect 27170 7098 27194 7100
rect 27250 7098 27256 7100
rect 27010 7046 27012 7098
rect 27192 7046 27194 7098
rect 26948 7044 26954 7046
rect 27010 7044 27034 7046
rect 27090 7044 27114 7046
rect 27170 7044 27194 7046
rect 27250 7044 27256 7046
rect 26948 7035 27256 7044
rect 25964 6996 26016 7002
rect 25964 6938 26016 6944
rect 25976 6798 26004 6938
rect 24584 6792 24636 6798
rect 24584 6734 24636 6740
rect 25320 6792 25372 6798
rect 25320 6734 25372 6740
rect 25964 6792 26016 6798
rect 25964 6734 26016 6740
rect 24596 6458 24624 6734
rect 24584 6452 24636 6458
rect 24584 6394 24636 6400
rect 25976 6322 26004 6734
rect 27344 6656 27396 6662
rect 27344 6598 27396 6604
rect 24308 6316 24360 6322
rect 24308 6258 24360 6264
rect 25964 6316 26016 6322
rect 25964 6258 26016 6264
rect 24320 5778 24348 6258
rect 24308 5772 24360 5778
rect 24308 5714 24360 5720
rect 25976 5710 26004 6258
rect 26948 6012 27256 6021
rect 26948 6010 26954 6012
rect 27010 6010 27034 6012
rect 27090 6010 27114 6012
rect 27170 6010 27194 6012
rect 27250 6010 27256 6012
rect 27010 5958 27012 6010
rect 27192 5958 27194 6010
rect 26948 5956 26954 5958
rect 27010 5956 27034 5958
rect 27090 5956 27114 5958
rect 27170 5956 27194 5958
rect 27250 5956 27256 5958
rect 26948 5947 27256 5956
rect 27356 5710 27384 6598
rect 27632 6458 27660 7346
rect 27724 6866 27752 8434
rect 27816 8430 27844 8842
rect 27908 8838 27936 9590
rect 28920 8974 28948 10610
rect 29736 10600 29788 10606
rect 29736 10542 29788 10548
rect 29748 10266 29776 10542
rect 29736 10260 29788 10266
rect 29736 10202 29788 10208
rect 30012 10192 30064 10198
rect 30012 10134 30064 10140
rect 29000 9920 29052 9926
rect 29000 9862 29052 9868
rect 29012 9654 29040 9862
rect 29000 9648 29052 9654
rect 29000 9590 29052 9596
rect 29828 9580 29880 9586
rect 29828 9522 29880 9528
rect 29368 9512 29420 9518
rect 29368 9454 29420 9460
rect 28908 8968 28960 8974
rect 28908 8910 28960 8916
rect 27896 8832 27948 8838
rect 27896 8774 27948 8780
rect 27988 8832 28040 8838
rect 27988 8774 28040 8780
rect 27908 8498 27936 8774
rect 28000 8498 28028 8774
rect 29380 8634 29408 9454
rect 29840 9178 29868 9522
rect 29828 9172 29880 9178
rect 29828 9114 29880 9120
rect 30024 9042 30052 10134
rect 31022 10024 31078 10033
rect 30196 9988 30248 9994
rect 31022 9959 31078 9968
rect 30196 9930 30248 9936
rect 30012 9036 30064 9042
rect 30012 8978 30064 8984
rect 29368 8628 29420 8634
rect 29368 8570 29420 8576
rect 27896 8492 27948 8498
rect 27896 8434 27948 8440
rect 27988 8492 28040 8498
rect 27988 8434 28040 8440
rect 28540 8492 28592 8498
rect 28540 8434 28592 8440
rect 27804 8424 27856 8430
rect 27804 8366 27856 8372
rect 27712 6860 27764 6866
rect 27712 6802 27764 6808
rect 27620 6452 27672 6458
rect 27620 6394 27672 6400
rect 27436 6112 27488 6118
rect 27436 6054 27488 6060
rect 22836 5704 22888 5710
rect 22836 5646 22888 5652
rect 25964 5704 26016 5710
rect 25964 5646 26016 5652
rect 27344 5704 27396 5710
rect 27344 5646 27396 5652
rect 27448 5574 27476 6054
rect 27724 5710 27752 6802
rect 27908 6730 27936 8434
rect 28552 7886 28580 8434
rect 28540 7880 28592 7886
rect 28540 7822 28592 7828
rect 28448 7744 28500 7750
rect 28448 7686 28500 7692
rect 28460 7478 28488 7686
rect 28552 7546 28580 7822
rect 28540 7540 28592 7546
rect 28540 7482 28592 7488
rect 28448 7472 28500 7478
rect 28448 7414 28500 7420
rect 30024 6866 30052 8978
rect 30208 8974 30236 9930
rect 30662 9820 30970 9829
rect 30662 9818 30668 9820
rect 30724 9818 30748 9820
rect 30804 9818 30828 9820
rect 30884 9818 30908 9820
rect 30964 9818 30970 9820
rect 30724 9766 30726 9818
rect 30906 9766 30908 9818
rect 30662 9764 30668 9766
rect 30724 9764 30748 9766
rect 30804 9764 30828 9766
rect 30884 9764 30908 9766
rect 30964 9764 30970 9766
rect 30662 9755 30970 9764
rect 31036 9722 31064 9959
rect 31024 9716 31076 9722
rect 31024 9658 31076 9664
rect 30196 8968 30248 8974
rect 30196 8910 30248 8916
rect 30662 8732 30970 8741
rect 30662 8730 30668 8732
rect 30724 8730 30748 8732
rect 30804 8730 30828 8732
rect 30884 8730 30908 8732
rect 30964 8730 30970 8732
rect 30724 8678 30726 8730
rect 30906 8678 30908 8730
rect 30662 8676 30668 8678
rect 30724 8676 30748 8678
rect 30804 8676 30828 8678
rect 30884 8676 30908 8678
rect 30964 8676 30970 8678
rect 30662 8667 30970 8676
rect 30662 7644 30970 7653
rect 30662 7642 30668 7644
rect 30724 7642 30748 7644
rect 30804 7642 30828 7644
rect 30884 7642 30908 7644
rect 30964 7642 30970 7644
rect 30724 7590 30726 7642
rect 30906 7590 30908 7642
rect 30662 7588 30668 7590
rect 30724 7588 30748 7590
rect 30804 7588 30828 7590
rect 30884 7588 30908 7590
rect 30964 7588 30970 7590
rect 30662 7579 30970 7588
rect 30012 6860 30064 6866
rect 30012 6802 30064 6808
rect 28816 6792 28868 6798
rect 28816 6734 28868 6740
rect 28908 6792 28960 6798
rect 28908 6734 28960 6740
rect 27896 6724 27948 6730
rect 27896 6666 27948 6672
rect 27908 5846 27936 6666
rect 28448 6656 28500 6662
rect 28448 6598 28500 6604
rect 28356 6452 28408 6458
rect 28356 6394 28408 6400
rect 27896 5840 27948 5846
rect 27896 5782 27948 5788
rect 27712 5704 27764 5710
rect 27712 5646 27764 5652
rect 27436 5568 27488 5574
rect 27436 5510 27488 5516
rect 23234 5468 23542 5477
rect 23234 5466 23240 5468
rect 23296 5466 23320 5468
rect 23376 5466 23400 5468
rect 23456 5466 23480 5468
rect 23536 5466 23542 5468
rect 23296 5414 23298 5466
rect 23478 5414 23480 5466
rect 23234 5412 23240 5414
rect 23296 5412 23320 5414
rect 23376 5412 23400 5414
rect 23456 5412 23480 5414
rect 23536 5412 23542 5414
rect 23234 5403 23542 5412
rect 27448 5234 27476 5510
rect 27724 5234 27752 5646
rect 27908 5642 27936 5782
rect 28368 5710 28396 6394
rect 28460 6186 28488 6598
rect 28828 6254 28856 6734
rect 28920 6390 28948 6734
rect 30662 6556 30970 6565
rect 30662 6554 30668 6556
rect 30724 6554 30748 6556
rect 30804 6554 30828 6556
rect 30884 6554 30908 6556
rect 30964 6554 30970 6556
rect 30724 6502 30726 6554
rect 30906 6502 30908 6554
rect 30662 6500 30668 6502
rect 30724 6500 30748 6502
rect 30804 6500 30828 6502
rect 30884 6500 30908 6502
rect 30964 6500 30970 6502
rect 30662 6491 30970 6500
rect 28908 6384 28960 6390
rect 28908 6326 28960 6332
rect 28816 6248 28868 6254
rect 28816 6190 28868 6196
rect 28448 6180 28500 6186
rect 28448 6122 28500 6128
rect 28356 5704 28408 5710
rect 28356 5646 28408 5652
rect 27896 5636 27948 5642
rect 27896 5578 27948 5584
rect 27908 5370 27936 5578
rect 27896 5364 27948 5370
rect 27896 5306 27948 5312
rect 28368 5302 28396 5646
rect 28356 5296 28408 5302
rect 28356 5238 28408 5244
rect 27436 5228 27488 5234
rect 27436 5170 27488 5176
rect 27712 5228 27764 5234
rect 27712 5170 27764 5176
rect 28460 5098 28488 6122
rect 28724 5772 28776 5778
rect 28724 5714 28776 5720
rect 28736 5234 28764 5714
rect 28828 5234 28856 6190
rect 28920 5914 28948 6326
rect 29092 6316 29144 6322
rect 29092 6258 29144 6264
rect 29104 5914 29132 6258
rect 29828 6112 29880 6118
rect 29828 6054 29880 6060
rect 31022 6080 31078 6089
rect 28908 5908 28960 5914
rect 28908 5850 28960 5856
rect 29092 5908 29144 5914
rect 29092 5850 29144 5856
rect 29840 5710 29868 6054
rect 31022 6015 31078 6024
rect 31036 5778 31064 6015
rect 31024 5772 31076 5778
rect 31024 5714 31076 5720
rect 29828 5704 29880 5710
rect 29828 5646 29880 5652
rect 30662 5468 30970 5477
rect 30662 5466 30668 5468
rect 30724 5466 30748 5468
rect 30804 5466 30828 5468
rect 30884 5466 30908 5468
rect 30964 5466 30970 5468
rect 30724 5414 30726 5466
rect 30906 5414 30908 5466
rect 30662 5412 30668 5414
rect 30724 5412 30748 5414
rect 30804 5412 30828 5414
rect 30884 5412 30908 5414
rect 30964 5412 30970 5414
rect 30662 5403 30970 5412
rect 28724 5228 28776 5234
rect 28724 5170 28776 5176
rect 28816 5228 28868 5234
rect 28816 5170 28868 5176
rect 28448 5092 28500 5098
rect 28448 5034 28500 5040
rect 28724 5024 28776 5030
rect 28724 4966 28776 4972
rect 26948 4924 27256 4933
rect 26948 4922 26954 4924
rect 27010 4922 27034 4924
rect 27090 4922 27114 4924
rect 27170 4922 27194 4924
rect 27250 4922 27256 4924
rect 27010 4870 27012 4922
rect 27192 4870 27194 4922
rect 26948 4868 26954 4870
rect 27010 4868 27034 4870
rect 27090 4868 27114 4870
rect 27170 4868 27194 4870
rect 27250 4868 27256 4870
rect 26948 4859 27256 4868
rect 20812 4684 20864 4690
rect 20812 4626 20864 4632
rect 17960 4616 18012 4622
rect 17960 4558 18012 4564
rect 19984 4616 20036 4622
rect 19984 4558 20036 4564
rect 15806 4380 16114 4389
rect 15806 4378 15812 4380
rect 15868 4378 15892 4380
rect 15948 4378 15972 4380
rect 16028 4378 16052 4380
rect 16108 4378 16114 4380
rect 15868 4326 15870 4378
rect 16050 4326 16052 4378
rect 15806 4324 15812 4326
rect 15868 4324 15892 4326
rect 15948 4324 15972 4326
rect 16028 4324 16052 4326
rect 16108 4324 16114 4326
rect 15806 4315 16114 4324
rect 23234 4380 23542 4389
rect 23234 4378 23240 4380
rect 23296 4378 23320 4380
rect 23376 4378 23400 4380
rect 23456 4378 23480 4380
rect 23536 4378 23542 4380
rect 23296 4326 23298 4378
rect 23478 4326 23480 4378
rect 23234 4324 23240 4326
rect 23296 4324 23320 4326
rect 23376 4324 23400 4326
rect 23456 4324 23480 4326
rect 23536 4324 23542 4326
rect 23234 4315 23542 4324
rect 14648 4276 14700 4282
rect 14648 4218 14700 4224
rect 14372 4208 14424 4214
rect 14372 4150 14424 4156
rect 14004 4140 14056 4146
rect 14004 4082 14056 4088
rect 4664 3836 4972 3845
rect 4664 3834 4670 3836
rect 4726 3834 4750 3836
rect 4806 3834 4830 3836
rect 4886 3834 4910 3836
rect 4966 3834 4972 3836
rect 4726 3782 4728 3834
rect 4908 3782 4910 3834
rect 4664 3780 4670 3782
rect 4726 3780 4750 3782
rect 4806 3780 4830 3782
rect 4886 3780 4910 3782
rect 4966 3780 4972 3782
rect 4664 3771 4972 3780
rect 12092 3836 12400 3845
rect 12092 3834 12098 3836
rect 12154 3834 12178 3836
rect 12234 3834 12258 3836
rect 12314 3834 12338 3836
rect 12394 3834 12400 3836
rect 12154 3782 12156 3834
rect 12336 3782 12338 3834
rect 12092 3780 12098 3782
rect 12154 3780 12178 3782
rect 12234 3780 12258 3782
rect 12314 3780 12338 3782
rect 12394 3780 12400 3782
rect 12092 3771 12400 3780
rect 19520 3836 19828 3845
rect 19520 3834 19526 3836
rect 19582 3834 19606 3836
rect 19662 3834 19686 3836
rect 19742 3834 19766 3836
rect 19822 3834 19828 3836
rect 19582 3782 19584 3834
rect 19764 3782 19766 3834
rect 19520 3780 19526 3782
rect 19582 3780 19606 3782
rect 19662 3780 19686 3782
rect 19742 3780 19766 3782
rect 19822 3780 19828 3782
rect 19520 3771 19828 3780
rect 26948 3836 27256 3845
rect 26948 3834 26954 3836
rect 27010 3834 27034 3836
rect 27090 3834 27114 3836
rect 27170 3834 27194 3836
rect 27250 3834 27256 3836
rect 27010 3782 27012 3834
rect 27192 3782 27194 3834
rect 26948 3780 26954 3782
rect 27010 3780 27034 3782
rect 27090 3780 27114 3782
rect 27170 3780 27194 3782
rect 27250 3780 27256 3782
rect 26948 3771 27256 3780
rect 8378 3292 8686 3301
rect 8378 3290 8384 3292
rect 8440 3290 8464 3292
rect 8520 3290 8544 3292
rect 8600 3290 8624 3292
rect 8680 3290 8686 3292
rect 8440 3238 8442 3290
rect 8622 3238 8624 3290
rect 8378 3236 8384 3238
rect 8440 3236 8464 3238
rect 8520 3236 8544 3238
rect 8600 3236 8624 3238
rect 8680 3236 8686 3238
rect 8378 3227 8686 3236
rect 15806 3292 16114 3301
rect 15806 3290 15812 3292
rect 15868 3290 15892 3292
rect 15948 3290 15972 3292
rect 16028 3290 16052 3292
rect 16108 3290 16114 3292
rect 15868 3238 15870 3290
rect 16050 3238 16052 3290
rect 15806 3236 15812 3238
rect 15868 3236 15892 3238
rect 15948 3236 15972 3238
rect 16028 3236 16052 3238
rect 16108 3236 16114 3238
rect 15806 3227 16114 3236
rect 23234 3292 23542 3301
rect 23234 3290 23240 3292
rect 23296 3290 23320 3292
rect 23376 3290 23400 3292
rect 23456 3290 23480 3292
rect 23536 3290 23542 3292
rect 23296 3238 23298 3290
rect 23478 3238 23480 3290
rect 23234 3236 23240 3238
rect 23296 3236 23320 3238
rect 23376 3236 23400 3238
rect 23456 3236 23480 3238
rect 23536 3236 23542 3238
rect 23234 3227 23542 3236
rect 4664 2748 4972 2757
rect 4664 2746 4670 2748
rect 4726 2746 4750 2748
rect 4806 2746 4830 2748
rect 4886 2746 4910 2748
rect 4966 2746 4972 2748
rect 4726 2694 4728 2746
rect 4908 2694 4910 2746
rect 4664 2692 4670 2694
rect 4726 2692 4750 2694
rect 4806 2692 4830 2694
rect 4886 2692 4910 2694
rect 4966 2692 4972 2694
rect 4664 2683 4972 2692
rect 12092 2748 12400 2757
rect 12092 2746 12098 2748
rect 12154 2746 12178 2748
rect 12234 2746 12258 2748
rect 12314 2746 12338 2748
rect 12394 2746 12400 2748
rect 12154 2694 12156 2746
rect 12336 2694 12338 2746
rect 12092 2692 12098 2694
rect 12154 2692 12178 2694
rect 12234 2692 12258 2694
rect 12314 2692 12338 2694
rect 12394 2692 12400 2694
rect 12092 2683 12400 2692
rect 19520 2748 19828 2757
rect 19520 2746 19526 2748
rect 19582 2746 19606 2748
rect 19662 2746 19686 2748
rect 19742 2746 19766 2748
rect 19822 2746 19828 2748
rect 19582 2694 19584 2746
rect 19764 2694 19766 2746
rect 19520 2692 19526 2694
rect 19582 2692 19606 2694
rect 19662 2692 19686 2694
rect 19742 2692 19766 2694
rect 19822 2692 19828 2694
rect 19520 2683 19828 2692
rect 26948 2748 27256 2757
rect 26948 2746 26954 2748
rect 27010 2746 27034 2748
rect 27090 2746 27114 2748
rect 27170 2746 27194 2748
rect 27250 2746 27256 2748
rect 27010 2694 27012 2746
rect 27192 2694 27194 2746
rect 26948 2692 26954 2694
rect 27010 2692 27034 2694
rect 27090 2692 27114 2694
rect 27170 2692 27194 2694
rect 27250 2692 27256 2694
rect 26948 2683 27256 2692
rect 28736 2446 28764 4966
rect 30662 4380 30970 4389
rect 30662 4378 30668 4380
rect 30724 4378 30748 4380
rect 30804 4378 30828 4380
rect 30884 4378 30908 4380
rect 30964 4378 30970 4380
rect 30724 4326 30726 4378
rect 30906 4326 30908 4378
rect 30662 4324 30668 4326
rect 30724 4324 30748 4326
rect 30804 4324 30828 4326
rect 30884 4324 30908 4326
rect 30964 4324 30970 4326
rect 30662 4315 30970 4324
rect 30662 3292 30970 3301
rect 30662 3290 30668 3292
rect 30724 3290 30748 3292
rect 30804 3290 30828 3292
rect 30884 3290 30908 3292
rect 30964 3290 30970 3292
rect 30724 3238 30726 3290
rect 30906 3238 30908 3290
rect 30662 3236 30668 3238
rect 30724 3236 30748 3238
rect 30804 3236 30828 3238
rect 30884 3236 30908 3238
rect 30964 3236 30970 3238
rect 30662 3227 30970 3236
rect 28724 2440 28776 2446
rect 28724 2382 28776 2388
rect 31024 2372 31076 2378
rect 31024 2314 31076 2320
rect 8378 2204 8686 2213
rect 8378 2202 8384 2204
rect 8440 2202 8464 2204
rect 8520 2202 8544 2204
rect 8600 2202 8624 2204
rect 8680 2202 8686 2204
rect 8440 2150 8442 2202
rect 8622 2150 8624 2202
rect 8378 2148 8384 2150
rect 8440 2148 8464 2150
rect 8520 2148 8544 2150
rect 8600 2148 8624 2150
rect 8680 2148 8686 2150
rect 8378 2139 8686 2148
rect 15806 2204 16114 2213
rect 15806 2202 15812 2204
rect 15868 2202 15892 2204
rect 15948 2202 15972 2204
rect 16028 2202 16052 2204
rect 16108 2202 16114 2204
rect 15868 2150 15870 2202
rect 16050 2150 16052 2202
rect 15806 2148 15812 2150
rect 15868 2148 15892 2150
rect 15948 2148 15972 2150
rect 16028 2148 16052 2150
rect 16108 2148 16114 2150
rect 15806 2139 16114 2148
rect 23234 2204 23542 2213
rect 23234 2202 23240 2204
rect 23296 2202 23320 2204
rect 23376 2202 23400 2204
rect 23456 2202 23480 2204
rect 23536 2202 23542 2204
rect 23296 2150 23298 2202
rect 23478 2150 23480 2202
rect 23234 2148 23240 2150
rect 23296 2148 23320 2150
rect 23376 2148 23400 2150
rect 23456 2148 23480 2150
rect 23536 2148 23542 2150
rect 23234 2139 23542 2148
rect 30662 2204 30970 2213
rect 30662 2202 30668 2204
rect 30724 2202 30748 2204
rect 30804 2202 30828 2204
rect 30884 2202 30908 2204
rect 30964 2202 30970 2204
rect 30724 2150 30726 2202
rect 30906 2150 30908 2202
rect 30662 2148 30668 2150
rect 30724 2148 30748 2150
rect 30804 2148 30828 2150
rect 30884 2148 30908 2150
rect 30964 2148 30970 2150
rect 30662 2139 30970 2148
rect 31036 2009 31064 2314
rect 31022 2000 31078 2009
rect 31022 1935 31078 1944
<< via2 >>
rect 8384 29402 8440 29404
rect 8464 29402 8520 29404
rect 8544 29402 8600 29404
rect 8624 29402 8680 29404
rect 8384 29350 8430 29402
rect 8430 29350 8440 29402
rect 8464 29350 8494 29402
rect 8494 29350 8506 29402
rect 8506 29350 8520 29402
rect 8544 29350 8558 29402
rect 8558 29350 8570 29402
rect 8570 29350 8600 29402
rect 8624 29350 8634 29402
rect 8634 29350 8680 29402
rect 8384 29348 8440 29350
rect 8464 29348 8520 29350
rect 8544 29348 8600 29350
rect 8624 29348 8680 29350
rect 15812 29402 15868 29404
rect 15892 29402 15948 29404
rect 15972 29402 16028 29404
rect 16052 29402 16108 29404
rect 15812 29350 15858 29402
rect 15858 29350 15868 29402
rect 15892 29350 15922 29402
rect 15922 29350 15934 29402
rect 15934 29350 15948 29402
rect 15972 29350 15986 29402
rect 15986 29350 15998 29402
rect 15998 29350 16028 29402
rect 16052 29350 16062 29402
rect 16062 29350 16108 29402
rect 15812 29348 15868 29350
rect 15892 29348 15948 29350
rect 15972 29348 16028 29350
rect 16052 29348 16108 29350
rect 4670 28858 4726 28860
rect 4750 28858 4806 28860
rect 4830 28858 4886 28860
rect 4910 28858 4966 28860
rect 4670 28806 4716 28858
rect 4716 28806 4726 28858
rect 4750 28806 4780 28858
rect 4780 28806 4792 28858
rect 4792 28806 4806 28858
rect 4830 28806 4844 28858
rect 4844 28806 4856 28858
rect 4856 28806 4886 28858
rect 4910 28806 4920 28858
rect 4920 28806 4966 28858
rect 4670 28804 4726 28806
rect 4750 28804 4806 28806
rect 4830 28804 4886 28806
rect 4910 28804 4966 28806
rect 12098 28858 12154 28860
rect 12178 28858 12234 28860
rect 12258 28858 12314 28860
rect 12338 28858 12394 28860
rect 12098 28806 12144 28858
rect 12144 28806 12154 28858
rect 12178 28806 12208 28858
rect 12208 28806 12220 28858
rect 12220 28806 12234 28858
rect 12258 28806 12272 28858
rect 12272 28806 12284 28858
rect 12284 28806 12314 28858
rect 12338 28806 12348 28858
rect 12348 28806 12394 28858
rect 12098 28804 12154 28806
rect 12178 28804 12234 28806
rect 12258 28804 12314 28806
rect 12338 28804 12394 28806
rect 4670 27770 4726 27772
rect 4750 27770 4806 27772
rect 4830 27770 4886 27772
rect 4910 27770 4966 27772
rect 4670 27718 4716 27770
rect 4716 27718 4726 27770
rect 4750 27718 4780 27770
rect 4780 27718 4792 27770
rect 4792 27718 4806 27770
rect 4830 27718 4844 27770
rect 4844 27718 4856 27770
rect 4856 27718 4886 27770
rect 4910 27718 4920 27770
rect 4920 27718 4966 27770
rect 4670 27716 4726 27718
rect 4750 27716 4806 27718
rect 4830 27716 4886 27718
rect 4910 27716 4966 27718
rect 4670 26682 4726 26684
rect 4750 26682 4806 26684
rect 4830 26682 4886 26684
rect 4910 26682 4966 26684
rect 4670 26630 4716 26682
rect 4716 26630 4726 26682
rect 4750 26630 4780 26682
rect 4780 26630 4792 26682
rect 4792 26630 4806 26682
rect 4830 26630 4844 26682
rect 4844 26630 4856 26682
rect 4856 26630 4886 26682
rect 4910 26630 4920 26682
rect 4920 26630 4966 26682
rect 4670 26628 4726 26630
rect 4750 26628 4806 26630
rect 4830 26628 4886 26630
rect 4910 26628 4966 26630
rect 4670 25594 4726 25596
rect 4750 25594 4806 25596
rect 4830 25594 4886 25596
rect 4910 25594 4966 25596
rect 4670 25542 4716 25594
rect 4716 25542 4726 25594
rect 4750 25542 4780 25594
rect 4780 25542 4792 25594
rect 4792 25542 4806 25594
rect 4830 25542 4844 25594
rect 4844 25542 4856 25594
rect 4856 25542 4886 25594
rect 4910 25542 4920 25594
rect 4920 25542 4966 25594
rect 4670 25540 4726 25542
rect 4750 25540 4806 25542
rect 4830 25540 4886 25542
rect 4910 25540 4966 25542
rect 4670 24506 4726 24508
rect 4750 24506 4806 24508
rect 4830 24506 4886 24508
rect 4910 24506 4966 24508
rect 4670 24454 4716 24506
rect 4716 24454 4726 24506
rect 4750 24454 4780 24506
rect 4780 24454 4792 24506
rect 4792 24454 4806 24506
rect 4830 24454 4844 24506
rect 4844 24454 4856 24506
rect 4856 24454 4886 24506
rect 4910 24454 4920 24506
rect 4920 24454 4966 24506
rect 4670 24452 4726 24454
rect 4750 24452 4806 24454
rect 4830 24452 4886 24454
rect 4910 24452 4966 24454
rect 4670 23418 4726 23420
rect 4750 23418 4806 23420
rect 4830 23418 4886 23420
rect 4910 23418 4966 23420
rect 4670 23366 4716 23418
rect 4716 23366 4726 23418
rect 4750 23366 4780 23418
rect 4780 23366 4792 23418
rect 4792 23366 4806 23418
rect 4830 23366 4844 23418
rect 4844 23366 4856 23418
rect 4856 23366 4886 23418
rect 4910 23366 4920 23418
rect 4920 23366 4966 23418
rect 4670 23364 4726 23366
rect 4750 23364 4806 23366
rect 4830 23364 4886 23366
rect 4910 23364 4966 23366
rect 4670 22330 4726 22332
rect 4750 22330 4806 22332
rect 4830 22330 4886 22332
rect 4910 22330 4966 22332
rect 4670 22278 4716 22330
rect 4716 22278 4726 22330
rect 4750 22278 4780 22330
rect 4780 22278 4792 22330
rect 4792 22278 4806 22330
rect 4830 22278 4844 22330
rect 4844 22278 4856 22330
rect 4856 22278 4886 22330
rect 4910 22278 4920 22330
rect 4920 22278 4966 22330
rect 4670 22276 4726 22278
rect 4750 22276 4806 22278
rect 4830 22276 4886 22278
rect 4910 22276 4966 22278
rect 4670 21242 4726 21244
rect 4750 21242 4806 21244
rect 4830 21242 4886 21244
rect 4910 21242 4966 21244
rect 4670 21190 4716 21242
rect 4716 21190 4726 21242
rect 4750 21190 4780 21242
rect 4780 21190 4792 21242
rect 4792 21190 4806 21242
rect 4830 21190 4844 21242
rect 4844 21190 4856 21242
rect 4856 21190 4886 21242
rect 4910 21190 4920 21242
rect 4920 21190 4966 21242
rect 4670 21188 4726 21190
rect 4750 21188 4806 21190
rect 4830 21188 4886 21190
rect 4910 21188 4966 21190
rect 4670 20154 4726 20156
rect 4750 20154 4806 20156
rect 4830 20154 4886 20156
rect 4910 20154 4966 20156
rect 4670 20102 4716 20154
rect 4716 20102 4726 20154
rect 4750 20102 4780 20154
rect 4780 20102 4792 20154
rect 4792 20102 4806 20154
rect 4830 20102 4844 20154
rect 4844 20102 4856 20154
rect 4856 20102 4886 20154
rect 4910 20102 4920 20154
rect 4920 20102 4966 20154
rect 4670 20100 4726 20102
rect 4750 20100 4806 20102
rect 4830 20100 4886 20102
rect 4910 20100 4966 20102
rect 4670 19066 4726 19068
rect 4750 19066 4806 19068
rect 4830 19066 4886 19068
rect 4910 19066 4966 19068
rect 4670 19014 4716 19066
rect 4716 19014 4726 19066
rect 4750 19014 4780 19066
rect 4780 19014 4792 19066
rect 4792 19014 4806 19066
rect 4830 19014 4844 19066
rect 4844 19014 4856 19066
rect 4856 19014 4886 19066
rect 4910 19014 4920 19066
rect 4920 19014 4966 19066
rect 4670 19012 4726 19014
rect 4750 19012 4806 19014
rect 4830 19012 4886 19014
rect 4910 19012 4966 19014
rect 4670 17978 4726 17980
rect 4750 17978 4806 17980
rect 4830 17978 4886 17980
rect 4910 17978 4966 17980
rect 4670 17926 4716 17978
rect 4716 17926 4726 17978
rect 4750 17926 4780 17978
rect 4780 17926 4792 17978
rect 4792 17926 4806 17978
rect 4830 17926 4844 17978
rect 4844 17926 4856 17978
rect 4856 17926 4886 17978
rect 4910 17926 4920 17978
rect 4920 17926 4966 17978
rect 4670 17924 4726 17926
rect 4750 17924 4806 17926
rect 4830 17924 4886 17926
rect 4910 17924 4966 17926
rect 8384 28314 8440 28316
rect 8464 28314 8520 28316
rect 8544 28314 8600 28316
rect 8624 28314 8680 28316
rect 8384 28262 8430 28314
rect 8430 28262 8440 28314
rect 8464 28262 8494 28314
rect 8494 28262 8506 28314
rect 8506 28262 8520 28314
rect 8544 28262 8558 28314
rect 8558 28262 8570 28314
rect 8570 28262 8600 28314
rect 8624 28262 8634 28314
rect 8634 28262 8680 28314
rect 8384 28260 8440 28262
rect 8464 28260 8520 28262
rect 8544 28260 8600 28262
rect 8624 28260 8680 28262
rect 8384 27226 8440 27228
rect 8464 27226 8520 27228
rect 8544 27226 8600 27228
rect 8624 27226 8680 27228
rect 8384 27174 8430 27226
rect 8430 27174 8440 27226
rect 8464 27174 8494 27226
rect 8494 27174 8506 27226
rect 8506 27174 8520 27226
rect 8544 27174 8558 27226
rect 8558 27174 8570 27226
rect 8570 27174 8600 27226
rect 8624 27174 8634 27226
rect 8634 27174 8680 27226
rect 8384 27172 8440 27174
rect 8464 27172 8520 27174
rect 8544 27172 8600 27174
rect 8624 27172 8680 27174
rect 12098 27770 12154 27772
rect 12178 27770 12234 27772
rect 12258 27770 12314 27772
rect 12338 27770 12394 27772
rect 12098 27718 12144 27770
rect 12144 27718 12154 27770
rect 12178 27718 12208 27770
rect 12208 27718 12220 27770
rect 12220 27718 12234 27770
rect 12258 27718 12272 27770
rect 12272 27718 12284 27770
rect 12284 27718 12314 27770
rect 12338 27718 12348 27770
rect 12348 27718 12394 27770
rect 12098 27716 12154 27718
rect 12178 27716 12234 27718
rect 12258 27716 12314 27718
rect 12338 27716 12394 27718
rect 12098 26682 12154 26684
rect 12178 26682 12234 26684
rect 12258 26682 12314 26684
rect 12338 26682 12394 26684
rect 12098 26630 12144 26682
rect 12144 26630 12154 26682
rect 12178 26630 12208 26682
rect 12208 26630 12220 26682
rect 12220 26630 12234 26682
rect 12258 26630 12272 26682
rect 12272 26630 12284 26682
rect 12284 26630 12314 26682
rect 12338 26630 12348 26682
rect 12348 26630 12394 26682
rect 12098 26628 12154 26630
rect 12178 26628 12234 26630
rect 12258 26628 12314 26630
rect 12338 26628 12394 26630
rect 8384 26138 8440 26140
rect 8464 26138 8520 26140
rect 8544 26138 8600 26140
rect 8624 26138 8680 26140
rect 8384 26086 8430 26138
rect 8430 26086 8440 26138
rect 8464 26086 8494 26138
rect 8494 26086 8506 26138
rect 8506 26086 8520 26138
rect 8544 26086 8558 26138
rect 8558 26086 8570 26138
rect 8570 26086 8600 26138
rect 8624 26086 8634 26138
rect 8634 26086 8680 26138
rect 8384 26084 8440 26086
rect 8464 26084 8520 26086
rect 8544 26084 8600 26086
rect 8624 26084 8680 26086
rect 8384 25050 8440 25052
rect 8464 25050 8520 25052
rect 8544 25050 8600 25052
rect 8624 25050 8680 25052
rect 8384 24998 8430 25050
rect 8430 24998 8440 25050
rect 8464 24998 8494 25050
rect 8494 24998 8506 25050
rect 8506 24998 8520 25050
rect 8544 24998 8558 25050
rect 8558 24998 8570 25050
rect 8570 24998 8600 25050
rect 8624 24998 8634 25050
rect 8634 24998 8680 25050
rect 8384 24996 8440 24998
rect 8464 24996 8520 24998
rect 8544 24996 8600 24998
rect 8624 24996 8680 24998
rect 8384 23962 8440 23964
rect 8464 23962 8520 23964
rect 8544 23962 8600 23964
rect 8624 23962 8680 23964
rect 8384 23910 8430 23962
rect 8430 23910 8440 23962
rect 8464 23910 8494 23962
rect 8494 23910 8506 23962
rect 8506 23910 8520 23962
rect 8544 23910 8558 23962
rect 8558 23910 8570 23962
rect 8570 23910 8600 23962
rect 8624 23910 8634 23962
rect 8634 23910 8680 23962
rect 8384 23908 8440 23910
rect 8464 23908 8520 23910
rect 8544 23908 8600 23910
rect 8624 23908 8680 23910
rect 8384 22874 8440 22876
rect 8464 22874 8520 22876
rect 8544 22874 8600 22876
rect 8624 22874 8680 22876
rect 8384 22822 8430 22874
rect 8430 22822 8440 22874
rect 8464 22822 8494 22874
rect 8494 22822 8506 22874
rect 8506 22822 8520 22874
rect 8544 22822 8558 22874
rect 8558 22822 8570 22874
rect 8570 22822 8600 22874
rect 8624 22822 8634 22874
rect 8634 22822 8680 22874
rect 8384 22820 8440 22822
rect 8464 22820 8520 22822
rect 8544 22820 8600 22822
rect 8624 22820 8680 22822
rect 8384 21786 8440 21788
rect 8464 21786 8520 21788
rect 8544 21786 8600 21788
rect 8624 21786 8680 21788
rect 8384 21734 8430 21786
rect 8430 21734 8440 21786
rect 8464 21734 8494 21786
rect 8494 21734 8506 21786
rect 8506 21734 8520 21786
rect 8544 21734 8558 21786
rect 8558 21734 8570 21786
rect 8570 21734 8600 21786
rect 8624 21734 8634 21786
rect 8634 21734 8680 21786
rect 8384 21732 8440 21734
rect 8464 21732 8520 21734
rect 8544 21732 8600 21734
rect 8624 21732 8680 21734
rect 4670 16890 4726 16892
rect 4750 16890 4806 16892
rect 4830 16890 4886 16892
rect 4910 16890 4966 16892
rect 4670 16838 4716 16890
rect 4716 16838 4726 16890
rect 4750 16838 4780 16890
rect 4780 16838 4792 16890
rect 4792 16838 4806 16890
rect 4830 16838 4844 16890
rect 4844 16838 4856 16890
rect 4856 16838 4886 16890
rect 4910 16838 4920 16890
rect 4920 16838 4966 16890
rect 4670 16836 4726 16838
rect 4750 16836 4806 16838
rect 4830 16836 4886 16838
rect 4910 16836 4966 16838
rect 4670 15802 4726 15804
rect 4750 15802 4806 15804
rect 4830 15802 4886 15804
rect 4910 15802 4966 15804
rect 4670 15750 4716 15802
rect 4716 15750 4726 15802
rect 4750 15750 4780 15802
rect 4780 15750 4792 15802
rect 4792 15750 4806 15802
rect 4830 15750 4844 15802
rect 4844 15750 4856 15802
rect 4856 15750 4886 15802
rect 4910 15750 4920 15802
rect 4920 15750 4966 15802
rect 4670 15748 4726 15750
rect 4750 15748 4806 15750
rect 4830 15748 4886 15750
rect 4910 15748 4966 15750
rect 4670 14714 4726 14716
rect 4750 14714 4806 14716
rect 4830 14714 4886 14716
rect 4910 14714 4966 14716
rect 4670 14662 4716 14714
rect 4716 14662 4726 14714
rect 4750 14662 4780 14714
rect 4780 14662 4792 14714
rect 4792 14662 4806 14714
rect 4830 14662 4844 14714
rect 4844 14662 4856 14714
rect 4856 14662 4886 14714
rect 4910 14662 4920 14714
rect 4920 14662 4966 14714
rect 4670 14660 4726 14662
rect 4750 14660 4806 14662
rect 4830 14660 4886 14662
rect 4910 14660 4966 14662
rect 4670 13626 4726 13628
rect 4750 13626 4806 13628
rect 4830 13626 4886 13628
rect 4910 13626 4966 13628
rect 4670 13574 4716 13626
rect 4716 13574 4726 13626
rect 4750 13574 4780 13626
rect 4780 13574 4792 13626
rect 4792 13574 4806 13626
rect 4830 13574 4844 13626
rect 4844 13574 4856 13626
rect 4856 13574 4886 13626
rect 4910 13574 4920 13626
rect 4920 13574 4966 13626
rect 4670 13572 4726 13574
rect 4750 13572 4806 13574
rect 4830 13572 4886 13574
rect 4910 13572 4966 13574
rect 4670 12538 4726 12540
rect 4750 12538 4806 12540
rect 4830 12538 4886 12540
rect 4910 12538 4966 12540
rect 4670 12486 4716 12538
rect 4716 12486 4726 12538
rect 4750 12486 4780 12538
rect 4780 12486 4792 12538
rect 4792 12486 4806 12538
rect 4830 12486 4844 12538
rect 4844 12486 4856 12538
rect 4856 12486 4886 12538
rect 4910 12486 4920 12538
rect 4920 12486 4966 12538
rect 4670 12484 4726 12486
rect 4750 12484 4806 12486
rect 4830 12484 4886 12486
rect 4910 12484 4966 12486
rect 4670 11450 4726 11452
rect 4750 11450 4806 11452
rect 4830 11450 4886 11452
rect 4910 11450 4966 11452
rect 4670 11398 4716 11450
rect 4716 11398 4726 11450
rect 4750 11398 4780 11450
rect 4780 11398 4792 11450
rect 4792 11398 4806 11450
rect 4830 11398 4844 11450
rect 4844 11398 4856 11450
rect 4856 11398 4886 11450
rect 4910 11398 4920 11450
rect 4920 11398 4966 11450
rect 4670 11396 4726 11398
rect 4750 11396 4806 11398
rect 4830 11396 4886 11398
rect 4910 11396 4966 11398
rect 4670 10362 4726 10364
rect 4750 10362 4806 10364
rect 4830 10362 4886 10364
rect 4910 10362 4966 10364
rect 4670 10310 4716 10362
rect 4716 10310 4726 10362
rect 4750 10310 4780 10362
rect 4780 10310 4792 10362
rect 4792 10310 4806 10362
rect 4830 10310 4844 10362
rect 4844 10310 4856 10362
rect 4856 10310 4886 10362
rect 4910 10310 4920 10362
rect 4920 10310 4966 10362
rect 4670 10308 4726 10310
rect 4750 10308 4806 10310
rect 4830 10308 4886 10310
rect 4910 10308 4966 10310
rect 4670 9274 4726 9276
rect 4750 9274 4806 9276
rect 4830 9274 4886 9276
rect 4910 9274 4966 9276
rect 4670 9222 4716 9274
rect 4716 9222 4726 9274
rect 4750 9222 4780 9274
rect 4780 9222 4792 9274
rect 4792 9222 4806 9274
rect 4830 9222 4844 9274
rect 4844 9222 4856 9274
rect 4856 9222 4886 9274
rect 4910 9222 4920 9274
rect 4920 9222 4966 9274
rect 4670 9220 4726 9222
rect 4750 9220 4806 9222
rect 4830 9220 4886 9222
rect 4910 9220 4966 9222
rect 4670 8186 4726 8188
rect 4750 8186 4806 8188
rect 4830 8186 4886 8188
rect 4910 8186 4966 8188
rect 4670 8134 4716 8186
rect 4716 8134 4726 8186
rect 4750 8134 4780 8186
rect 4780 8134 4792 8186
rect 4792 8134 4806 8186
rect 4830 8134 4844 8186
rect 4844 8134 4856 8186
rect 4856 8134 4886 8186
rect 4910 8134 4920 8186
rect 4920 8134 4966 8186
rect 4670 8132 4726 8134
rect 4750 8132 4806 8134
rect 4830 8132 4886 8134
rect 4910 8132 4966 8134
rect 4670 7098 4726 7100
rect 4750 7098 4806 7100
rect 4830 7098 4886 7100
rect 4910 7098 4966 7100
rect 4670 7046 4716 7098
rect 4716 7046 4726 7098
rect 4750 7046 4780 7098
rect 4780 7046 4792 7098
rect 4792 7046 4806 7098
rect 4830 7046 4844 7098
rect 4844 7046 4856 7098
rect 4856 7046 4886 7098
rect 4910 7046 4920 7098
rect 4920 7046 4966 7098
rect 4670 7044 4726 7046
rect 4750 7044 4806 7046
rect 4830 7044 4886 7046
rect 4910 7044 4966 7046
rect 8384 20698 8440 20700
rect 8464 20698 8520 20700
rect 8544 20698 8600 20700
rect 8624 20698 8680 20700
rect 8384 20646 8430 20698
rect 8430 20646 8440 20698
rect 8464 20646 8494 20698
rect 8494 20646 8506 20698
rect 8506 20646 8520 20698
rect 8544 20646 8558 20698
rect 8558 20646 8570 20698
rect 8570 20646 8600 20698
rect 8624 20646 8634 20698
rect 8634 20646 8680 20698
rect 8384 20644 8440 20646
rect 8464 20644 8520 20646
rect 8544 20644 8600 20646
rect 8624 20644 8680 20646
rect 8384 19610 8440 19612
rect 8464 19610 8520 19612
rect 8544 19610 8600 19612
rect 8624 19610 8680 19612
rect 8384 19558 8430 19610
rect 8430 19558 8440 19610
rect 8464 19558 8494 19610
rect 8494 19558 8506 19610
rect 8506 19558 8520 19610
rect 8544 19558 8558 19610
rect 8558 19558 8570 19610
rect 8570 19558 8600 19610
rect 8624 19558 8634 19610
rect 8634 19558 8680 19610
rect 8384 19556 8440 19558
rect 8464 19556 8520 19558
rect 8544 19556 8600 19558
rect 8624 19556 8680 19558
rect 8384 18522 8440 18524
rect 8464 18522 8520 18524
rect 8544 18522 8600 18524
rect 8624 18522 8680 18524
rect 8384 18470 8430 18522
rect 8430 18470 8440 18522
rect 8464 18470 8494 18522
rect 8494 18470 8506 18522
rect 8506 18470 8520 18522
rect 8544 18470 8558 18522
rect 8558 18470 8570 18522
rect 8570 18470 8600 18522
rect 8624 18470 8634 18522
rect 8634 18470 8680 18522
rect 8384 18468 8440 18470
rect 8464 18468 8520 18470
rect 8544 18468 8600 18470
rect 8624 18468 8680 18470
rect 8384 17434 8440 17436
rect 8464 17434 8520 17436
rect 8544 17434 8600 17436
rect 8624 17434 8680 17436
rect 8384 17382 8430 17434
rect 8430 17382 8440 17434
rect 8464 17382 8494 17434
rect 8494 17382 8506 17434
rect 8506 17382 8520 17434
rect 8544 17382 8558 17434
rect 8558 17382 8570 17434
rect 8570 17382 8600 17434
rect 8624 17382 8634 17434
rect 8634 17382 8680 17434
rect 8384 17380 8440 17382
rect 8464 17380 8520 17382
rect 8544 17380 8600 17382
rect 8624 17380 8680 17382
rect 8384 16346 8440 16348
rect 8464 16346 8520 16348
rect 8544 16346 8600 16348
rect 8624 16346 8680 16348
rect 8384 16294 8430 16346
rect 8430 16294 8440 16346
rect 8464 16294 8494 16346
rect 8494 16294 8506 16346
rect 8506 16294 8520 16346
rect 8544 16294 8558 16346
rect 8558 16294 8570 16346
rect 8570 16294 8600 16346
rect 8624 16294 8634 16346
rect 8634 16294 8680 16346
rect 8384 16292 8440 16294
rect 8464 16292 8520 16294
rect 8544 16292 8600 16294
rect 8624 16292 8680 16294
rect 12098 25594 12154 25596
rect 12178 25594 12234 25596
rect 12258 25594 12314 25596
rect 12338 25594 12394 25596
rect 12098 25542 12144 25594
rect 12144 25542 12154 25594
rect 12178 25542 12208 25594
rect 12208 25542 12220 25594
rect 12220 25542 12234 25594
rect 12258 25542 12272 25594
rect 12272 25542 12284 25594
rect 12284 25542 12314 25594
rect 12338 25542 12348 25594
rect 12348 25542 12394 25594
rect 12098 25540 12154 25542
rect 12178 25540 12234 25542
rect 12258 25540 12314 25542
rect 12338 25540 12394 25542
rect 12098 24506 12154 24508
rect 12178 24506 12234 24508
rect 12258 24506 12314 24508
rect 12338 24506 12394 24508
rect 12098 24454 12144 24506
rect 12144 24454 12154 24506
rect 12178 24454 12208 24506
rect 12208 24454 12220 24506
rect 12220 24454 12234 24506
rect 12258 24454 12272 24506
rect 12272 24454 12284 24506
rect 12284 24454 12314 24506
rect 12338 24454 12348 24506
rect 12348 24454 12394 24506
rect 12098 24452 12154 24454
rect 12178 24452 12234 24454
rect 12258 24452 12314 24454
rect 12338 24452 12394 24454
rect 12098 23418 12154 23420
rect 12178 23418 12234 23420
rect 12258 23418 12314 23420
rect 12338 23418 12394 23420
rect 12098 23366 12144 23418
rect 12144 23366 12154 23418
rect 12178 23366 12208 23418
rect 12208 23366 12220 23418
rect 12220 23366 12234 23418
rect 12258 23366 12272 23418
rect 12272 23366 12284 23418
rect 12284 23366 12314 23418
rect 12338 23366 12348 23418
rect 12348 23366 12394 23418
rect 12098 23364 12154 23366
rect 12178 23364 12234 23366
rect 12258 23364 12314 23366
rect 12338 23364 12394 23366
rect 12098 22330 12154 22332
rect 12178 22330 12234 22332
rect 12258 22330 12314 22332
rect 12338 22330 12394 22332
rect 12098 22278 12144 22330
rect 12144 22278 12154 22330
rect 12178 22278 12208 22330
rect 12208 22278 12220 22330
rect 12220 22278 12234 22330
rect 12258 22278 12272 22330
rect 12272 22278 12284 22330
rect 12284 22278 12314 22330
rect 12338 22278 12348 22330
rect 12348 22278 12394 22330
rect 12098 22276 12154 22278
rect 12178 22276 12234 22278
rect 12258 22276 12314 22278
rect 12338 22276 12394 22278
rect 12098 21242 12154 21244
rect 12178 21242 12234 21244
rect 12258 21242 12314 21244
rect 12338 21242 12394 21244
rect 12098 21190 12144 21242
rect 12144 21190 12154 21242
rect 12178 21190 12208 21242
rect 12208 21190 12220 21242
rect 12220 21190 12234 21242
rect 12258 21190 12272 21242
rect 12272 21190 12284 21242
rect 12284 21190 12314 21242
rect 12338 21190 12348 21242
rect 12348 21190 12394 21242
rect 12098 21188 12154 21190
rect 12178 21188 12234 21190
rect 12258 21188 12314 21190
rect 12338 21188 12394 21190
rect 12098 20154 12154 20156
rect 12178 20154 12234 20156
rect 12258 20154 12314 20156
rect 12338 20154 12394 20156
rect 12098 20102 12144 20154
rect 12144 20102 12154 20154
rect 12178 20102 12208 20154
rect 12208 20102 12220 20154
rect 12220 20102 12234 20154
rect 12258 20102 12272 20154
rect 12272 20102 12284 20154
rect 12284 20102 12314 20154
rect 12338 20102 12348 20154
rect 12348 20102 12394 20154
rect 12098 20100 12154 20102
rect 12178 20100 12234 20102
rect 12258 20100 12314 20102
rect 12338 20100 12394 20102
rect 12098 19066 12154 19068
rect 12178 19066 12234 19068
rect 12258 19066 12314 19068
rect 12338 19066 12394 19068
rect 12098 19014 12144 19066
rect 12144 19014 12154 19066
rect 12178 19014 12208 19066
rect 12208 19014 12220 19066
rect 12220 19014 12234 19066
rect 12258 19014 12272 19066
rect 12272 19014 12284 19066
rect 12284 19014 12314 19066
rect 12338 19014 12348 19066
rect 12348 19014 12394 19066
rect 12098 19012 12154 19014
rect 12178 19012 12234 19014
rect 12258 19012 12314 19014
rect 12338 19012 12394 19014
rect 8384 15258 8440 15260
rect 8464 15258 8520 15260
rect 8544 15258 8600 15260
rect 8624 15258 8680 15260
rect 8384 15206 8430 15258
rect 8430 15206 8440 15258
rect 8464 15206 8494 15258
rect 8494 15206 8506 15258
rect 8506 15206 8520 15258
rect 8544 15206 8558 15258
rect 8558 15206 8570 15258
rect 8570 15206 8600 15258
rect 8624 15206 8634 15258
rect 8634 15206 8680 15258
rect 8384 15204 8440 15206
rect 8464 15204 8520 15206
rect 8544 15204 8600 15206
rect 8624 15204 8680 15206
rect 8384 14170 8440 14172
rect 8464 14170 8520 14172
rect 8544 14170 8600 14172
rect 8624 14170 8680 14172
rect 8384 14118 8430 14170
rect 8430 14118 8440 14170
rect 8464 14118 8494 14170
rect 8494 14118 8506 14170
rect 8506 14118 8520 14170
rect 8544 14118 8558 14170
rect 8558 14118 8570 14170
rect 8570 14118 8600 14170
rect 8624 14118 8634 14170
rect 8634 14118 8680 14170
rect 8384 14116 8440 14118
rect 8464 14116 8520 14118
rect 8544 14116 8600 14118
rect 8624 14116 8680 14118
rect 8384 13082 8440 13084
rect 8464 13082 8520 13084
rect 8544 13082 8600 13084
rect 8624 13082 8680 13084
rect 8384 13030 8430 13082
rect 8430 13030 8440 13082
rect 8464 13030 8494 13082
rect 8494 13030 8506 13082
rect 8506 13030 8520 13082
rect 8544 13030 8558 13082
rect 8558 13030 8570 13082
rect 8570 13030 8600 13082
rect 8624 13030 8634 13082
rect 8634 13030 8680 13082
rect 8384 13028 8440 13030
rect 8464 13028 8520 13030
rect 8544 13028 8600 13030
rect 8624 13028 8680 13030
rect 8384 11994 8440 11996
rect 8464 11994 8520 11996
rect 8544 11994 8600 11996
rect 8624 11994 8680 11996
rect 8384 11942 8430 11994
rect 8430 11942 8440 11994
rect 8464 11942 8494 11994
rect 8494 11942 8506 11994
rect 8506 11942 8520 11994
rect 8544 11942 8558 11994
rect 8558 11942 8570 11994
rect 8570 11942 8600 11994
rect 8624 11942 8634 11994
rect 8634 11942 8680 11994
rect 8384 11940 8440 11942
rect 8464 11940 8520 11942
rect 8544 11940 8600 11942
rect 8624 11940 8680 11942
rect 8384 10906 8440 10908
rect 8464 10906 8520 10908
rect 8544 10906 8600 10908
rect 8624 10906 8680 10908
rect 8384 10854 8430 10906
rect 8430 10854 8440 10906
rect 8464 10854 8494 10906
rect 8494 10854 8506 10906
rect 8506 10854 8520 10906
rect 8544 10854 8558 10906
rect 8558 10854 8570 10906
rect 8570 10854 8600 10906
rect 8624 10854 8634 10906
rect 8634 10854 8680 10906
rect 8384 10852 8440 10854
rect 8464 10852 8520 10854
rect 8544 10852 8600 10854
rect 8624 10852 8680 10854
rect 8384 9818 8440 9820
rect 8464 9818 8520 9820
rect 8544 9818 8600 9820
rect 8624 9818 8680 9820
rect 8384 9766 8430 9818
rect 8430 9766 8440 9818
rect 8464 9766 8494 9818
rect 8494 9766 8506 9818
rect 8506 9766 8520 9818
rect 8544 9766 8558 9818
rect 8558 9766 8570 9818
rect 8570 9766 8600 9818
rect 8624 9766 8634 9818
rect 8634 9766 8680 9818
rect 8384 9764 8440 9766
rect 8464 9764 8520 9766
rect 8544 9764 8600 9766
rect 8624 9764 8680 9766
rect 8384 8730 8440 8732
rect 8464 8730 8520 8732
rect 8544 8730 8600 8732
rect 8624 8730 8680 8732
rect 8384 8678 8430 8730
rect 8430 8678 8440 8730
rect 8464 8678 8494 8730
rect 8494 8678 8506 8730
rect 8506 8678 8520 8730
rect 8544 8678 8558 8730
rect 8558 8678 8570 8730
rect 8570 8678 8600 8730
rect 8624 8678 8634 8730
rect 8634 8678 8680 8730
rect 8384 8676 8440 8678
rect 8464 8676 8520 8678
rect 8544 8676 8600 8678
rect 8624 8676 8680 8678
rect 8384 7642 8440 7644
rect 8464 7642 8520 7644
rect 8544 7642 8600 7644
rect 8624 7642 8680 7644
rect 8384 7590 8430 7642
rect 8430 7590 8440 7642
rect 8464 7590 8494 7642
rect 8494 7590 8506 7642
rect 8506 7590 8520 7642
rect 8544 7590 8558 7642
rect 8558 7590 8570 7642
rect 8570 7590 8600 7642
rect 8624 7590 8634 7642
rect 8634 7590 8680 7642
rect 8384 7588 8440 7590
rect 8464 7588 8520 7590
rect 8544 7588 8600 7590
rect 8624 7588 8680 7590
rect 8384 6554 8440 6556
rect 8464 6554 8520 6556
rect 8544 6554 8600 6556
rect 8624 6554 8680 6556
rect 8384 6502 8430 6554
rect 8430 6502 8440 6554
rect 8464 6502 8494 6554
rect 8494 6502 8506 6554
rect 8506 6502 8520 6554
rect 8544 6502 8558 6554
rect 8558 6502 8570 6554
rect 8570 6502 8600 6554
rect 8624 6502 8634 6554
rect 8634 6502 8680 6554
rect 8384 6500 8440 6502
rect 8464 6500 8520 6502
rect 8544 6500 8600 6502
rect 8624 6500 8680 6502
rect 12098 17978 12154 17980
rect 12178 17978 12234 17980
rect 12258 17978 12314 17980
rect 12338 17978 12394 17980
rect 12098 17926 12144 17978
rect 12144 17926 12154 17978
rect 12178 17926 12208 17978
rect 12208 17926 12220 17978
rect 12220 17926 12234 17978
rect 12258 17926 12272 17978
rect 12272 17926 12284 17978
rect 12284 17926 12314 17978
rect 12338 17926 12348 17978
rect 12348 17926 12394 17978
rect 12098 17924 12154 17926
rect 12178 17924 12234 17926
rect 12258 17924 12314 17926
rect 12338 17924 12394 17926
rect 12098 16890 12154 16892
rect 12178 16890 12234 16892
rect 12258 16890 12314 16892
rect 12338 16890 12394 16892
rect 12098 16838 12144 16890
rect 12144 16838 12154 16890
rect 12178 16838 12208 16890
rect 12208 16838 12220 16890
rect 12220 16838 12234 16890
rect 12258 16838 12272 16890
rect 12272 16838 12284 16890
rect 12284 16838 12314 16890
rect 12338 16838 12348 16890
rect 12348 16838 12394 16890
rect 12098 16836 12154 16838
rect 12178 16836 12234 16838
rect 12258 16836 12314 16838
rect 12338 16836 12394 16838
rect 12098 15802 12154 15804
rect 12178 15802 12234 15804
rect 12258 15802 12314 15804
rect 12338 15802 12394 15804
rect 12098 15750 12144 15802
rect 12144 15750 12154 15802
rect 12178 15750 12208 15802
rect 12208 15750 12220 15802
rect 12220 15750 12234 15802
rect 12258 15750 12272 15802
rect 12272 15750 12284 15802
rect 12284 15750 12314 15802
rect 12338 15750 12348 15802
rect 12348 15750 12394 15802
rect 12098 15748 12154 15750
rect 12178 15748 12234 15750
rect 12258 15748 12314 15750
rect 12338 15748 12394 15750
rect 12098 14714 12154 14716
rect 12178 14714 12234 14716
rect 12258 14714 12314 14716
rect 12338 14714 12394 14716
rect 12098 14662 12144 14714
rect 12144 14662 12154 14714
rect 12178 14662 12208 14714
rect 12208 14662 12220 14714
rect 12220 14662 12234 14714
rect 12258 14662 12272 14714
rect 12272 14662 12284 14714
rect 12284 14662 12314 14714
rect 12338 14662 12348 14714
rect 12348 14662 12394 14714
rect 12098 14660 12154 14662
rect 12178 14660 12234 14662
rect 12258 14660 12314 14662
rect 12338 14660 12394 14662
rect 12098 13626 12154 13628
rect 12178 13626 12234 13628
rect 12258 13626 12314 13628
rect 12338 13626 12394 13628
rect 12098 13574 12144 13626
rect 12144 13574 12154 13626
rect 12178 13574 12208 13626
rect 12208 13574 12220 13626
rect 12220 13574 12234 13626
rect 12258 13574 12272 13626
rect 12272 13574 12284 13626
rect 12284 13574 12314 13626
rect 12338 13574 12348 13626
rect 12348 13574 12394 13626
rect 12098 13572 12154 13574
rect 12178 13572 12234 13574
rect 12258 13572 12314 13574
rect 12338 13572 12394 13574
rect 12098 12538 12154 12540
rect 12178 12538 12234 12540
rect 12258 12538 12314 12540
rect 12338 12538 12394 12540
rect 12098 12486 12144 12538
rect 12144 12486 12154 12538
rect 12178 12486 12208 12538
rect 12208 12486 12220 12538
rect 12220 12486 12234 12538
rect 12258 12486 12272 12538
rect 12272 12486 12284 12538
rect 12284 12486 12314 12538
rect 12338 12486 12348 12538
rect 12348 12486 12394 12538
rect 12098 12484 12154 12486
rect 12178 12484 12234 12486
rect 12258 12484 12314 12486
rect 12338 12484 12394 12486
rect 12098 11450 12154 11452
rect 12178 11450 12234 11452
rect 12258 11450 12314 11452
rect 12338 11450 12394 11452
rect 12098 11398 12144 11450
rect 12144 11398 12154 11450
rect 12178 11398 12208 11450
rect 12208 11398 12220 11450
rect 12220 11398 12234 11450
rect 12258 11398 12272 11450
rect 12272 11398 12284 11450
rect 12284 11398 12314 11450
rect 12338 11398 12348 11450
rect 12348 11398 12394 11450
rect 12098 11396 12154 11398
rect 12178 11396 12234 11398
rect 12258 11396 12314 11398
rect 12338 11396 12394 11398
rect 12098 10362 12154 10364
rect 12178 10362 12234 10364
rect 12258 10362 12314 10364
rect 12338 10362 12394 10364
rect 12098 10310 12144 10362
rect 12144 10310 12154 10362
rect 12178 10310 12208 10362
rect 12208 10310 12220 10362
rect 12220 10310 12234 10362
rect 12258 10310 12272 10362
rect 12272 10310 12284 10362
rect 12284 10310 12314 10362
rect 12338 10310 12348 10362
rect 12348 10310 12394 10362
rect 12098 10308 12154 10310
rect 12178 10308 12234 10310
rect 12258 10308 12314 10310
rect 12338 10308 12394 10310
rect 12098 9274 12154 9276
rect 12178 9274 12234 9276
rect 12258 9274 12314 9276
rect 12338 9274 12394 9276
rect 12098 9222 12144 9274
rect 12144 9222 12154 9274
rect 12178 9222 12208 9274
rect 12208 9222 12220 9274
rect 12220 9222 12234 9274
rect 12258 9222 12272 9274
rect 12272 9222 12284 9274
rect 12284 9222 12314 9274
rect 12338 9222 12348 9274
rect 12348 9222 12394 9274
rect 12098 9220 12154 9222
rect 12178 9220 12234 9222
rect 12258 9220 12314 9222
rect 12338 9220 12394 9222
rect 12098 8186 12154 8188
rect 12178 8186 12234 8188
rect 12258 8186 12314 8188
rect 12338 8186 12394 8188
rect 12098 8134 12144 8186
rect 12144 8134 12154 8186
rect 12178 8134 12208 8186
rect 12208 8134 12220 8186
rect 12220 8134 12234 8186
rect 12258 8134 12272 8186
rect 12272 8134 12284 8186
rect 12284 8134 12314 8186
rect 12338 8134 12348 8186
rect 12348 8134 12394 8186
rect 12098 8132 12154 8134
rect 12178 8132 12234 8134
rect 12258 8132 12314 8134
rect 12338 8132 12394 8134
rect 12098 7098 12154 7100
rect 12178 7098 12234 7100
rect 12258 7098 12314 7100
rect 12338 7098 12394 7100
rect 12098 7046 12144 7098
rect 12144 7046 12154 7098
rect 12178 7046 12208 7098
rect 12208 7046 12220 7098
rect 12220 7046 12234 7098
rect 12258 7046 12272 7098
rect 12272 7046 12284 7098
rect 12284 7046 12314 7098
rect 12338 7046 12348 7098
rect 12348 7046 12394 7098
rect 12098 7044 12154 7046
rect 12178 7044 12234 7046
rect 12258 7044 12314 7046
rect 12338 7044 12394 7046
rect 4670 6010 4726 6012
rect 4750 6010 4806 6012
rect 4830 6010 4886 6012
rect 4910 6010 4966 6012
rect 4670 5958 4716 6010
rect 4716 5958 4726 6010
rect 4750 5958 4780 6010
rect 4780 5958 4792 6010
rect 4792 5958 4806 6010
rect 4830 5958 4844 6010
rect 4844 5958 4856 6010
rect 4856 5958 4886 6010
rect 4910 5958 4920 6010
rect 4920 5958 4966 6010
rect 4670 5956 4726 5958
rect 4750 5956 4806 5958
rect 4830 5956 4886 5958
rect 4910 5956 4966 5958
rect 12098 6010 12154 6012
rect 12178 6010 12234 6012
rect 12258 6010 12314 6012
rect 12338 6010 12394 6012
rect 12098 5958 12144 6010
rect 12144 5958 12154 6010
rect 12178 5958 12208 6010
rect 12208 5958 12220 6010
rect 12220 5958 12234 6010
rect 12258 5958 12272 6010
rect 12272 5958 12284 6010
rect 12284 5958 12314 6010
rect 12338 5958 12348 6010
rect 12348 5958 12394 6010
rect 12098 5956 12154 5958
rect 12178 5956 12234 5958
rect 12258 5956 12314 5958
rect 12338 5956 12394 5958
rect 23240 29402 23296 29404
rect 23320 29402 23376 29404
rect 23400 29402 23456 29404
rect 23480 29402 23536 29404
rect 23240 29350 23286 29402
rect 23286 29350 23296 29402
rect 23320 29350 23350 29402
rect 23350 29350 23362 29402
rect 23362 29350 23376 29402
rect 23400 29350 23414 29402
rect 23414 29350 23426 29402
rect 23426 29350 23456 29402
rect 23480 29350 23490 29402
rect 23490 29350 23536 29402
rect 23240 29348 23296 29350
rect 23320 29348 23376 29350
rect 23400 29348 23456 29350
rect 23480 29348 23536 29350
rect 31022 29688 31078 29744
rect 30668 29402 30724 29404
rect 30748 29402 30804 29404
rect 30828 29402 30884 29404
rect 30908 29402 30964 29404
rect 30668 29350 30714 29402
rect 30714 29350 30724 29402
rect 30748 29350 30778 29402
rect 30778 29350 30790 29402
rect 30790 29350 30804 29402
rect 30828 29350 30842 29402
rect 30842 29350 30854 29402
rect 30854 29350 30884 29402
rect 30908 29350 30918 29402
rect 30918 29350 30964 29402
rect 30668 29348 30724 29350
rect 30748 29348 30804 29350
rect 30828 29348 30884 29350
rect 30908 29348 30964 29350
rect 19526 28858 19582 28860
rect 19606 28858 19662 28860
rect 19686 28858 19742 28860
rect 19766 28858 19822 28860
rect 19526 28806 19572 28858
rect 19572 28806 19582 28858
rect 19606 28806 19636 28858
rect 19636 28806 19648 28858
rect 19648 28806 19662 28858
rect 19686 28806 19700 28858
rect 19700 28806 19712 28858
rect 19712 28806 19742 28858
rect 19766 28806 19776 28858
rect 19776 28806 19822 28858
rect 19526 28804 19582 28806
rect 19606 28804 19662 28806
rect 19686 28804 19742 28806
rect 19766 28804 19822 28806
rect 15812 28314 15868 28316
rect 15892 28314 15948 28316
rect 15972 28314 16028 28316
rect 16052 28314 16108 28316
rect 15812 28262 15858 28314
rect 15858 28262 15868 28314
rect 15892 28262 15922 28314
rect 15922 28262 15934 28314
rect 15934 28262 15948 28314
rect 15972 28262 15986 28314
rect 15986 28262 15998 28314
rect 15998 28262 16028 28314
rect 16052 28262 16062 28314
rect 16062 28262 16108 28314
rect 15812 28260 15868 28262
rect 15892 28260 15948 28262
rect 15972 28260 16028 28262
rect 16052 28260 16108 28262
rect 15812 27226 15868 27228
rect 15892 27226 15948 27228
rect 15972 27226 16028 27228
rect 16052 27226 16108 27228
rect 15812 27174 15858 27226
rect 15858 27174 15868 27226
rect 15892 27174 15922 27226
rect 15922 27174 15934 27226
rect 15934 27174 15948 27226
rect 15972 27174 15986 27226
rect 15986 27174 15998 27226
rect 15998 27174 16028 27226
rect 16052 27174 16062 27226
rect 16062 27174 16108 27226
rect 15812 27172 15868 27174
rect 15892 27172 15948 27174
rect 15972 27172 16028 27174
rect 16052 27172 16108 27174
rect 15812 26138 15868 26140
rect 15892 26138 15948 26140
rect 15972 26138 16028 26140
rect 16052 26138 16108 26140
rect 15812 26086 15858 26138
rect 15858 26086 15868 26138
rect 15892 26086 15922 26138
rect 15922 26086 15934 26138
rect 15934 26086 15948 26138
rect 15972 26086 15986 26138
rect 15986 26086 15998 26138
rect 15998 26086 16028 26138
rect 16052 26086 16062 26138
rect 16062 26086 16108 26138
rect 15812 26084 15868 26086
rect 15892 26084 15948 26086
rect 15972 26084 16028 26086
rect 16052 26084 16108 26086
rect 15812 25050 15868 25052
rect 15892 25050 15948 25052
rect 15972 25050 16028 25052
rect 16052 25050 16108 25052
rect 15812 24998 15858 25050
rect 15858 24998 15868 25050
rect 15892 24998 15922 25050
rect 15922 24998 15934 25050
rect 15934 24998 15948 25050
rect 15972 24998 15986 25050
rect 15986 24998 15998 25050
rect 15998 24998 16028 25050
rect 16052 24998 16062 25050
rect 16062 24998 16108 25050
rect 15812 24996 15868 24998
rect 15892 24996 15948 24998
rect 15972 24996 16028 24998
rect 16052 24996 16108 24998
rect 15812 23962 15868 23964
rect 15892 23962 15948 23964
rect 15972 23962 16028 23964
rect 16052 23962 16108 23964
rect 15812 23910 15858 23962
rect 15858 23910 15868 23962
rect 15892 23910 15922 23962
rect 15922 23910 15934 23962
rect 15934 23910 15948 23962
rect 15972 23910 15986 23962
rect 15986 23910 15998 23962
rect 15998 23910 16028 23962
rect 16052 23910 16062 23962
rect 16062 23910 16108 23962
rect 15812 23908 15868 23910
rect 15892 23908 15948 23910
rect 15972 23908 16028 23910
rect 16052 23908 16108 23910
rect 15812 22874 15868 22876
rect 15892 22874 15948 22876
rect 15972 22874 16028 22876
rect 16052 22874 16108 22876
rect 15812 22822 15858 22874
rect 15858 22822 15868 22874
rect 15892 22822 15922 22874
rect 15922 22822 15934 22874
rect 15934 22822 15948 22874
rect 15972 22822 15986 22874
rect 15986 22822 15998 22874
rect 15998 22822 16028 22874
rect 16052 22822 16062 22874
rect 16062 22822 16108 22874
rect 15812 22820 15868 22822
rect 15892 22820 15948 22822
rect 15972 22820 16028 22822
rect 16052 22820 16108 22822
rect 15812 21786 15868 21788
rect 15892 21786 15948 21788
rect 15972 21786 16028 21788
rect 16052 21786 16108 21788
rect 15812 21734 15858 21786
rect 15858 21734 15868 21786
rect 15892 21734 15922 21786
rect 15922 21734 15934 21786
rect 15934 21734 15948 21786
rect 15972 21734 15986 21786
rect 15986 21734 15998 21786
rect 15998 21734 16028 21786
rect 16052 21734 16062 21786
rect 16062 21734 16108 21786
rect 15812 21732 15868 21734
rect 15892 21732 15948 21734
rect 15972 21732 16028 21734
rect 16052 21732 16108 21734
rect 15812 20698 15868 20700
rect 15892 20698 15948 20700
rect 15972 20698 16028 20700
rect 16052 20698 16108 20700
rect 15812 20646 15858 20698
rect 15858 20646 15868 20698
rect 15892 20646 15922 20698
rect 15922 20646 15934 20698
rect 15934 20646 15948 20698
rect 15972 20646 15986 20698
rect 15986 20646 15998 20698
rect 15998 20646 16028 20698
rect 16052 20646 16062 20698
rect 16062 20646 16108 20698
rect 15812 20644 15868 20646
rect 15892 20644 15948 20646
rect 15972 20644 16028 20646
rect 16052 20644 16108 20646
rect 15812 19610 15868 19612
rect 15892 19610 15948 19612
rect 15972 19610 16028 19612
rect 16052 19610 16108 19612
rect 15812 19558 15858 19610
rect 15858 19558 15868 19610
rect 15892 19558 15922 19610
rect 15922 19558 15934 19610
rect 15934 19558 15948 19610
rect 15972 19558 15986 19610
rect 15986 19558 15998 19610
rect 15998 19558 16028 19610
rect 16052 19558 16062 19610
rect 16062 19558 16108 19610
rect 15812 19556 15868 19558
rect 15892 19556 15948 19558
rect 15972 19556 16028 19558
rect 16052 19556 16108 19558
rect 15812 18522 15868 18524
rect 15892 18522 15948 18524
rect 15972 18522 16028 18524
rect 16052 18522 16108 18524
rect 15812 18470 15858 18522
rect 15858 18470 15868 18522
rect 15892 18470 15922 18522
rect 15922 18470 15934 18522
rect 15934 18470 15948 18522
rect 15972 18470 15986 18522
rect 15986 18470 15998 18522
rect 15998 18470 16028 18522
rect 16052 18470 16062 18522
rect 16062 18470 16108 18522
rect 15812 18468 15868 18470
rect 15892 18468 15948 18470
rect 15972 18468 16028 18470
rect 16052 18468 16108 18470
rect 15812 17434 15868 17436
rect 15892 17434 15948 17436
rect 15972 17434 16028 17436
rect 16052 17434 16108 17436
rect 15812 17382 15858 17434
rect 15858 17382 15868 17434
rect 15892 17382 15922 17434
rect 15922 17382 15934 17434
rect 15934 17382 15948 17434
rect 15972 17382 15986 17434
rect 15986 17382 15998 17434
rect 15998 17382 16028 17434
rect 16052 17382 16062 17434
rect 16062 17382 16108 17434
rect 15812 17380 15868 17382
rect 15892 17380 15948 17382
rect 15972 17380 16028 17382
rect 16052 17380 16108 17382
rect 15812 16346 15868 16348
rect 15892 16346 15948 16348
rect 15972 16346 16028 16348
rect 16052 16346 16108 16348
rect 15812 16294 15858 16346
rect 15858 16294 15868 16346
rect 15892 16294 15922 16346
rect 15922 16294 15934 16346
rect 15934 16294 15948 16346
rect 15972 16294 15986 16346
rect 15986 16294 15998 16346
rect 15998 16294 16028 16346
rect 16052 16294 16062 16346
rect 16062 16294 16108 16346
rect 15812 16292 15868 16294
rect 15892 16292 15948 16294
rect 15972 16292 16028 16294
rect 16052 16292 16108 16294
rect 15812 15258 15868 15260
rect 15892 15258 15948 15260
rect 15972 15258 16028 15260
rect 16052 15258 16108 15260
rect 15812 15206 15858 15258
rect 15858 15206 15868 15258
rect 15892 15206 15922 15258
rect 15922 15206 15934 15258
rect 15934 15206 15948 15258
rect 15972 15206 15986 15258
rect 15986 15206 15998 15258
rect 15998 15206 16028 15258
rect 16052 15206 16062 15258
rect 16062 15206 16108 15258
rect 15812 15204 15868 15206
rect 15892 15204 15948 15206
rect 15972 15204 16028 15206
rect 16052 15204 16108 15206
rect 15812 14170 15868 14172
rect 15892 14170 15948 14172
rect 15972 14170 16028 14172
rect 16052 14170 16108 14172
rect 15812 14118 15858 14170
rect 15858 14118 15868 14170
rect 15892 14118 15922 14170
rect 15922 14118 15934 14170
rect 15934 14118 15948 14170
rect 15972 14118 15986 14170
rect 15986 14118 15998 14170
rect 15998 14118 16028 14170
rect 16052 14118 16062 14170
rect 16062 14118 16108 14170
rect 15812 14116 15868 14118
rect 15892 14116 15948 14118
rect 15972 14116 16028 14118
rect 16052 14116 16108 14118
rect 19526 27770 19582 27772
rect 19606 27770 19662 27772
rect 19686 27770 19742 27772
rect 19766 27770 19822 27772
rect 19526 27718 19572 27770
rect 19572 27718 19582 27770
rect 19606 27718 19636 27770
rect 19636 27718 19648 27770
rect 19648 27718 19662 27770
rect 19686 27718 19700 27770
rect 19700 27718 19712 27770
rect 19712 27718 19742 27770
rect 19766 27718 19776 27770
rect 19776 27718 19822 27770
rect 19526 27716 19582 27718
rect 19606 27716 19662 27718
rect 19686 27716 19742 27718
rect 19766 27716 19822 27718
rect 19526 26682 19582 26684
rect 19606 26682 19662 26684
rect 19686 26682 19742 26684
rect 19766 26682 19822 26684
rect 19526 26630 19572 26682
rect 19572 26630 19582 26682
rect 19606 26630 19636 26682
rect 19636 26630 19648 26682
rect 19648 26630 19662 26682
rect 19686 26630 19700 26682
rect 19700 26630 19712 26682
rect 19712 26630 19742 26682
rect 19766 26630 19776 26682
rect 19776 26630 19822 26682
rect 19526 26628 19582 26630
rect 19606 26628 19662 26630
rect 19686 26628 19742 26630
rect 19766 26628 19822 26630
rect 19526 25594 19582 25596
rect 19606 25594 19662 25596
rect 19686 25594 19742 25596
rect 19766 25594 19822 25596
rect 19526 25542 19572 25594
rect 19572 25542 19582 25594
rect 19606 25542 19636 25594
rect 19636 25542 19648 25594
rect 19648 25542 19662 25594
rect 19686 25542 19700 25594
rect 19700 25542 19712 25594
rect 19712 25542 19742 25594
rect 19766 25542 19776 25594
rect 19776 25542 19822 25594
rect 19526 25540 19582 25542
rect 19606 25540 19662 25542
rect 19686 25540 19742 25542
rect 19766 25540 19822 25542
rect 19526 24506 19582 24508
rect 19606 24506 19662 24508
rect 19686 24506 19742 24508
rect 19766 24506 19822 24508
rect 19526 24454 19572 24506
rect 19572 24454 19582 24506
rect 19606 24454 19636 24506
rect 19636 24454 19648 24506
rect 19648 24454 19662 24506
rect 19686 24454 19700 24506
rect 19700 24454 19712 24506
rect 19712 24454 19742 24506
rect 19766 24454 19776 24506
rect 19776 24454 19822 24506
rect 19526 24452 19582 24454
rect 19606 24452 19662 24454
rect 19686 24452 19742 24454
rect 19766 24452 19822 24454
rect 19526 23418 19582 23420
rect 19606 23418 19662 23420
rect 19686 23418 19742 23420
rect 19766 23418 19822 23420
rect 19526 23366 19572 23418
rect 19572 23366 19582 23418
rect 19606 23366 19636 23418
rect 19636 23366 19648 23418
rect 19648 23366 19662 23418
rect 19686 23366 19700 23418
rect 19700 23366 19712 23418
rect 19712 23366 19742 23418
rect 19766 23366 19776 23418
rect 19776 23366 19822 23418
rect 19526 23364 19582 23366
rect 19606 23364 19662 23366
rect 19686 23364 19742 23366
rect 19766 23364 19822 23366
rect 19526 22330 19582 22332
rect 19606 22330 19662 22332
rect 19686 22330 19742 22332
rect 19766 22330 19822 22332
rect 19526 22278 19572 22330
rect 19572 22278 19582 22330
rect 19606 22278 19636 22330
rect 19636 22278 19648 22330
rect 19648 22278 19662 22330
rect 19686 22278 19700 22330
rect 19700 22278 19712 22330
rect 19712 22278 19742 22330
rect 19766 22278 19776 22330
rect 19776 22278 19822 22330
rect 19526 22276 19582 22278
rect 19606 22276 19662 22278
rect 19686 22276 19742 22278
rect 19766 22276 19822 22278
rect 19526 21242 19582 21244
rect 19606 21242 19662 21244
rect 19686 21242 19742 21244
rect 19766 21242 19822 21244
rect 19526 21190 19572 21242
rect 19572 21190 19582 21242
rect 19606 21190 19636 21242
rect 19636 21190 19648 21242
rect 19648 21190 19662 21242
rect 19686 21190 19700 21242
rect 19700 21190 19712 21242
rect 19712 21190 19742 21242
rect 19766 21190 19776 21242
rect 19776 21190 19822 21242
rect 19526 21188 19582 21190
rect 19606 21188 19662 21190
rect 19686 21188 19742 21190
rect 19766 21188 19822 21190
rect 19526 20154 19582 20156
rect 19606 20154 19662 20156
rect 19686 20154 19742 20156
rect 19766 20154 19822 20156
rect 19526 20102 19572 20154
rect 19572 20102 19582 20154
rect 19606 20102 19636 20154
rect 19636 20102 19648 20154
rect 19648 20102 19662 20154
rect 19686 20102 19700 20154
rect 19700 20102 19712 20154
rect 19712 20102 19742 20154
rect 19766 20102 19776 20154
rect 19776 20102 19822 20154
rect 19526 20100 19582 20102
rect 19606 20100 19662 20102
rect 19686 20100 19742 20102
rect 19766 20100 19822 20102
rect 19526 19066 19582 19068
rect 19606 19066 19662 19068
rect 19686 19066 19742 19068
rect 19766 19066 19822 19068
rect 19526 19014 19572 19066
rect 19572 19014 19582 19066
rect 19606 19014 19636 19066
rect 19636 19014 19648 19066
rect 19648 19014 19662 19066
rect 19686 19014 19700 19066
rect 19700 19014 19712 19066
rect 19712 19014 19742 19066
rect 19766 19014 19776 19066
rect 19776 19014 19822 19066
rect 19526 19012 19582 19014
rect 19606 19012 19662 19014
rect 19686 19012 19742 19014
rect 19766 19012 19822 19014
rect 19526 17978 19582 17980
rect 19606 17978 19662 17980
rect 19686 17978 19742 17980
rect 19766 17978 19822 17980
rect 19526 17926 19572 17978
rect 19572 17926 19582 17978
rect 19606 17926 19636 17978
rect 19636 17926 19648 17978
rect 19648 17926 19662 17978
rect 19686 17926 19700 17978
rect 19700 17926 19712 17978
rect 19712 17926 19742 17978
rect 19766 17926 19776 17978
rect 19776 17926 19822 17978
rect 19526 17924 19582 17926
rect 19606 17924 19662 17926
rect 19686 17924 19742 17926
rect 19766 17924 19822 17926
rect 19526 16890 19582 16892
rect 19606 16890 19662 16892
rect 19686 16890 19742 16892
rect 19766 16890 19822 16892
rect 19526 16838 19572 16890
rect 19572 16838 19582 16890
rect 19606 16838 19636 16890
rect 19636 16838 19648 16890
rect 19648 16838 19662 16890
rect 19686 16838 19700 16890
rect 19700 16838 19712 16890
rect 19712 16838 19742 16890
rect 19766 16838 19776 16890
rect 19776 16838 19822 16890
rect 19526 16836 19582 16838
rect 19606 16836 19662 16838
rect 19686 16836 19742 16838
rect 19766 16836 19822 16838
rect 15812 13082 15868 13084
rect 15892 13082 15948 13084
rect 15972 13082 16028 13084
rect 16052 13082 16108 13084
rect 15812 13030 15858 13082
rect 15858 13030 15868 13082
rect 15892 13030 15922 13082
rect 15922 13030 15934 13082
rect 15934 13030 15948 13082
rect 15972 13030 15986 13082
rect 15986 13030 15998 13082
rect 15998 13030 16028 13082
rect 16052 13030 16062 13082
rect 16062 13030 16108 13082
rect 15812 13028 15868 13030
rect 15892 13028 15948 13030
rect 15972 13028 16028 13030
rect 16052 13028 16108 13030
rect 15812 11994 15868 11996
rect 15892 11994 15948 11996
rect 15972 11994 16028 11996
rect 16052 11994 16108 11996
rect 15812 11942 15858 11994
rect 15858 11942 15868 11994
rect 15892 11942 15922 11994
rect 15922 11942 15934 11994
rect 15934 11942 15948 11994
rect 15972 11942 15986 11994
rect 15986 11942 15998 11994
rect 15998 11942 16028 11994
rect 16052 11942 16062 11994
rect 16062 11942 16108 11994
rect 15812 11940 15868 11942
rect 15892 11940 15948 11942
rect 15972 11940 16028 11942
rect 16052 11940 16108 11942
rect 15812 10906 15868 10908
rect 15892 10906 15948 10908
rect 15972 10906 16028 10908
rect 16052 10906 16108 10908
rect 15812 10854 15858 10906
rect 15858 10854 15868 10906
rect 15892 10854 15922 10906
rect 15922 10854 15934 10906
rect 15934 10854 15948 10906
rect 15972 10854 15986 10906
rect 15986 10854 15998 10906
rect 15998 10854 16028 10906
rect 16052 10854 16062 10906
rect 16062 10854 16108 10906
rect 15812 10852 15868 10854
rect 15892 10852 15948 10854
rect 15972 10852 16028 10854
rect 16052 10852 16108 10854
rect 15812 9818 15868 9820
rect 15892 9818 15948 9820
rect 15972 9818 16028 9820
rect 16052 9818 16108 9820
rect 15812 9766 15858 9818
rect 15858 9766 15868 9818
rect 15892 9766 15922 9818
rect 15922 9766 15934 9818
rect 15934 9766 15948 9818
rect 15972 9766 15986 9818
rect 15986 9766 15998 9818
rect 15998 9766 16028 9818
rect 16052 9766 16062 9818
rect 16062 9766 16108 9818
rect 15812 9764 15868 9766
rect 15892 9764 15948 9766
rect 15972 9764 16028 9766
rect 16052 9764 16108 9766
rect 15812 8730 15868 8732
rect 15892 8730 15948 8732
rect 15972 8730 16028 8732
rect 16052 8730 16108 8732
rect 15812 8678 15858 8730
rect 15858 8678 15868 8730
rect 15892 8678 15922 8730
rect 15922 8678 15934 8730
rect 15934 8678 15948 8730
rect 15972 8678 15986 8730
rect 15986 8678 15998 8730
rect 15998 8678 16028 8730
rect 16052 8678 16062 8730
rect 16062 8678 16108 8730
rect 15812 8676 15868 8678
rect 15892 8676 15948 8678
rect 15972 8676 16028 8678
rect 16052 8676 16108 8678
rect 15812 7642 15868 7644
rect 15892 7642 15948 7644
rect 15972 7642 16028 7644
rect 16052 7642 16108 7644
rect 15812 7590 15858 7642
rect 15858 7590 15868 7642
rect 15892 7590 15922 7642
rect 15922 7590 15934 7642
rect 15934 7590 15948 7642
rect 15972 7590 15986 7642
rect 15986 7590 15998 7642
rect 15998 7590 16028 7642
rect 16052 7590 16062 7642
rect 16062 7590 16108 7642
rect 15812 7588 15868 7590
rect 15892 7588 15948 7590
rect 15972 7588 16028 7590
rect 16052 7588 16108 7590
rect 8384 5466 8440 5468
rect 8464 5466 8520 5468
rect 8544 5466 8600 5468
rect 8624 5466 8680 5468
rect 8384 5414 8430 5466
rect 8430 5414 8440 5466
rect 8464 5414 8494 5466
rect 8494 5414 8506 5466
rect 8506 5414 8520 5466
rect 8544 5414 8558 5466
rect 8558 5414 8570 5466
rect 8570 5414 8600 5466
rect 8624 5414 8634 5466
rect 8634 5414 8680 5466
rect 8384 5412 8440 5414
rect 8464 5412 8520 5414
rect 8544 5412 8600 5414
rect 8624 5412 8680 5414
rect 19526 15802 19582 15804
rect 19606 15802 19662 15804
rect 19686 15802 19742 15804
rect 19766 15802 19822 15804
rect 19526 15750 19572 15802
rect 19572 15750 19582 15802
rect 19606 15750 19636 15802
rect 19636 15750 19648 15802
rect 19648 15750 19662 15802
rect 19686 15750 19700 15802
rect 19700 15750 19712 15802
rect 19712 15750 19742 15802
rect 19766 15750 19776 15802
rect 19776 15750 19822 15802
rect 19526 15748 19582 15750
rect 19606 15748 19662 15750
rect 19686 15748 19742 15750
rect 19766 15748 19822 15750
rect 23240 28314 23296 28316
rect 23320 28314 23376 28316
rect 23400 28314 23456 28316
rect 23480 28314 23536 28316
rect 23240 28262 23286 28314
rect 23286 28262 23296 28314
rect 23320 28262 23350 28314
rect 23350 28262 23362 28314
rect 23362 28262 23376 28314
rect 23400 28262 23414 28314
rect 23414 28262 23426 28314
rect 23426 28262 23456 28314
rect 23480 28262 23490 28314
rect 23490 28262 23536 28314
rect 23240 28260 23296 28262
rect 23320 28260 23376 28262
rect 23400 28260 23456 28262
rect 23480 28260 23536 28262
rect 23240 27226 23296 27228
rect 23320 27226 23376 27228
rect 23400 27226 23456 27228
rect 23480 27226 23536 27228
rect 23240 27174 23286 27226
rect 23286 27174 23296 27226
rect 23320 27174 23350 27226
rect 23350 27174 23362 27226
rect 23362 27174 23376 27226
rect 23400 27174 23414 27226
rect 23414 27174 23426 27226
rect 23426 27174 23456 27226
rect 23480 27174 23490 27226
rect 23490 27174 23536 27226
rect 23240 27172 23296 27174
rect 23320 27172 23376 27174
rect 23400 27172 23456 27174
rect 23480 27172 23536 27174
rect 23240 26138 23296 26140
rect 23320 26138 23376 26140
rect 23400 26138 23456 26140
rect 23480 26138 23536 26140
rect 23240 26086 23286 26138
rect 23286 26086 23296 26138
rect 23320 26086 23350 26138
rect 23350 26086 23362 26138
rect 23362 26086 23376 26138
rect 23400 26086 23414 26138
rect 23414 26086 23426 26138
rect 23426 26086 23456 26138
rect 23480 26086 23490 26138
rect 23490 26086 23536 26138
rect 23240 26084 23296 26086
rect 23320 26084 23376 26086
rect 23400 26084 23456 26086
rect 23480 26084 23536 26086
rect 23240 25050 23296 25052
rect 23320 25050 23376 25052
rect 23400 25050 23456 25052
rect 23480 25050 23536 25052
rect 23240 24998 23286 25050
rect 23286 24998 23296 25050
rect 23320 24998 23350 25050
rect 23350 24998 23362 25050
rect 23362 24998 23376 25050
rect 23400 24998 23414 25050
rect 23414 24998 23426 25050
rect 23426 24998 23456 25050
rect 23480 24998 23490 25050
rect 23490 24998 23536 25050
rect 23240 24996 23296 24998
rect 23320 24996 23376 24998
rect 23400 24996 23456 24998
rect 23480 24996 23536 24998
rect 23240 23962 23296 23964
rect 23320 23962 23376 23964
rect 23400 23962 23456 23964
rect 23480 23962 23536 23964
rect 23240 23910 23286 23962
rect 23286 23910 23296 23962
rect 23320 23910 23350 23962
rect 23350 23910 23362 23962
rect 23362 23910 23376 23962
rect 23400 23910 23414 23962
rect 23414 23910 23426 23962
rect 23426 23910 23456 23962
rect 23480 23910 23490 23962
rect 23490 23910 23536 23962
rect 23240 23908 23296 23910
rect 23320 23908 23376 23910
rect 23400 23908 23456 23910
rect 23480 23908 23536 23910
rect 23240 22874 23296 22876
rect 23320 22874 23376 22876
rect 23400 22874 23456 22876
rect 23480 22874 23536 22876
rect 23240 22822 23286 22874
rect 23286 22822 23296 22874
rect 23320 22822 23350 22874
rect 23350 22822 23362 22874
rect 23362 22822 23376 22874
rect 23400 22822 23414 22874
rect 23414 22822 23426 22874
rect 23426 22822 23456 22874
rect 23480 22822 23490 22874
rect 23490 22822 23536 22874
rect 23240 22820 23296 22822
rect 23320 22820 23376 22822
rect 23400 22820 23456 22822
rect 23480 22820 23536 22822
rect 23240 21786 23296 21788
rect 23320 21786 23376 21788
rect 23400 21786 23456 21788
rect 23480 21786 23536 21788
rect 23240 21734 23286 21786
rect 23286 21734 23296 21786
rect 23320 21734 23350 21786
rect 23350 21734 23362 21786
rect 23362 21734 23376 21786
rect 23400 21734 23414 21786
rect 23414 21734 23426 21786
rect 23426 21734 23456 21786
rect 23480 21734 23490 21786
rect 23490 21734 23536 21786
rect 23240 21732 23296 21734
rect 23320 21732 23376 21734
rect 23400 21732 23456 21734
rect 23480 21732 23536 21734
rect 23240 20698 23296 20700
rect 23320 20698 23376 20700
rect 23400 20698 23456 20700
rect 23480 20698 23536 20700
rect 23240 20646 23286 20698
rect 23286 20646 23296 20698
rect 23320 20646 23350 20698
rect 23350 20646 23362 20698
rect 23362 20646 23376 20698
rect 23400 20646 23414 20698
rect 23414 20646 23426 20698
rect 23426 20646 23456 20698
rect 23480 20646 23490 20698
rect 23490 20646 23536 20698
rect 23240 20644 23296 20646
rect 23320 20644 23376 20646
rect 23400 20644 23456 20646
rect 23480 20644 23536 20646
rect 23240 19610 23296 19612
rect 23320 19610 23376 19612
rect 23400 19610 23456 19612
rect 23480 19610 23536 19612
rect 23240 19558 23286 19610
rect 23286 19558 23296 19610
rect 23320 19558 23350 19610
rect 23350 19558 23362 19610
rect 23362 19558 23376 19610
rect 23400 19558 23414 19610
rect 23414 19558 23426 19610
rect 23426 19558 23456 19610
rect 23480 19558 23490 19610
rect 23490 19558 23536 19610
rect 23240 19556 23296 19558
rect 23320 19556 23376 19558
rect 23400 19556 23456 19558
rect 23480 19556 23536 19558
rect 23240 18522 23296 18524
rect 23320 18522 23376 18524
rect 23400 18522 23456 18524
rect 23480 18522 23536 18524
rect 23240 18470 23286 18522
rect 23286 18470 23296 18522
rect 23320 18470 23350 18522
rect 23350 18470 23362 18522
rect 23362 18470 23376 18522
rect 23400 18470 23414 18522
rect 23414 18470 23426 18522
rect 23426 18470 23456 18522
rect 23480 18470 23490 18522
rect 23490 18470 23536 18522
rect 23240 18468 23296 18470
rect 23320 18468 23376 18470
rect 23400 18468 23456 18470
rect 23480 18468 23536 18470
rect 19526 14714 19582 14716
rect 19606 14714 19662 14716
rect 19686 14714 19742 14716
rect 19766 14714 19822 14716
rect 19526 14662 19572 14714
rect 19572 14662 19582 14714
rect 19606 14662 19636 14714
rect 19636 14662 19648 14714
rect 19648 14662 19662 14714
rect 19686 14662 19700 14714
rect 19700 14662 19712 14714
rect 19712 14662 19742 14714
rect 19766 14662 19776 14714
rect 19776 14662 19822 14714
rect 19526 14660 19582 14662
rect 19606 14660 19662 14662
rect 19686 14660 19742 14662
rect 19766 14660 19822 14662
rect 23240 17434 23296 17436
rect 23320 17434 23376 17436
rect 23400 17434 23456 17436
rect 23480 17434 23536 17436
rect 23240 17382 23286 17434
rect 23286 17382 23296 17434
rect 23320 17382 23350 17434
rect 23350 17382 23362 17434
rect 23362 17382 23376 17434
rect 23400 17382 23414 17434
rect 23414 17382 23426 17434
rect 23426 17382 23456 17434
rect 23480 17382 23490 17434
rect 23490 17382 23536 17434
rect 23240 17380 23296 17382
rect 23320 17380 23376 17382
rect 23400 17380 23456 17382
rect 23480 17380 23536 17382
rect 19526 13626 19582 13628
rect 19606 13626 19662 13628
rect 19686 13626 19742 13628
rect 19766 13626 19822 13628
rect 19526 13574 19572 13626
rect 19572 13574 19582 13626
rect 19606 13574 19636 13626
rect 19636 13574 19648 13626
rect 19648 13574 19662 13626
rect 19686 13574 19700 13626
rect 19700 13574 19712 13626
rect 19712 13574 19742 13626
rect 19766 13574 19776 13626
rect 19776 13574 19822 13626
rect 19526 13572 19582 13574
rect 19606 13572 19662 13574
rect 19686 13572 19742 13574
rect 19766 13572 19822 13574
rect 19526 12538 19582 12540
rect 19606 12538 19662 12540
rect 19686 12538 19742 12540
rect 19766 12538 19822 12540
rect 19526 12486 19572 12538
rect 19572 12486 19582 12538
rect 19606 12486 19636 12538
rect 19636 12486 19648 12538
rect 19648 12486 19662 12538
rect 19686 12486 19700 12538
rect 19700 12486 19712 12538
rect 19712 12486 19742 12538
rect 19766 12486 19776 12538
rect 19776 12486 19822 12538
rect 19526 12484 19582 12486
rect 19606 12484 19662 12486
rect 19686 12484 19742 12486
rect 19766 12484 19822 12486
rect 19526 11450 19582 11452
rect 19606 11450 19662 11452
rect 19686 11450 19742 11452
rect 19766 11450 19822 11452
rect 19526 11398 19572 11450
rect 19572 11398 19582 11450
rect 19606 11398 19636 11450
rect 19636 11398 19648 11450
rect 19648 11398 19662 11450
rect 19686 11398 19700 11450
rect 19700 11398 19712 11450
rect 19712 11398 19742 11450
rect 19766 11398 19776 11450
rect 19776 11398 19822 11450
rect 19526 11396 19582 11398
rect 19606 11396 19662 11398
rect 19686 11396 19742 11398
rect 19766 11396 19822 11398
rect 23240 16346 23296 16348
rect 23320 16346 23376 16348
rect 23400 16346 23456 16348
rect 23480 16346 23536 16348
rect 23240 16294 23286 16346
rect 23286 16294 23296 16346
rect 23320 16294 23350 16346
rect 23350 16294 23362 16346
rect 23362 16294 23376 16346
rect 23400 16294 23414 16346
rect 23414 16294 23426 16346
rect 23426 16294 23456 16346
rect 23480 16294 23490 16346
rect 23490 16294 23536 16346
rect 23240 16292 23296 16294
rect 23320 16292 23376 16294
rect 23400 16292 23456 16294
rect 23480 16292 23536 16294
rect 26954 28858 27010 28860
rect 27034 28858 27090 28860
rect 27114 28858 27170 28860
rect 27194 28858 27250 28860
rect 26954 28806 27000 28858
rect 27000 28806 27010 28858
rect 27034 28806 27064 28858
rect 27064 28806 27076 28858
rect 27076 28806 27090 28858
rect 27114 28806 27128 28858
rect 27128 28806 27140 28858
rect 27140 28806 27170 28858
rect 27194 28806 27204 28858
rect 27204 28806 27250 28858
rect 26954 28804 27010 28806
rect 27034 28804 27090 28806
rect 27114 28804 27170 28806
rect 27194 28804 27250 28806
rect 26954 27770 27010 27772
rect 27034 27770 27090 27772
rect 27114 27770 27170 27772
rect 27194 27770 27250 27772
rect 26954 27718 27000 27770
rect 27000 27718 27010 27770
rect 27034 27718 27064 27770
rect 27064 27718 27076 27770
rect 27076 27718 27090 27770
rect 27114 27718 27128 27770
rect 27128 27718 27140 27770
rect 27140 27718 27170 27770
rect 27194 27718 27204 27770
rect 27204 27718 27250 27770
rect 26954 27716 27010 27718
rect 27034 27716 27090 27718
rect 27114 27716 27170 27718
rect 27194 27716 27250 27718
rect 26954 26682 27010 26684
rect 27034 26682 27090 26684
rect 27114 26682 27170 26684
rect 27194 26682 27250 26684
rect 26954 26630 27000 26682
rect 27000 26630 27010 26682
rect 27034 26630 27064 26682
rect 27064 26630 27076 26682
rect 27076 26630 27090 26682
rect 27114 26630 27128 26682
rect 27128 26630 27140 26682
rect 27140 26630 27170 26682
rect 27194 26630 27204 26682
rect 27204 26630 27250 26682
rect 26954 26628 27010 26630
rect 27034 26628 27090 26630
rect 27114 26628 27170 26630
rect 27194 26628 27250 26630
rect 26954 25594 27010 25596
rect 27034 25594 27090 25596
rect 27114 25594 27170 25596
rect 27194 25594 27250 25596
rect 26954 25542 27000 25594
rect 27000 25542 27010 25594
rect 27034 25542 27064 25594
rect 27064 25542 27076 25594
rect 27076 25542 27090 25594
rect 27114 25542 27128 25594
rect 27128 25542 27140 25594
rect 27140 25542 27170 25594
rect 27194 25542 27204 25594
rect 27204 25542 27250 25594
rect 26954 25540 27010 25542
rect 27034 25540 27090 25542
rect 27114 25540 27170 25542
rect 27194 25540 27250 25542
rect 26954 24506 27010 24508
rect 27034 24506 27090 24508
rect 27114 24506 27170 24508
rect 27194 24506 27250 24508
rect 26954 24454 27000 24506
rect 27000 24454 27010 24506
rect 27034 24454 27064 24506
rect 27064 24454 27076 24506
rect 27076 24454 27090 24506
rect 27114 24454 27128 24506
rect 27128 24454 27140 24506
rect 27140 24454 27170 24506
rect 27194 24454 27204 24506
rect 27204 24454 27250 24506
rect 26954 24452 27010 24454
rect 27034 24452 27090 24454
rect 27114 24452 27170 24454
rect 27194 24452 27250 24454
rect 26954 23418 27010 23420
rect 27034 23418 27090 23420
rect 27114 23418 27170 23420
rect 27194 23418 27250 23420
rect 26954 23366 27000 23418
rect 27000 23366 27010 23418
rect 27034 23366 27064 23418
rect 27064 23366 27076 23418
rect 27076 23366 27090 23418
rect 27114 23366 27128 23418
rect 27128 23366 27140 23418
rect 27140 23366 27170 23418
rect 27194 23366 27204 23418
rect 27204 23366 27250 23418
rect 26954 23364 27010 23366
rect 27034 23364 27090 23366
rect 27114 23364 27170 23366
rect 27194 23364 27250 23366
rect 26954 22330 27010 22332
rect 27034 22330 27090 22332
rect 27114 22330 27170 22332
rect 27194 22330 27250 22332
rect 26954 22278 27000 22330
rect 27000 22278 27010 22330
rect 27034 22278 27064 22330
rect 27064 22278 27076 22330
rect 27076 22278 27090 22330
rect 27114 22278 27128 22330
rect 27128 22278 27140 22330
rect 27140 22278 27170 22330
rect 27194 22278 27204 22330
rect 27204 22278 27250 22330
rect 26954 22276 27010 22278
rect 27034 22276 27090 22278
rect 27114 22276 27170 22278
rect 27194 22276 27250 22278
rect 30668 28314 30724 28316
rect 30748 28314 30804 28316
rect 30828 28314 30884 28316
rect 30908 28314 30964 28316
rect 30668 28262 30714 28314
rect 30714 28262 30724 28314
rect 30748 28262 30778 28314
rect 30778 28262 30790 28314
rect 30790 28262 30804 28314
rect 30828 28262 30842 28314
rect 30842 28262 30854 28314
rect 30854 28262 30884 28314
rect 30908 28262 30918 28314
rect 30918 28262 30964 28314
rect 30668 28260 30724 28262
rect 30748 28260 30804 28262
rect 30828 28260 30884 28262
rect 30908 28260 30964 28262
rect 30668 27226 30724 27228
rect 30748 27226 30804 27228
rect 30828 27226 30884 27228
rect 30908 27226 30964 27228
rect 30668 27174 30714 27226
rect 30714 27174 30724 27226
rect 30748 27174 30778 27226
rect 30778 27174 30790 27226
rect 30790 27174 30804 27226
rect 30828 27174 30842 27226
rect 30842 27174 30854 27226
rect 30854 27174 30884 27226
rect 30908 27174 30918 27226
rect 30918 27174 30964 27226
rect 30668 27172 30724 27174
rect 30748 27172 30804 27174
rect 30828 27172 30884 27174
rect 30908 27172 30964 27174
rect 30668 26138 30724 26140
rect 30748 26138 30804 26140
rect 30828 26138 30884 26140
rect 30908 26138 30964 26140
rect 30668 26086 30714 26138
rect 30714 26086 30724 26138
rect 30748 26086 30778 26138
rect 30778 26086 30790 26138
rect 30790 26086 30804 26138
rect 30828 26086 30842 26138
rect 30842 26086 30854 26138
rect 30854 26086 30884 26138
rect 30908 26086 30918 26138
rect 30918 26086 30964 26138
rect 30668 26084 30724 26086
rect 30748 26084 30804 26086
rect 30828 26084 30884 26086
rect 30908 26084 30964 26086
rect 31022 25744 31078 25800
rect 26954 21242 27010 21244
rect 27034 21242 27090 21244
rect 27114 21242 27170 21244
rect 27194 21242 27250 21244
rect 26954 21190 27000 21242
rect 27000 21190 27010 21242
rect 27034 21190 27064 21242
rect 27064 21190 27076 21242
rect 27076 21190 27090 21242
rect 27114 21190 27128 21242
rect 27128 21190 27140 21242
rect 27140 21190 27170 21242
rect 27194 21190 27204 21242
rect 27204 21190 27250 21242
rect 26954 21188 27010 21190
rect 27034 21188 27090 21190
rect 27114 21188 27170 21190
rect 27194 21188 27250 21190
rect 26954 20154 27010 20156
rect 27034 20154 27090 20156
rect 27114 20154 27170 20156
rect 27194 20154 27250 20156
rect 26954 20102 27000 20154
rect 27000 20102 27010 20154
rect 27034 20102 27064 20154
rect 27064 20102 27076 20154
rect 27076 20102 27090 20154
rect 27114 20102 27128 20154
rect 27128 20102 27140 20154
rect 27140 20102 27170 20154
rect 27194 20102 27204 20154
rect 27204 20102 27250 20154
rect 26954 20100 27010 20102
rect 27034 20100 27090 20102
rect 27114 20100 27170 20102
rect 27194 20100 27250 20102
rect 26954 19066 27010 19068
rect 27034 19066 27090 19068
rect 27114 19066 27170 19068
rect 27194 19066 27250 19068
rect 26954 19014 27000 19066
rect 27000 19014 27010 19066
rect 27034 19014 27064 19066
rect 27064 19014 27076 19066
rect 27076 19014 27090 19066
rect 27114 19014 27128 19066
rect 27128 19014 27140 19066
rect 27140 19014 27170 19066
rect 27194 19014 27204 19066
rect 27204 19014 27250 19066
rect 26954 19012 27010 19014
rect 27034 19012 27090 19014
rect 27114 19012 27170 19014
rect 27194 19012 27250 19014
rect 30668 25050 30724 25052
rect 30748 25050 30804 25052
rect 30828 25050 30884 25052
rect 30908 25050 30964 25052
rect 30668 24998 30714 25050
rect 30714 24998 30724 25050
rect 30748 24998 30778 25050
rect 30778 24998 30790 25050
rect 30790 24998 30804 25050
rect 30828 24998 30842 25050
rect 30842 24998 30854 25050
rect 30854 24998 30884 25050
rect 30908 24998 30918 25050
rect 30918 24998 30964 25050
rect 30668 24996 30724 24998
rect 30748 24996 30804 24998
rect 30828 24996 30884 24998
rect 30908 24996 30964 24998
rect 30668 23962 30724 23964
rect 30748 23962 30804 23964
rect 30828 23962 30884 23964
rect 30908 23962 30964 23964
rect 30668 23910 30714 23962
rect 30714 23910 30724 23962
rect 30748 23910 30778 23962
rect 30778 23910 30790 23962
rect 30790 23910 30804 23962
rect 30828 23910 30842 23962
rect 30842 23910 30854 23962
rect 30854 23910 30884 23962
rect 30908 23910 30918 23962
rect 30918 23910 30964 23962
rect 30668 23908 30724 23910
rect 30748 23908 30804 23910
rect 30828 23908 30884 23910
rect 30908 23908 30964 23910
rect 30668 22874 30724 22876
rect 30748 22874 30804 22876
rect 30828 22874 30884 22876
rect 30908 22874 30964 22876
rect 30668 22822 30714 22874
rect 30714 22822 30724 22874
rect 30748 22822 30778 22874
rect 30778 22822 30790 22874
rect 30790 22822 30804 22874
rect 30828 22822 30842 22874
rect 30842 22822 30854 22874
rect 30854 22822 30884 22874
rect 30908 22822 30918 22874
rect 30918 22822 30964 22874
rect 30668 22820 30724 22822
rect 30748 22820 30804 22822
rect 30828 22820 30884 22822
rect 30908 22820 30964 22822
rect 31022 21956 31078 21992
rect 31022 21936 31024 21956
rect 31024 21936 31076 21956
rect 31076 21936 31078 21956
rect 30668 21786 30724 21788
rect 30748 21786 30804 21788
rect 30828 21786 30884 21788
rect 30908 21786 30964 21788
rect 30668 21734 30714 21786
rect 30714 21734 30724 21786
rect 30748 21734 30778 21786
rect 30778 21734 30790 21786
rect 30790 21734 30804 21786
rect 30828 21734 30842 21786
rect 30842 21734 30854 21786
rect 30854 21734 30884 21786
rect 30908 21734 30918 21786
rect 30918 21734 30964 21786
rect 30668 21732 30724 21734
rect 30748 21732 30804 21734
rect 30828 21732 30884 21734
rect 30908 21732 30964 21734
rect 30668 20698 30724 20700
rect 30748 20698 30804 20700
rect 30828 20698 30884 20700
rect 30908 20698 30964 20700
rect 30668 20646 30714 20698
rect 30714 20646 30724 20698
rect 30748 20646 30778 20698
rect 30778 20646 30790 20698
rect 30790 20646 30804 20698
rect 30828 20646 30842 20698
rect 30842 20646 30854 20698
rect 30854 20646 30884 20698
rect 30908 20646 30918 20698
rect 30918 20646 30964 20698
rect 30668 20644 30724 20646
rect 30748 20644 30804 20646
rect 30828 20644 30884 20646
rect 30908 20644 30964 20646
rect 30668 19610 30724 19612
rect 30748 19610 30804 19612
rect 30828 19610 30884 19612
rect 30908 19610 30964 19612
rect 30668 19558 30714 19610
rect 30714 19558 30724 19610
rect 30748 19558 30778 19610
rect 30778 19558 30790 19610
rect 30790 19558 30804 19610
rect 30828 19558 30842 19610
rect 30842 19558 30854 19610
rect 30854 19558 30884 19610
rect 30908 19558 30918 19610
rect 30918 19558 30964 19610
rect 30668 19556 30724 19558
rect 30748 19556 30804 19558
rect 30828 19556 30884 19558
rect 30908 19556 30964 19558
rect 23240 15258 23296 15260
rect 23320 15258 23376 15260
rect 23400 15258 23456 15260
rect 23480 15258 23536 15260
rect 23240 15206 23286 15258
rect 23286 15206 23296 15258
rect 23320 15206 23350 15258
rect 23350 15206 23362 15258
rect 23362 15206 23376 15258
rect 23400 15206 23414 15258
rect 23414 15206 23426 15258
rect 23426 15206 23456 15258
rect 23480 15206 23490 15258
rect 23490 15206 23536 15258
rect 23240 15204 23296 15206
rect 23320 15204 23376 15206
rect 23400 15204 23456 15206
rect 23480 15204 23536 15206
rect 23240 14170 23296 14172
rect 23320 14170 23376 14172
rect 23400 14170 23456 14172
rect 23480 14170 23536 14172
rect 23240 14118 23286 14170
rect 23286 14118 23296 14170
rect 23320 14118 23350 14170
rect 23350 14118 23362 14170
rect 23362 14118 23376 14170
rect 23400 14118 23414 14170
rect 23414 14118 23426 14170
rect 23426 14118 23456 14170
rect 23480 14118 23490 14170
rect 23490 14118 23536 14170
rect 23240 14116 23296 14118
rect 23320 14116 23376 14118
rect 23400 14116 23456 14118
rect 23480 14116 23536 14118
rect 23240 13082 23296 13084
rect 23320 13082 23376 13084
rect 23400 13082 23456 13084
rect 23480 13082 23536 13084
rect 23240 13030 23286 13082
rect 23286 13030 23296 13082
rect 23320 13030 23350 13082
rect 23350 13030 23362 13082
rect 23362 13030 23376 13082
rect 23400 13030 23414 13082
rect 23414 13030 23426 13082
rect 23426 13030 23456 13082
rect 23480 13030 23490 13082
rect 23490 13030 23536 13082
rect 23240 13028 23296 13030
rect 23320 13028 23376 13030
rect 23400 13028 23456 13030
rect 23480 13028 23536 13030
rect 19526 10362 19582 10364
rect 19606 10362 19662 10364
rect 19686 10362 19742 10364
rect 19766 10362 19822 10364
rect 19526 10310 19572 10362
rect 19572 10310 19582 10362
rect 19606 10310 19636 10362
rect 19636 10310 19648 10362
rect 19648 10310 19662 10362
rect 19686 10310 19700 10362
rect 19700 10310 19712 10362
rect 19712 10310 19742 10362
rect 19766 10310 19776 10362
rect 19776 10310 19822 10362
rect 19526 10308 19582 10310
rect 19606 10308 19662 10310
rect 19686 10308 19742 10310
rect 19766 10308 19822 10310
rect 23240 11994 23296 11996
rect 23320 11994 23376 11996
rect 23400 11994 23456 11996
rect 23480 11994 23536 11996
rect 23240 11942 23286 11994
rect 23286 11942 23296 11994
rect 23320 11942 23350 11994
rect 23350 11942 23362 11994
rect 23362 11942 23376 11994
rect 23400 11942 23414 11994
rect 23414 11942 23426 11994
rect 23426 11942 23456 11994
rect 23480 11942 23490 11994
rect 23490 11942 23536 11994
rect 23240 11940 23296 11942
rect 23320 11940 23376 11942
rect 23400 11940 23456 11942
rect 23480 11940 23536 11942
rect 23240 10906 23296 10908
rect 23320 10906 23376 10908
rect 23400 10906 23456 10908
rect 23480 10906 23536 10908
rect 23240 10854 23286 10906
rect 23286 10854 23296 10906
rect 23320 10854 23350 10906
rect 23350 10854 23362 10906
rect 23362 10854 23376 10906
rect 23400 10854 23414 10906
rect 23414 10854 23426 10906
rect 23426 10854 23456 10906
rect 23480 10854 23490 10906
rect 23490 10854 23536 10906
rect 23240 10852 23296 10854
rect 23320 10852 23376 10854
rect 23400 10852 23456 10854
rect 23480 10852 23536 10854
rect 23240 9818 23296 9820
rect 23320 9818 23376 9820
rect 23400 9818 23456 9820
rect 23480 9818 23536 9820
rect 23240 9766 23286 9818
rect 23286 9766 23296 9818
rect 23320 9766 23350 9818
rect 23350 9766 23362 9818
rect 23362 9766 23376 9818
rect 23400 9766 23414 9818
rect 23414 9766 23426 9818
rect 23426 9766 23456 9818
rect 23480 9766 23490 9818
rect 23490 9766 23536 9818
rect 23240 9764 23296 9766
rect 23320 9764 23376 9766
rect 23400 9764 23456 9766
rect 23480 9764 23536 9766
rect 19526 9274 19582 9276
rect 19606 9274 19662 9276
rect 19686 9274 19742 9276
rect 19766 9274 19822 9276
rect 19526 9222 19572 9274
rect 19572 9222 19582 9274
rect 19606 9222 19636 9274
rect 19636 9222 19648 9274
rect 19648 9222 19662 9274
rect 19686 9222 19700 9274
rect 19700 9222 19712 9274
rect 19712 9222 19742 9274
rect 19766 9222 19776 9274
rect 19776 9222 19822 9274
rect 19526 9220 19582 9222
rect 19606 9220 19662 9222
rect 19686 9220 19742 9222
rect 19766 9220 19822 9222
rect 26954 17978 27010 17980
rect 27034 17978 27090 17980
rect 27114 17978 27170 17980
rect 27194 17978 27250 17980
rect 26954 17926 27000 17978
rect 27000 17926 27010 17978
rect 27034 17926 27064 17978
rect 27064 17926 27076 17978
rect 27076 17926 27090 17978
rect 27114 17926 27128 17978
rect 27128 17926 27140 17978
rect 27140 17926 27170 17978
rect 27194 17926 27204 17978
rect 27204 17926 27250 17978
rect 26954 17924 27010 17926
rect 27034 17924 27090 17926
rect 27114 17924 27170 17926
rect 27194 17924 27250 17926
rect 26954 16890 27010 16892
rect 27034 16890 27090 16892
rect 27114 16890 27170 16892
rect 27194 16890 27250 16892
rect 26954 16838 27000 16890
rect 27000 16838 27010 16890
rect 27034 16838 27064 16890
rect 27064 16838 27076 16890
rect 27076 16838 27090 16890
rect 27114 16838 27128 16890
rect 27128 16838 27140 16890
rect 27140 16838 27170 16890
rect 27194 16838 27204 16890
rect 27204 16838 27250 16890
rect 26954 16836 27010 16838
rect 27034 16836 27090 16838
rect 27114 16836 27170 16838
rect 27194 16836 27250 16838
rect 26954 15802 27010 15804
rect 27034 15802 27090 15804
rect 27114 15802 27170 15804
rect 27194 15802 27250 15804
rect 26954 15750 27000 15802
rect 27000 15750 27010 15802
rect 27034 15750 27064 15802
rect 27064 15750 27076 15802
rect 27076 15750 27090 15802
rect 27114 15750 27128 15802
rect 27128 15750 27140 15802
rect 27140 15750 27170 15802
rect 27194 15750 27204 15802
rect 27204 15750 27250 15802
rect 26954 15748 27010 15750
rect 27034 15748 27090 15750
rect 27114 15748 27170 15750
rect 27194 15748 27250 15750
rect 26954 14714 27010 14716
rect 27034 14714 27090 14716
rect 27114 14714 27170 14716
rect 27194 14714 27250 14716
rect 26954 14662 27000 14714
rect 27000 14662 27010 14714
rect 27034 14662 27064 14714
rect 27064 14662 27076 14714
rect 27076 14662 27090 14714
rect 27114 14662 27128 14714
rect 27128 14662 27140 14714
rect 27140 14662 27170 14714
rect 27194 14662 27204 14714
rect 27204 14662 27250 14714
rect 26954 14660 27010 14662
rect 27034 14660 27090 14662
rect 27114 14660 27170 14662
rect 27194 14660 27250 14662
rect 26954 13626 27010 13628
rect 27034 13626 27090 13628
rect 27114 13626 27170 13628
rect 27194 13626 27250 13628
rect 26954 13574 27000 13626
rect 27000 13574 27010 13626
rect 27034 13574 27064 13626
rect 27064 13574 27076 13626
rect 27076 13574 27090 13626
rect 27114 13574 27128 13626
rect 27128 13574 27140 13626
rect 27140 13574 27170 13626
rect 27194 13574 27204 13626
rect 27204 13574 27250 13626
rect 26954 13572 27010 13574
rect 27034 13572 27090 13574
rect 27114 13572 27170 13574
rect 27194 13572 27250 13574
rect 26954 12538 27010 12540
rect 27034 12538 27090 12540
rect 27114 12538 27170 12540
rect 27194 12538 27250 12540
rect 26954 12486 27000 12538
rect 27000 12486 27010 12538
rect 27034 12486 27064 12538
rect 27064 12486 27076 12538
rect 27076 12486 27090 12538
rect 27114 12486 27128 12538
rect 27128 12486 27140 12538
rect 27140 12486 27170 12538
rect 27194 12486 27204 12538
rect 27204 12486 27250 12538
rect 26954 12484 27010 12486
rect 27034 12484 27090 12486
rect 27114 12484 27170 12486
rect 27194 12484 27250 12486
rect 26954 11450 27010 11452
rect 27034 11450 27090 11452
rect 27114 11450 27170 11452
rect 27194 11450 27250 11452
rect 26954 11398 27000 11450
rect 27000 11398 27010 11450
rect 27034 11398 27064 11450
rect 27064 11398 27076 11450
rect 27076 11398 27090 11450
rect 27114 11398 27128 11450
rect 27128 11398 27140 11450
rect 27140 11398 27170 11450
rect 27194 11398 27204 11450
rect 27204 11398 27250 11450
rect 26954 11396 27010 11398
rect 27034 11396 27090 11398
rect 27114 11396 27170 11398
rect 27194 11396 27250 11398
rect 26954 10362 27010 10364
rect 27034 10362 27090 10364
rect 27114 10362 27170 10364
rect 27194 10362 27250 10364
rect 26954 10310 27000 10362
rect 27000 10310 27010 10362
rect 27034 10310 27064 10362
rect 27064 10310 27076 10362
rect 27076 10310 27090 10362
rect 27114 10310 27128 10362
rect 27128 10310 27140 10362
rect 27140 10310 27170 10362
rect 27194 10310 27204 10362
rect 27204 10310 27250 10362
rect 26954 10308 27010 10310
rect 27034 10308 27090 10310
rect 27114 10308 27170 10310
rect 27194 10308 27250 10310
rect 30668 18522 30724 18524
rect 30748 18522 30804 18524
rect 30828 18522 30884 18524
rect 30908 18522 30964 18524
rect 30668 18470 30714 18522
rect 30714 18470 30724 18522
rect 30748 18470 30778 18522
rect 30778 18470 30790 18522
rect 30790 18470 30804 18522
rect 30828 18470 30842 18522
rect 30842 18470 30854 18522
rect 30854 18470 30884 18522
rect 30908 18470 30918 18522
rect 30918 18470 30964 18522
rect 30668 18468 30724 18470
rect 30748 18468 30804 18470
rect 30828 18468 30884 18470
rect 30908 18468 30964 18470
rect 31022 17856 31078 17912
rect 30668 17434 30724 17436
rect 30748 17434 30804 17436
rect 30828 17434 30884 17436
rect 30908 17434 30964 17436
rect 30668 17382 30714 17434
rect 30714 17382 30724 17434
rect 30748 17382 30778 17434
rect 30778 17382 30790 17434
rect 30790 17382 30804 17434
rect 30828 17382 30842 17434
rect 30842 17382 30854 17434
rect 30854 17382 30884 17434
rect 30908 17382 30918 17434
rect 30918 17382 30964 17434
rect 30668 17380 30724 17382
rect 30748 17380 30804 17382
rect 30828 17380 30884 17382
rect 30908 17380 30964 17382
rect 30668 16346 30724 16348
rect 30748 16346 30804 16348
rect 30828 16346 30884 16348
rect 30908 16346 30964 16348
rect 30668 16294 30714 16346
rect 30714 16294 30724 16346
rect 30748 16294 30778 16346
rect 30778 16294 30790 16346
rect 30790 16294 30804 16346
rect 30828 16294 30842 16346
rect 30842 16294 30854 16346
rect 30854 16294 30884 16346
rect 30908 16294 30918 16346
rect 30918 16294 30964 16346
rect 30668 16292 30724 16294
rect 30748 16292 30804 16294
rect 30828 16292 30884 16294
rect 30908 16292 30964 16294
rect 30668 15258 30724 15260
rect 30748 15258 30804 15260
rect 30828 15258 30884 15260
rect 30908 15258 30964 15260
rect 30668 15206 30714 15258
rect 30714 15206 30724 15258
rect 30748 15206 30778 15258
rect 30778 15206 30790 15258
rect 30790 15206 30804 15258
rect 30828 15206 30842 15258
rect 30842 15206 30854 15258
rect 30854 15206 30884 15258
rect 30908 15206 30918 15258
rect 30918 15206 30964 15258
rect 30668 15204 30724 15206
rect 30748 15204 30804 15206
rect 30828 15204 30884 15206
rect 30908 15204 30964 15206
rect 30668 14170 30724 14172
rect 30748 14170 30804 14172
rect 30828 14170 30884 14172
rect 30908 14170 30964 14172
rect 30668 14118 30714 14170
rect 30714 14118 30724 14170
rect 30748 14118 30778 14170
rect 30778 14118 30790 14170
rect 30790 14118 30804 14170
rect 30828 14118 30842 14170
rect 30842 14118 30854 14170
rect 30854 14118 30884 14170
rect 30908 14118 30918 14170
rect 30918 14118 30964 14170
rect 30668 14116 30724 14118
rect 30748 14116 30804 14118
rect 30828 14116 30884 14118
rect 30908 14116 30964 14118
rect 31022 13912 31078 13968
rect 30668 13082 30724 13084
rect 30748 13082 30804 13084
rect 30828 13082 30884 13084
rect 30908 13082 30964 13084
rect 30668 13030 30714 13082
rect 30714 13030 30724 13082
rect 30748 13030 30778 13082
rect 30778 13030 30790 13082
rect 30790 13030 30804 13082
rect 30828 13030 30842 13082
rect 30842 13030 30854 13082
rect 30854 13030 30884 13082
rect 30908 13030 30918 13082
rect 30918 13030 30964 13082
rect 30668 13028 30724 13030
rect 30748 13028 30804 13030
rect 30828 13028 30884 13030
rect 30908 13028 30964 13030
rect 30668 11994 30724 11996
rect 30748 11994 30804 11996
rect 30828 11994 30884 11996
rect 30908 11994 30964 11996
rect 30668 11942 30714 11994
rect 30714 11942 30724 11994
rect 30748 11942 30778 11994
rect 30778 11942 30790 11994
rect 30790 11942 30804 11994
rect 30828 11942 30842 11994
rect 30842 11942 30854 11994
rect 30854 11942 30884 11994
rect 30908 11942 30918 11994
rect 30918 11942 30964 11994
rect 30668 11940 30724 11942
rect 30748 11940 30804 11942
rect 30828 11940 30884 11942
rect 30908 11940 30964 11942
rect 30668 10906 30724 10908
rect 30748 10906 30804 10908
rect 30828 10906 30884 10908
rect 30908 10906 30964 10908
rect 30668 10854 30714 10906
rect 30714 10854 30724 10906
rect 30748 10854 30778 10906
rect 30778 10854 30790 10906
rect 30790 10854 30804 10906
rect 30828 10854 30842 10906
rect 30842 10854 30854 10906
rect 30854 10854 30884 10906
rect 30908 10854 30918 10906
rect 30918 10854 30964 10906
rect 30668 10852 30724 10854
rect 30748 10852 30804 10854
rect 30828 10852 30884 10854
rect 30908 10852 30964 10854
rect 26954 9274 27010 9276
rect 27034 9274 27090 9276
rect 27114 9274 27170 9276
rect 27194 9274 27250 9276
rect 26954 9222 27000 9274
rect 27000 9222 27010 9274
rect 27034 9222 27064 9274
rect 27064 9222 27076 9274
rect 27076 9222 27090 9274
rect 27114 9222 27128 9274
rect 27128 9222 27140 9274
rect 27140 9222 27170 9274
rect 27194 9222 27204 9274
rect 27204 9222 27250 9274
rect 26954 9220 27010 9222
rect 27034 9220 27090 9222
rect 27114 9220 27170 9222
rect 27194 9220 27250 9222
rect 19526 8186 19582 8188
rect 19606 8186 19662 8188
rect 19686 8186 19742 8188
rect 19766 8186 19822 8188
rect 19526 8134 19572 8186
rect 19572 8134 19582 8186
rect 19606 8134 19636 8186
rect 19636 8134 19648 8186
rect 19648 8134 19662 8186
rect 19686 8134 19700 8186
rect 19700 8134 19712 8186
rect 19712 8134 19742 8186
rect 19766 8134 19776 8186
rect 19776 8134 19822 8186
rect 19526 8132 19582 8134
rect 19606 8132 19662 8134
rect 19686 8132 19742 8134
rect 19766 8132 19822 8134
rect 15812 6554 15868 6556
rect 15892 6554 15948 6556
rect 15972 6554 16028 6556
rect 16052 6554 16108 6556
rect 15812 6502 15858 6554
rect 15858 6502 15868 6554
rect 15892 6502 15922 6554
rect 15922 6502 15934 6554
rect 15934 6502 15948 6554
rect 15972 6502 15986 6554
rect 15986 6502 15998 6554
rect 15998 6502 16028 6554
rect 16052 6502 16062 6554
rect 16062 6502 16108 6554
rect 15812 6500 15868 6502
rect 15892 6500 15948 6502
rect 15972 6500 16028 6502
rect 16052 6500 16108 6502
rect 15812 5466 15868 5468
rect 15892 5466 15948 5468
rect 15972 5466 16028 5468
rect 16052 5466 16108 5468
rect 15812 5414 15858 5466
rect 15858 5414 15868 5466
rect 15892 5414 15922 5466
rect 15922 5414 15934 5466
rect 15934 5414 15948 5466
rect 15972 5414 15986 5466
rect 15986 5414 15998 5466
rect 15998 5414 16028 5466
rect 16052 5414 16062 5466
rect 16062 5414 16108 5466
rect 15812 5412 15868 5414
rect 15892 5412 15948 5414
rect 15972 5412 16028 5414
rect 16052 5412 16108 5414
rect 4670 4922 4726 4924
rect 4750 4922 4806 4924
rect 4830 4922 4886 4924
rect 4910 4922 4966 4924
rect 4670 4870 4716 4922
rect 4716 4870 4726 4922
rect 4750 4870 4780 4922
rect 4780 4870 4792 4922
rect 4792 4870 4806 4922
rect 4830 4870 4844 4922
rect 4844 4870 4856 4922
rect 4856 4870 4886 4922
rect 4910 4870 4920 4922
rect 4920 4870 4966 4922
rect 4670 4868 4726 4870
rect 4750 4868 4806 4870
rect 4830 4868 4886 4870
rect 4910 4868 4966 4870
rect 12098 4922 12154 4924
rect 12178 4922 12234 4924
rect 12258 4922 12314 4924
rect 12338 4922 12394 4924
rect 12098 4870 12144 4922
rect 12144 4870 12154 4922
rect 12178 4870 12208 4922
rect 12208 4870 12220 4922
rect 12220 4870 12234 4922
rect 12258 4870 12272 4922
rect 12272 4870 12284 4922
rect 12284 4870 12314 4922
rect 12338 4870 12348 4922
rect 12348 4870 12394 4922
rect 12098 4868 12154 4870
rect 12178 4868 12234 4870
rect 12258 4868 12314 4870
rect 12338 4868 12394 4870
rect 8384 4378 8440 4380
rect 8464 4378 8520 4380
rect 8544 4378 8600 4380
rect 8624 4378 8680 4380
rect 8384 4326 8430 4378
rect 8430 4326 8440 4378
rect 8464 4326 8494 4378
rect 8494 4326 8506 4378
rect 8506 4326 8520 4378
rect 8544 4326 8558 4378
rect 8558 4326 8570 4378
rect 8570 4326 8600 4378
rect 8624 4326 8634 4378
rect 8634 4326 8680 4378
rect 8384 4324 8440 4326
rect 8464 4324 8520 4326
rect 8544 4324 8600 4326
rect 8624 4324 8680 4326
rect 23240 8730 23296 8732
rect 23320 8730 23376 8732
rect 23400 8730 23456 8732
rect 23480 8730 23536 8732
rect 23240 8678 23286 8730
rect 23286 8678 23296 8730
rect 23320 8678 23350 8730
rect 23350 8678 23362 8730
rect 23362 8678 23376 8730
rect 23400 8678 23414 8730
rect 23414 8678 23426 8730
rect 23426 8678 23456 8730
rect 23480 8678 23490 8730
rect 23490 8678 23536 8730
rect 23240 8676 23296 8678
rect 23320 8676 23376 8678
rect 23400 8676 23456 8678
rect 23480 8676 23536 8678
rect 19526 7098 19582 7100
rect 19606 7098 19662 7100
rect 19686 7098 19742 7100
rect 19766 7098 19822 7100
rect 19526 7046 19572 7098
rect 19572 7046 19582 7098
rect 19606 7046 19636 7098
rect 19636 7046 19648 7098
rect 19648 7046 19662 7098
rect 19686 7046 19700 7098
rect 19700 7046 19712 7098
rect 19712 7046 19742 7098
rect 19766 7046 19776 7098
rect 19776 7046 19822 7098
rect 19526 7044 19582 7046
rect 19606 7044 19662 7046
rect 19686 7044 19742 7046
rect 19766 7044 19822 7046
rect 19526 6010 19582 6012
rect 19606 6010 19662 6012
rect 19686 6010 19742 6012
rect 19766 6010 19822 6012
rect 19526 5958 19572 6010
rect 19572 5958 19582 6010
rect 19606 5958 19636 6010
rect 19636 5958 19648 6010
rect 19648 5958 19662 6010
rect 19686 5958 19700 6010
rect 19700 5958 19712 6010
rect 19712 5958 19742 6010
rect 19766 5958 19776 6010
rect 19776 5958 19822 6010
rect 19526 5956 19582 5958
rect 19606 5956 19662 5958
rect 19686 5956 19742 5958
rect 19766 5956 19822 5958
rect 26954 8186 27010 8188
rect 27034 8186 27090 8188
rect 27114 8186 27170 8188
rect 27194 8186 27250 8188
rect 26954 8134 27000 8186
rect 27000 8134 27010 8186
rect 27034 8134 27064 8186
rect 27064 8134 27076 8186
rect 27076 8134 27090 8186
rect 27114 8134 27128 8186
rect 27128 8134 27140 8186
rect 27140 8134 27170 8186
rect 27194 8134 27204 8186
rect 27204 8134 27250 8186
rect 26954 8132 27010 8134
rect 27034 8132 27090 8134
rect 27114 8132 27170 8134
rect 27194 8132 27250 8134
rect 23240 7642 23296 7644
rect 23320 7642 23376 7644
rect 23400 7642 23456 7644
rect 23480 7642 23536 7644
rect 23240 7590 23286 7642
rect 23286 7590 23296 7642
rect 23320 7590 23350 7642
rect 23350 7590 23362 7642
rect 23362 7590 23376 7642
rect 23400 7590 23414 7642
rect 23414 7590 23426 7642
rect 23426 7590 23456 7642
rect 23480 7590 23490 7642
rect 23490 7590 23536 7642
rect 23240 7588 23296 7590
rect 23320 7588 23376 7590
rect 23400 7588 23456 7590
rect 23480 7588 23536 7590
rect 19526 4922 19582 4924
rect 19606 4922 19662 4924
rect 19686 4922 19742 4924
rect 19766 4922 19822 4924
rect 19526 4870 19572 4922
rect 19572 4870 19582 4922
rect 19606 4870 19636 4922
rect 19636 4870 19648 4922
rect 19648 4870 19662 4922
rect 19686 4870 19700 4922
rect 19700 4870 19712 4922
rect 19712 4870 19742 4922
rect 19766 4870 19776 4922
rect 19776 4870 19822 4922
rect 19526 4868 19582 4870
rect 19606 4868 19662 4870
rect 19686 4868 19742 4870
rect 19766 4868 19822 4870
rect 23240 6554 23296 6556
rect 23320 6554 23376 6556
rect 23400 6554 23456 6556
rect 23480 6554 23536 6556
rect 23240 6502 23286 6554
rect 23286 6502 23296 6554
rect 23320 6502 23350 6554
rect 23350 6502 23362 6554
rect 23362 6502 23376 6554
rect 23400 6502 23414 6554
rect 23414 6502 23426 6554
rect 23426 6502 23456 6554
rect 23480 6502 23490 6554
rect 23490 6502 23536 6554
rect 23240 6500 23296 6502
rect 23320 6500 23376 6502
rect 23400 6500 23456 6502
rect 23480 6500 23536 6502
rect 26954 7098 27010 7100
rect 27034 7098 27090 7100
rect 27114 7098 27170 7100
rect 27194 7098 27250 7100
rect 26954 7046 27000 7098
rect 27000 7046 27010 7098
rect 27034 7046 27064 7098
rect 27064 7046 27076 7098
rect 27076 7046 27090 7098
rect 27114 7046 27128 7098
rect 27128 7046 27140 7098
rect 27140 7046 27170 7098
rect 27194 7046 27204 7098
rect 27204 7046 27250 7098
rect 26954 7044 27010 7046
rect 27034 7044 27090 7046
rect 27114 7044 27170 7046
rect 27194 7044 27250 7046
rect 26954 6010 27010 6012
rect 27034 6010 27090 6012
rect 27114 6010 27170 6012
rect 27194 6010 27250 6012
rect 26954 5958 27000 6010
rect 27000 5958 27010 6010
rect 27034 5958 27064 6010
rect 27064 5958 27076 6010
rect 27076 5958 27090 6010
rect 27114 5958 27128 6010
rect 27128 5958 27140 6010
rect 27140 5958 27170 6010
rect 27194 5958 27204 6010
rect 27204 5958 27250 6010
rect 26954 5956 27010 5958
rect 27034 5956 27090 5958
rect 27114 5956 27170 5958
rect 27194 5956 27250 5958
rect 31022 9968 31078 10024
rect 30668 9818 30724 9820
rect 30748 9818 30804 9820
rect 30828 9818 30884 9820
rect 30908 9818 30964 9820
rect 30668 9766 30714 9818
rect 30714 9766 30724 9818
rect 30748 9766 30778 9818
rect 30778 9766 30790 9818
rect 30790 9766 30804 9818
rect 30828 9766 30842 9818
rect 30842 9766 30854 9818
rect 30854 9766 30884 9818
rect 30908 9766 30918 9818
rect 30918 9766 30964 9818
rect 30668 9764 30724 9766
rect 30748 9764 30804 9766
rect 30828 9764 30884 9766
rect 30908 9764 30964 9766
rect 30668 8730 30724 8732
rect 30748 8730 30804 8732
rect 30828 8730 30884 8732
rect 30908 8730 30964 8732
rect 30668 8678 30714 8730
rect 30714 8678 30724 8730
rect 30748 8678 30778 8730
rect 30778 8678 30790 8730
rect 30790 8678 30804 8730
rect 30828 8678 30842 8730
rect 30842 8678 30854 8730
rect 30854 8678 30884 8730
rect 30908 8678 30918 8730
rect 30918 8678 30964 8730
rect 30668 8676 30724 8678
rect 30748 8676 30804 8678
rect 30828 8676 30884 8678
rect 30908 8676 30964 8678
rect 30668 7642 30724 7644
rect 30748 7642 30804 7644
rect 30828 7642 30884 7644
rect 30908 7642 30964 7644
rect 30668 7590 30714 7642
rect 30714 7590 30724 7642
rect 30748 7590 30778 7642
rect 30778 7590 30790 7642
rect 30790 7590 30804 7642
rect 30828 7590 30842 7642
rect 30842 7590 30854 7642
rect 30854 7590 30884 7642
rect 30908 7590 30918 7642
rect 30918 7590 30964 7642
rect 30668 7588 30724 7590
rect 30748 7588 30804 7590
rect 30828 7588 30884 7590
rect 30908 7588 30964 7590
rect 23240 5466 23296 5468
rect 23320 5466 23376 5468
rect 23400 5466 23456 5468
rect 23480 5466 23536 5468
rect 23240 5414 23286 5466
rect 23286 5414 23296 5466
rect 23320 5414 23350 5466
rect 23350 5414 23362 5466
rect 23362 5414 23376 5466
rect 23400 5414 23414 5466
rect 23414 5414 23426 5466
rect 23426 5414 23456 5466
rect 23480 5414 23490 5466
rect 23490 5414 23536 5466
rect 23240 5412 23296 5414
rect 23320 5412 23376 5414
rect 23400 5412 23456 5414
rect 23480 5412 23536 5414
rect 30668 6554 30724 6556
rect 30748 6554 30804 6556
rect 30828 6554 30884 6556
rect 30908 6554 30964 6556
rect 30668 6502 30714 6554
rect 30714 6502 30724 6554
rect 30748 6502 30778 6554
rect 30778 6502 30790 6554
rect 30790 6502 30804 6554
rect 30828 6502 30842 6554
rect 30842 6502 30854 6554
rect 30854 6502 30884 6554
rect 30908 6502 30918 6554
rect 30918 6502 30964 6554
rect 30668 6500 30724 6502
rect 30748 6500 30804 6502
rect 30828 6500 30884 6502
rect 30908 6500 30964 6502
rect 31022 6024 31078 6080
rect 30668 5466 30724 5468
rect 30748 5466 30804 5468
rect 30828 5466 30884 5468
rect 30908 5466 30964 5468
rect 30668 5414 30714 5466
rect 30714 5414 30724 5466
rect 30748 5414 30778 5466
rect 30778 5414 30790 5466
rect 30790 5414 30804 5466
rect 30828 5414 30842 5466
rect 30842 5414 30854 5466
rect 30854 5414 30884 5466
rect 30908 5414 30918 5466
rect 30918 5414 30964 5466
rect 30668 5412 30724 5414
rect 30748 5412 30804 5414
rect 30828 5412 30884 5414
rect 30908 5412 30964 5414
rect 26954 4922 27010 4924
rect 27034 4922 27090 4924
rect 27114 4922 27170 4924
rect 27194 4922 27250 4924
rect 26954 4870 27000 4922
rect 27000 4870 27010 4922
rect 27034 4870 27064 4922
rect 27064 4870 27076 4922
rect 27076 4870 27090 4922
rect 27114 4870 27128 4922
rect 27128 4870 27140 4922
rect 27140 4870 27170 4922
rect 27194 4870 27204 4922
rect 27204 4870 27250 4922
rect 26954 4868 27010 4870
rect 27034 4868 27090 4870
rect 27114 4868 27170 4870
rect 27194 4868 27250 4870
rect 15812 4378 15868 4380
rect 15892 4378 15948 4380
rect 15972 4378 16028 4380
rect 16052 4378 16108 4380
rect 15812 4326 15858 4378
rect 15858 4326 15868 4378
rect 15892 4326 15922 4378
rect 15922 4326 15934 4378
rect 15934 4326 15948 4378
rect 15972 4326 15986 4378
rect 15986 4326 15998 4378
rect 15998 4326 16028 4378
rect 16052 4326 16062 4378
rect 16062 4326 16108 4378
rect 15812 4324 15868 4326
rect 15892 4324 15948 4326
rect 15972 4324 16028 4326
rect 16052 4324 16108 4326
rect 23240 4378 23296 4380
rect 23320 4378 23376 4380
rect 23400 4378 23456 4380
rect 23480 4378 23536 4380
rect 23240 4326 23286 4378
rect 23286 4326 23296 4378
rect 23320 4326 23350 4378
rect 23350 4326 23362 4378
rect 23362 4326 23376 4378
rect 23400 4326 23414 4378
rect 23414 4326 23426 4378
rect 23426 4326 23456 4378
rect 23480 4326 23490 4378
rect 23490 4326 23536 4378
rect 23240 4324 23296 4326
rect 23320 4324 23376 4326
rect 23400 4324 23456 4326
rect 23480 4324 23536 4326
rect 4670 3834 4726 3836
rect 4750 3834 4806 3836
rect 4830 3834 4886 3836
rect 4910 3834 4966 3836
rect 4670 3782 4716 3834
rect 4716 3782 4726 3834
rect 4750 3782 4780 3834
rect 4780 3782 4792 3834
rect 4792 3782 4806 3834
rect 4830 3782 4844 3834
rect 4844 3782 4856 3834
rect 4856 3782 4886 3834
rect 4910 3782 4920 3834
rect 4920 3782 4966 3834
rect 4670 3780 4726 3782
rect 4750 3780 4806 3782
rect 4830 3780 4886 3782
rect 4910 3780 4966 3782
rect 12098 3834 12154 3836
rect 12178 3834 12234 3836
rect 12258 3834 12314 3836
rect 12338 3834 12394 3836
rect 12098 3782 12144 3834
rect 12144 3782 12154 3834
rect 12178 3782 12208 3834
rect 12208 3782 12220 3834
rect 12220 3782 12234 3834
rect 12258 3782 12272 3834
rect 12272 3782 12284 3834
rect 12284 3782 12314 3834
rect 12338 3782 12348 3834
rect 12348 3782 12394 3834
rect 12098 3780 12154 3782
rect 12178 3780 12234 3782
rect 12258 3780 12314 3782
rect 12338 3780 12394 3782
rect 19526 3834 19582 3836
rect 19606 3834 19662 3836
rect 19686 3834 19742 3836
rect 19766 3834 19822 3836
rect 19526 3782 19572 3834
rect 19572 3782 19582 3834
rect 19606 3782 19636 3834
rect 19636 3782 19648 3834
rect 19648 3782 19662 3834
rect 19686 3782 19700 3834
rect 19700 3782 19712 3834
rect 19712 3782 19742 3834
rect 19766 3782 19776 3834
rect 19776 3782 19822 3834
rect 19526 3780 19582 3782
rect 19606 3780 19662 3782
rect 19686 3780 19742 3782
rect 19766 3780 19822 3782
rect 26954 3834 27010 3836
rect 27034 3834 27090 3836
rect 27114 3834 27170 3836
rect 27194 3834 27250 3836
rect 26954 3782 27000 3834
rect 27000 3782 27010 3834
rect 27034 3782 27064 3834
rect 27064 3782 27076 3834
rect 27076 3782 27090 3834
rect 27114 3782 27128 3834
rect 27128 3782 27140 3834
rect 27140 3782 27170 3834
rect 27194 3782 27204 3834
rect 27204 3782 27250 3834
rect 26954 3780 27010 3782
rect 27034 3780 27090 3782
rect 27114 3780 27170 3782
rect 27194 3780 27250 3782
rect 8384 3290 8440 3292
rect 8464 3290 8520 3292
rect 8544 3290 8600 3292
rect 8624 3290 8680 3292
rect 8384 3238 8430 3290
rect 8430 3238 8440 3290
rect 8464 3238 8494 3290
rect 8494 3238 8506 3290
rect 8506 3238 8520 3290
rect 8544 3238 8558 3290
rect 8558 3238 8570 3290
rect 8570 3238 8600 3290
rect 8624 3238 8634 3290
rect 8634 3238 8680 3290
rect 8384 3236 8440 3238
rect 8464 3236 8520 3238
rect 8544 3236 8600 3238
rect 8624 3236 8680 3238
rect 15812 3290 15868 3292
rect 15892 3290 15948 3292
rect 15972 3290 16028 3292
rect 16052 3290 16108 3292
rect 15812 3238 15858 3290
rect 15858 3238 15868 3290
rect 15892 3238 15922 3290
rect 15922 3238 15934 3290
rect 15934 3238 15948 3290
rect 15972 3238 15986 3290
rect 15986 3238 15998 3290
rect 15998 3238 16028 3290
rect 16052 3238 16062 3290
rect 16062 3238 16108 3290
rect 15812 3236 15868 3238
rect 15892 3236 15948 3238
rect 15972 3236 16028 3238
rect 16052 3236 16108 3238
rect 23240 3290 23296 3292
rect 23320 3290 23376 3292
rect 23400 3290 23456 3292
rect 23480 3290 23536 3292
rect 23240 3238 23286 3290
rect 23286 3238 23296 3290
rect 23320 3238 23350 3290
rect 23350 3238 23362 3290
rect 23362 3238 23376 3290
rect 23400 3238 23414 3290
rect 23414 3238 23426 3290
rect 23426 3238 23456 3290
rect 23480 3238 23490 3290
rect 23490 3238 23536 3290
rect 23240 3236 23296 3238
rect 23320 3236 23376 3238
rect 23400 3236 23456 3238
rect 23480 3236 23536 3238
rect 4670 2746 4726 2748
rect 4750 2746 4806 2748
rect 4830 2746 4886 2748
rect 4910 2746 4966 2748
rect 4670 2694 4716 2746
rect 4716 2694 4726 2746
rect 4750 2694 4780 2746
rect 4780 2694 4792 2746
rect 4792 2694 4806 2746
rect 4830 2694 4844 2746
rect 4844 2694 4856 2746
rect 4856 2694 4886 2746
rect 4910 2694 4920 2746
rect 4920 2694 4966 2746
rect 4670 2692 4726 2694
rect 4750 2692 4806 2694
rect 4830 2692 4886 2694
rect 4910 2692 4966 2694
rect 12098 2746 12154 2748
rect 12178 2746 12234 2748
rect 12258 2746 12314 2748
rect 12338 2746 12394 2748
rect 12098 2694 12144 2746
rect 12144 2694 12154 2746
rect 12178 2694 12208 2746
rect 12208 2694 12220 2746
rect 12220 2694 12234 2746
rect 12258 2694 12272 2746
rect 12272 2694 12284 2746
rect 12284 2694 12314 2746
rect 12338 2694 12348 2746
rect 12348 2694 12394 2746
rect 12098 2692 12154 2694
rect 12178 2692 12234 2694
rect 12258 2692 12314 2694
rect 12338 2692 12394 2694
rect 19526 2746 19582 2748
rect 19606 2746 19662 2748
rect 19686 2746 19742 2748
rect 19766 2746 19822 2748
rect 19526 2694 19572 2746
rect 19572 2694 19582 2746
rect 19606 2694 19636 2746
rect 19636 2694 19648 2746
rect 19648 2694 19662 2746
rect 19686 2694 19700 2746
rect 19700 2694 19712 2746
rect 19712 2694 19742 2746
rect 19766 2694 19776 2746
rect 19776 2694 19822 2746
rect 19526 2692 19582 2694
rect 19606 2692 19662 2694
rect 19686 2692 19742 2694
rect 19766 2692 19822 2694
rect 26954 2746 27010 2748
rect 27034 2746 27090 2748
rect 27114 2746 27170 2748
rect 27194 2746 27250 2748
rect 26954 2694 27000 2746
rect 27000 2694 27010 2746
rect 27034 2694 27064 2746
rect 27064 2694 27076 2746
rect 27076 2694 27090 2746
rect 27114 2694 27128 2746
rect 27128 2694 27140 2746
rect 27140 2694 27170 2746
rect 27194 2694 27204 2746
rect 27204 2694 27250 2746
rect 26954 2692 27010 2694
rect 27034 2692 27090 2694
rect 27114 2692 27170 2694
rect 27194 2692 27250 2694
rect 30668 4378 30724 4380
rect 30748 4378 30804 4380
rect 30828 4378 30884 4380
rect 30908 4378 30964 4380
rect 30668 4326 30714 4378
rect 30714 4326 30724 4378
rect 30748 4326 30778 4378
rect 30778 4326 30790 4378
rect 30790 4326 30804 4378
rect 30828 4326 30842 4378
rect 30842 4326 30854 4378
rect 30854 4326 30884 4378
rect 30908 4326 30918 4378
rect 30918 4326 30964 4378
rect 30668 4324 30724 4326
rect 30748 4324 30804 4326
rect 30828 4324 30884 4326
rect 30908 4324 30964 4326
rect 30668 3290 30724 3292
rect 30748 3290 30804 3292
rect 30828 3290 30884 3292
rect 30908 3290 30964 3292
rect 30668 3238 30714 3290
rect 30714 3238 30724 3290
rect 30748 3238 30778 3290
rect 30778 3238 30790 3290
rect 30790 3238 30804 3290
rect 30828 3238 30842 3290
rect 30842 3238 30854 3290
rect 30854 3238 30884 3290
rect 30908 3238 30918 3290
rect 30918 3238 30964 3290
rect 30668 3236 30724 3238
rect 30748 3236 30804 3238
rect 30828 3236 30884 3238
rect 30908 3236 30964 3238
rect 8384 2202 8440 2204
rect 8464 2202 8520 2204
rect 8544 2202 8600 2204
rect 8624 2202 8680 2204
rect 8384 2150 8430 2202
rect 8430 2150 8440 2202
rect 8464 2150 8494 2202
rect 8494 2150 8506 2202
rect 8506 2150 8520 2202
rect 8544 2150 8558 2202
rect 8558 2150 8570 2202
rect 8570 2150 8600 2202
rect 8624 2150 8634 2202
rect 8634 2150 8680 2202
rect 8384 2148 8440 2150
rect 8464 2148 8520 2150
rect 8544 2148 8600 2150
rect 8624 2148 8680 2150
rect 15812 2202 15868 2204
rect 15892 2202 15948 2204
rect 15972 2202 16028 2204
rect 16052 2202 16108 2204
rect 15812 2150 15858 2202
rect 15858 2150 15868 2202
rect 15892 2150 15922 2202
rect 15922 2150 15934 2202
rect 15934 2150 15948 2202
rect 15972 2150 15986 2202
rect 15986 2150 15998 2202
rect 15998 2150 16028 2202
rect 16052 2150 16062 2202
rect 16062 2150 16108 2202
rect 15812 2148 15868 2150
rect 15892 2148 15948 2150
rect 15972 2148 16028 2150
rect 16052 2148 16108 2150
rect 23240 2202 23296 2204
rect 23320 2202 23376 2204
rect 23400 2202 23456 2204
rect 23480 2202 23536 2204
rect 23240 2150 23286 2202
rect 23286 2150 23296 2202
rect 23320 2150 23350 2202
rect 23350 2150 23362 2202
rect 23362 2150 23376 2202
rect 23400 2150 23414 2202
rect 23414 2150 23426 2202
rect 23426 2150 23456 2202
rect 23480 2150 23490 2202
rect 23490 2150 23536 2202
rect 23240 2148 23296 2150
rect 23320 2148 23376 2150
rect 23400 2148 23456 2150
rect 23480 2148 23536 2150
rect 30668 2202 30724 2204
rect 30748 2202 30804 2204
rect 30828 2202 30884 2204
rect 30908 2202 30964 2204
rect 30668 2150 30714 2202
rect 30714 2150 30724 2202
rect 30748 2150 30778 2202
rect 30778 2150 30790 2202
rect 30790 2150 30804 2202
rect 30828 2150 30842 2202
rect 30842 2150 30854 2202
rect 30854 2150 30884 2202
rect 30908 2150 30918 2202
rect 30918 2150 30964 2202
rect 30668 2148 30724 2150
rect 30748 2148 30804 2150
rect 30828 2148 30884 2150
rect 30908 2148 30964 2150
rect 31022 1944 31078 2000
<< metal3 >>
rect 31017 29746 31083 29749
rect 31200 29746 32000 29776
rect 31017 29744 32000 29746
rect 31017 29688 31022 29744
rect 31078 29688 32000 29744
rect 31017 29686 32000 29688
rect 31017 29683 31083 29686
rect 31200 29656 32000 29686
rect 8374 29408 8690 29409
rect 8374 29344 8380 29408
rect 8444 29344 8460 29408
rect 8524 29344 8540 29408
rect 8604 29344 8620 29408
rect 8684 29344 8690 29408
rect 8374 29343 8690 29344
rect 15802 29408 16118 29409
rect 15802 29344 15808 29408
rect 15872 29344 15888 29408
rect 15952 29344 15968 29408
rect 16032 29344 16048 29408
rect 16112 29344 16118 29408
rect 15802 29343 16118 29344
rect 23230 29408 23546 29409
rect 23230 29344 23236 29408
rect 23300 29344 23316 29408
rect 23380 29344 23396 29408
rect 23460 29344 23476 29408
rect 23540 29344 23546 29408
rect 23230 29343 23546 29344
rect 30658 29408 30974 29409
rect 30658 29344 30664 29408
rect 30728 29344 30744 29408
rect 30808 29344 30824 29408
rect 30888 29344 30904 29408
rect 30968 29344 30974 29408
rect 30658 29343 30974 29344
rect 4660 28864 4976 28865
rect 4660 28800 4666 28864
rect 4730 28800 4746 28864
rect 4810 28800 4826 28864
rect 4890 28800 4906 28864
rect 4970 28800 4976 28864
rect 4660 28799 4976 28800
rect 12088 28864 12404 28865
rect 12088 28800 12094 28864
rect 12158 28800 12174 28864
rect 12238 28800 12254 28864
rect 12318 28800 12334 28864
rect 12398 28800 12404 28864
rect 12088 28799 12404 28800
rect 19516 28864 19832 28865
rect 19516 28800 19522 28864
rect 19586 28800 19602 28864
rect 19666 28800 19682 28864
rect 19746 28800 19762 28864
rect 19826 28800 19832 28864
rect 19516 28799 19832 28800
rect 26944 28864 27260 28865
rect 26944 28800 26950 28864
rect 27014 28800 27030 28864
rect 27094 28800 27110 28864
rect 27174 28800 27190 28864
rect 27254 28800 27260 28864
rect 26944 28799 27260 28800
rect 8374 28320 8690 28321
rect 8374 28256 8380 28320
rect 8444 28256 8460 28320
rect 8524 28256 8540 28320
rect 8604 28256 8620 28320
rect 8684 28256 8690 28320
rect 8374 28255 8690 28256
rect 15802 28320 16118 28321
rect 15802 28256 15808 28320
rect 15872 28256 15888 28320
rect 15952 28256 15968 28320
rect 16032 28256 16048 28320
rect 16112 28256 16118 28320
rect 15802 28255 16118 28256
rect 23230 28320 23546 28321
rect 23230 28256 23236 28320
rect 23300 28256 23316 28320
rect 23380 28256 23396 28320
rect 23460 28256 23476 28320
rect 23540 28256 23546 28320
rect 23230 28255 23546 28256
rect 30658 28320 30974 28321
rect 30658 28256 30664 28320
rect 30728 28256 30744 28320
rect 30808 28256 30824 28320
rect 30888 28256 30904 28320
rect 30968 28256 30974 28320
rect 30658 28255 30974 28256
rect 4660 27776 4976 27777
rect 4660 27712 4666 27776
rect 4730 27712 4746 27776
rect 4810 27712 4826 27776
rect 4890 27712 4906 27776
rect 4970 27712 4976 27776
rect 4660 27711 4976 27712
rect 12088 27776 12404 27777
rect 12088 27712 12094 27776
rect 12158 27712 12174 27776
rect 12238 27712 12254 27776
rect 12318 27712 12334 27776
rect 12398 27712 12404 27776
rect 12088 27711 12404 27712
rect 19516 27776 19832 27777
rect 19516 27712 19522 27776
rect 19586 27712 19602 27776
rect 19666 27712 19682 27776
rect 19746 27712 19762 27776
rect 19826 27712 19832 27776
rect 19516 27711 19832 27712
rect 26944 27776 27260 27777
rect 26944 27712 26950 27776
rect 27014 27712 27030 27776
rect 27094 27712 27110 27776
rect 27174 27712 27190 27776
rect 27254 27712 27260 27776
rect 26944 27711 27260 27712
rect 8374 27232 8690 27233
rect 8374 27168 8380 27232
rect 8444 27168 8460 27232
rect 8524 27168 8540 27232
rect 8604 27168 8620 27232
rect 8684 27168 8690 27232
rect 8374 27167 8690 27168
rect 15802 27232 16118 27233
rect 15802 27168 15808 27232
rect 15872 27168 15888 27232
rect 15952 27168 15968 27232
rect 16032 27168 16048 27232
rect 16112 27168 16118 27232
rect 15802 27167 16118 27168
rect 23230 27232 23546 27233
rect 23230 27168 23236 27232
rect 23300 27168 23316 27232
rect 23380 27168 23396 27232
rect 23460 27168 23476 27232
rect 23540 27168 23546 27232
rect 23230 27167 23546 27168
rect 30658 27232 30974 27233
rect 30658 27168 30664 27232
rect 30728 27168 30744 27232
rect 30808 27168 30824 27232
rect 30888 27168 30904 27232
rect 30968 27168 30974 27232
rect 30658 27167 30974 27168
rect 4660 26688 4976 26689
rect 4660 26624 4666 26688
rect 4730 26624 4746 26688
rect 4810 26624 4826 26688
rect 4890 26624 4906 26688
rect 4970 26624 4976 26688
rect 4660 26623 4976 26624
rect 12088 26688 12404 26689
rect 12088 26624 12094 26688
rect 12158 26624 12174 26688
rect 12238 26624 12254 26688
rect 12318 26624 12334 26688
rect 12398 26624 12404 26688
rect 12088 26623 12404 26624
rect 19516 26688 19832 26689
rect 19516 26624 19522 26688
rect 19586 26624 19602 26688
rect 19666 26624 19682 26688
rect 19746 26624 19762 26688
rect 19826 26624 19832 26688
rect 19516 26623 19832 26624
rect 26944 26688 27260 26689
rect 26944 26624 26950 26688
rect 27014 26624 27030 26688
rect 27094 26624 27110 26688
rect 27174 26624 27190 26688
rect 27254 26624 27260 26688
rect 26944 26623 27260 26624
rect 8374 26144 8690 26145
rect 8374 26080 8380 26144
rect 8444 26080 8460 26144
rect 8524 26080 8540 26144
rect 8604 26080 8620 26144
rect 8684 26080 8690 26144
rect 8374 26079 8690 26080
rect 15802 26144 16118 26145
rect 15802 26080 15808 26144
rect 15872 26080 15888 26144
rect 15952 26080 15968 26144
rect 16032 26080 16048 26144
rect 16112 26080 16118 26144
rect 15802 26079 16118 26080
rect 23230 26144 23546 26145
rect 23230 26080 23236 26144
rect 23300 26080 23316 26144
rect 23380 26080 23396 26144
rect 23460 26080 23476 26144
rect 23540 26080 23546 26144
rect 23230 26079 23546 26080
rect 30658 26144 30974 26145
rect 30658 26080 30664 26144
rect 30728 26080 30744 26144
rect 30808 26080 30824 26144
rect 30888 26080 30904 26144
rect 30968 26080 30974 26144
rect 30658 26079 30974 26080
rect 31017 25802 31083 25805
rect 31200 25802 32000 25832
rect 31017 25800 32000 25802
rect 31017 25744 31022 25800
rect 31078 25744 32000 25800
rect 31017 25742 32000 25744
rect 31017 25739 31083 25742
rect 31200 25712 32000 25742
rect 4660 25600 4976 25601
rect 4660 25536 4666 25600
rect 4730 25536 4746 25600
rect 4810 25536 4826 25600
rect 4890 25536 4906 25600
rect 4970 25536 4976 25600
rect 4660 25535 4976 25536
rect 12088 25600 12404 25601
rect 12088 25536 12094 25600
rect 12158 25536 12174 25600
rect 12238 25536 12254 25600
rect 12318 25536 12334 25600
rect 12398 25536 12404 25600
rect 12088 25535 12404 25536
rect 19516 25600 19832 25601
rect 19516 25536 19522 25600
rect 19586 25536 19602 25600
rect 19666 25536 19682 25600
rect 19746 25536 19762 25600
rect 19826 25536 19832 25600
rect 19516 25535 19832 25536
rect 26944 25600 27260 25601
rect 26944 25536 26950 25600
rect 27014 25536 27030 25600
rect 27094 25536 27110 25600
rect 27174 25536 27190 25600
rect 27254 25536 27260 25600
rect 26944 25535 27260 25536
rect 8374 25056 8690 25057
rect 8374 24992 8380 25056
rect 8444 24992 8460 25056
rect 8524 24992 8540 25056
rect 8604 24992 8620 25056
rect 8684 24992 8690 25056
rect 8374 24991 8690 24992
rect 15802 25056 16118 25057
rect 15802 24992 15808 25056
rect 15872 24992 15888 25056
rect 15952 24992 15968 25056
rect 16032 24992 16048 25056
rect 16112 24992 16118 25056
rect 15802 24991 16118 24992
rect 23230 25056 23546 25057
rect 23230 24992 23236 25056
rect 23300 24992 23316 25056
rect 23380 24992 23396 25056
rect 23460 24992 23476 25056
rect 23540 24992 23546 25056
rect 23230 24991 23546 24992
rect 30658 25056 30974 25057
rect 30658 24992 30664 25056
rect 30728 24992 30744 25056
rect 30808 24992 30824 25056
rect 30888 24992 30904 25056
rect 30968 24992 30974 25056
rect 30658 24991 30974 24992
rect 4660 24512 4976 24513
rect 4660 24448 4666 24512
rect 4730 24448 4746 24512
rect 4810 24448 4826 24512
rect 4890 24448 4906 24512
rect 4970 24448 4976 24512
rect 4660 24447 4976 24448
rect 12088 24512 12404 24513
rect 12088 24448 12094 24512
rect 12158 24448 12174 24512
rect 12238 24448 12254 24512
rect 12318 24448 12334 24512
rect 12398 24448 12404 24512
rect 12088 24447 12404 24448
rect 19516 24512 19832 24513
rect 19516 24448 19522 24512
rect 19586 24448 19602 24512
rect 19666 24448 19682 24512
rect 19746 24448 19762 24512
rect 19826 24448 19832 24512
rect 19516 24447 19832 24448
rect 26944 24512 27260 24513
rect 26944 24448 26950 24512
rect 27014 24448 27030 24512
rect 27094 24448 27110 24512
rect 27174 24448 27190 24512
rect 27254 24448 27260 24512
rect 26944 24447 27260 24448
rect 8374 23968 8690 23969
rect 8374 23904 8380 23968
rect 8444 23904 8460 23968
rect 8524 23904 8540 23968
rect 8604 23904 8620 23968
rect 8684 23904 8690 23968
rect 8374 23903 8690 23904
rect 15802 23968 16118 23969
rect 15802 23904 15808 23968
rect 15872 23904 15888 23968
rect 15952 23904 15968 23968
rect 16032 23904 16048 23968
rect 16112 23904 16118 23968
rect 15802 23903 16118 23904
rect 23230 23968 23546 23969
rect 23230 23904 23236 23968
rect 23300 23904 23316 23968
rect 23380 23904 23396 23968
rect 23460 23904 23476 23968
rect 23540 23904 23546 23968
rect 23230 23903 23546 23904
rect 30658 23968 30974 23969
rect 30658 23904 30664 23968
rect 30728 23904 30744 23968
rect 30808 23904 30824 23968
rect 30888 23904 30904 23968
rect 30968 23904 30974 23968
rect 30658 23903 30974 23904
rect 4660 23424 4976 23425
rect 4660 23360 4666 23424
rect 4730 23360 4746 23424
rect 4810 23360 4826 23424
rect 4890 23360 4906 23424
rect 4970 23360 4976 23424
rect 4660 23359 4976 23360
rect 12088 23424 12404 23425
rect 12088 23360 12094 23424
rect 12158 23360 12174 23424
rect 12238 23360 12254 23424
rect 12318 23360 12334 23424
rect 12398 23360 12404 23424
rect 12088 23359 12404 23360
rect 19516 23424 19832 23425
rect 19516 23360 19522 23424
rect 19586 23360 19602 23424
rect 19666 23360 19682 23424
rect 19746 23360 19762 23424
rect 19826 23360 19832 23424
rect 19516 23359 19832 23360
rect 26944 23424 27260 23425
rect 26944 23360 26950 23424
rect 27014 23360 27030 23424
rect 27094 23360 27110 23424
rect 27174 23360 27190 23424
rect 27254 23360 27260 23424
rect 26944 23359 27260 23360
rect 8374 22880 8690 22881
rect 8374 22816 8380 22880
rect 8444 22816 8460 22880
rect 8524 22816 8540 22880
rect 8604 22816 8620 22880
rect 8684 22816 8690 22880
rect 8374 22815 8690 22816
rect 15802 22880 16118 22881
rect 15802 22816 15808 22880
rect 15872 22816 15888 22880
rect 15952 22816 15968 22880
rect 16032 22816 16048 22880
rect 16112 22816 16118 22880
rect 15802 22815 16118 22816
rect 23230 22880 23546 22881
rect 23230 22816 23236 22880
rect 23300 22816 23316 22880
rect 23380 22816 23396 22880
rect 23460 22816 23476 22880
rect 23540 22816 23546 22880
rect 23230 22815 23546 22816
rect 30658 22880 30974 22881
rect 30658 22816 30664 22880
rect 30728 22816 30744 22880
rect 30808 22816 30824 22880
rect 30888 22816 30904 22880
rect 30968 22816 30974 22880
rect 30658 22815 30974 22816
rect 4660 22336 4976 22337
rect 4660 22272 4666 22336
rect 4730 22272 4746 22336
rect 4810 22272 4826 22336
rect 4890 22272 4906 22336
rect 4970 22272 4976 22336
rect 4660 22271 4976 22272
rect 12088 22336 12404 22337
rect 12088 22272 12094 22336
rect 12158 22272 12174 22336
rect 12238 22272 12254 22336
rect 12318 22272 12334 22336
rect 12398 22272 12404 22336
rect 12088 22271 12404 22272
rect 19516 22336 19832 22337
rect 19516 22272 19522 22336
rect 19586 22272 19602 22336
rect 19666 22272 19682 22336
rect 19746 22272 19762 22336
rect 19826 22272 19832 22336
rect 19516 22271 19832 22272
rect 26944 22336 27260 22337
rect 26944 22272 26950 22336
rect 27014 22272 27030 22336
rect 27094 22272 27110 22336
rect 27174 22272 27190 22336
rect 27254 22272 27260 22336
rect 26944 22271 27260 22272
rect 31017 21994 31083 21997
rect 31017 21992 31218 21994
rect 31017 21936 31022 21992
rect 31078 21936 31218 21992
rect 31017 21934 31218 21936
rect 31017 21931 31083 21934
rect 31158 21888 31218 21934
rect 31158 21798 32000 21888
rect 8374 21792 8690 21793
rect 8374 21728 8380 21792
rect 8444 21728 8460 21792
rect 8524 21728 8540 21792
rect 8604 21728 8620 21792
rect 8684 21728 8690 21792
rect 8374 21727 8690 21728
rect 15802 21792 16118 21793
rect 15802 21728 15808 21792
rect 15872 21728 15888 21792
rect 15952 21728 15968 21792
rect 16032 21728 16048 21792
rect 16112 21728 16118 21792
rect 15802 21727 16118 21728
rect 23230 21792 23546 21793
rect 23230 21728 23236 21792
rect 23300 21728 23316 21792
rect 23380 21728 23396 21792
rect 23460 21728 23476 21792
rect 23540 21728 23546 21792
rect 23230 21727 23546 21728
rect 30658 21792 30974 21793
rect 30658 21728 30664 21792
rect 30728 21728 30744 21792
rect 30808 21728 30824 21792
rect 30888 21728 30904 21792
rect 30968 21728 30974 21792
rect 31200 21768 32000 21798
rect 30658 21727 30974 21728
rect 4660 21248 4976 21249
rect 4660 21184 4666 21248
rect 4730 21184 4746 21248
rect 4810 21184 4826 21248
rect 4890 21184 4906 21248
rect 4970 21184 4976 21248
rect 4660 21183 4976 21184
rect 12088 21248 12404 21249
rect 12088 21184 12094 21248
rect 12158 21184 12174 21248
rect 12238 21184 12254 21248
rect 12318 21184 12334 21248
rect 12398 21184 12404 21248
rect 12088 21183 12404 21184
rect 19516 21248 19832 21249
rect 19516 21184 19522 21248
rect 19586 21184 19602 21248
rect 19666 21184 19682 21248
rect 19746 21184 19762 21248
rect 19826 21184 19832 21248
rect 19516 21183 19832 21184
rect 26944 21248 27260 21249
rect 26944 21184 26950 21248
rect 27014 21184 27030 21248
rect 27094 21184 27110 21248
rect 27174 21184 27190 21248
rect 27254 21184 27260 21248
rect 26944 21183 27260 21184
rect 8374 20704 8690 20705
rect 8374 20640 8380 20704
rect 8444 20640 8460 20704
rect 8524 20640 8540 20704
rect 8604 20640 8620 20704
rect 8684 20640 8690 20704
rect 8374 20639 8690 20640
rect 15802 20704 16118 20705
rect 15802 20640 15808 20704
rect 15872 20640 15888 20704
rect 15952 20640 15968 20704
rect 16032 20640 16048 20704
rect 16112 20640 16118 20704
rect 15802 20639 16118 20640
rect 23230 20704 23546 20705
rect 23230 20640 23236 20704
rect 23300 20640 23316 20704
rect 23380 20640 23396 20704
rect 23460 20640 23476 20704
rect 23540 20640 23546 20704
rect 23230 20639 23546 20640
rect 30658 20704 30974 20705
rect 30658 20640 30664 20704
rect 30728 20640 30744 20704
rect 30808 20640 30824 20704
rect 30888 20640 30904 20704
rect 30968 20640 30974 20704
rect 30658 20639 30974 20640
rect 4660 20160 4976 20161
rect 4660 20096 4666 20160
rect 4730 20096 4746 20160
rect 4810 20096 4826 20160
rect 4890 20096 4906 20160
rect 4970 20096 4976 20160
rect 4660 20095 4976 20096
rect 12088 20160 12404 20161
rect 12088 20096 12094 20160
rect 12158 20096 12174 20160
rect 12238 20096 12254 20160
rect 12318 20096 12334 20160
rect 12398 20096 12404 20160
rect 12088 20095 12404 20096
rect 19516 20160 19832 20161
rect 19516 20096 19522 20160
rect 19586 20096 19602 20160
rect 19666 20096 19682 20160
rect 19746 20096 19762 20160
rect 19826 20096 19832 20160
rect 19516 20095 19832 20096
rect 26944 20160 27260 20161
rect 26944 20096 26950 20160
rect 27014 20096 27030 20160
rect 27094 20096 27110 20160
rect 27174 20096 27190 20160
rect 27254 20096 27260 20160
rect 26944 20095 27260 20096
rect 8374 19616 8690 19617
rect 8374 19552 8380 19616
rect 8444 19552 8460 19616
rect 8524 19552 8540 19616
rect 8604 19552 8620 19616
rect 8684 19552 8690 19616
rect 8374 19551 8690 19552
rect 15802 19616 16118 19617
rect 15802 19552 15808 19616
rect 15872 19552 15888 19616
rect 15952 19552 15968 19616
rect 16032 19552 16048 19616
rect 16112 19552 16118 19616
rect 15802 19551 16118 19552
rect 23230 19616 23546 19617
rect 23230 19552 23236 19616
rect 23300 19552 23316 19616
rect 23380 19552 23396 19616
rect 23460 19552 23476 19616
rect 23540 19552 23546 19616
rect 23230 19551 23546 19552
rect 30658 19616 30974 19617
rect 30658 19552 30664 19616
rect 30728 19552 30744 19616
rect 30808 19552 30824 19616
rect 30888 19552 30904 19616
rect 30968 19552 30974 19616
rect 30658 19551 30974 19552
rect 4660 19072 4976 19073
rect 4660 19008 4666 19072
rect 4730 19008 4746 19072
rect 4810 19008 4826 19072
rect 4890 19008 4906 19072
rect 4970 19008 4976 19072
rect 4660 19007 4976 19008
rect 12088 19072 12404 19073
rect 12088 19008 12094 19072
rect 12158 19008 12174 19072
rect 12238 19008 12254 19072
rect 12318 19008 12334 19072
rect 12398 19008 12404 19072
rect 12088 19007 12404 19008
rect 19516 19072 19832 19073
rect 19516 19008 19522 19072
rect 19586 19008 19602 19072
rect 19666 19008 19682 19072
rect 19746 19008 19762 19072
rect 19826 19008 19832 19072
rect 19516 19007 19832 19008
rect 26944 19072 27260 19073
rect 26944 19008 26950 19072
rect 27014 19008 27030 19072
rect 27094 19008 27110 19072
rect 27174 19008 27190 19072
rect 27254 19008 27260 19072
rect 26944 19007 27260 19008
rect 8374 18528 8690 18529
rect 8374 18464 8380 18528
rect 8444 18464 8460 18528
rect 8524 18464 8540 18528
rect 8604 18464 8620 18528
rect 8684 18464 8690 18528
rect 8374 18463 8690 18464
rect 15802 18528 16118 18529
rect 15802 18464 15808 18528
rect 15872 18464 15888 18528
rect 15952 18464 15968 18528
rect 16032 18464 16048 18528
rect 16112 18464 16118 18528
rect 15802 18463 16118 18464
rect 23230 18528 23546 18529
rect 23230 18464 23236 18528
rect 23300 18464 23316 18528
rect 23380 18464 23396 18528
rect 23460 18464 23476 18528
rect 23540 18464 23546 18528
rect 23230 18463 23546 18464
rect 30658 18528 30974 18529
rect 30658 18464 30664 18528
rect 30728 18464 30744 18528
rect 30808 18464 30824 18528
rect 30888 18464 30904 18528
rect 30968 18464 30974 18528
rect 30658 18463 30974 18464
rect 4660 17984 4976 17985
rect 4660 17920 4666 17984
rect 4730 17920 4746 17984
rect 4810 17920 4826 17984
rect 4890 17920 4906 17984
rect 4970 17920 4976 17984
rect 4660 17919 4976 17920
rect 12088 17984 12404 17985
rect 12088 17920 12094 17984
rect 12158 17920 12174 17984
rect 12238 17920 12254 17984
rect 12318 17920 12334 17984
rect 12398 17920 12404 17984
rect 12088 17919 12404 17920
rect 19516 17984 19832 17985
rect 19516 17920 19522 17984
rect 19586 17920 19602 17984
rect 19666 17920 19682 17984
rect 19746 17920 19762 17984
rect 19826 17920 19832 17984
rect 19516 17919 19832 17920
rect 26944 17984 27260 17985
rect 26944 17920 26950 17984
rect 27014 17920 27030 17984
rect 27094 17920 27110 17984
rect 27174 17920 27190 17984
rect 27254 17920 27260 17984
rect 26944 17919 27260 17920
rect 31017 17914 31083 17917
rect 31200 17914 32000 17944
rect 31017 17912 32000 17914
rect 31017 17856 31022 17912
rect 31078 17856 32000 17912
rect 31017 17854 32000 17856
rect 31017 17851 31083 17854
rect 31200 17824 32000 17854
rect 8374 17440 8690 17441
rect 8374 17376 8380 17440
rect 8444 17376 8460 17440
rect 8524 17376 8540 17440
rect 8604 17376 8620 17440
rect 8684 17376 8690 17440
rect 8374 17375 8690 17376
rect 15802 17440 16118 17441
rect 15802 17376 15808 17440
rect 15872 17376 15888 17440
rect 15952 17376 15968 17440
rect 16032 17376 16048 17440
rect 16112 17376 16118 17440
rect 15802 17375 16118 17376
rect 23230 17440 23546 17441
rect 23230 17376 23236 17440
rect 23300 17376 23316 17440
rect 23380 17376 23396 17440
rect 23460 17376 23476 17440
rect 23540 17376 23546 17440
rect 23230 17375 23546 17376
rect 30658 17440 30974 17441
rect 30658 17376 30664 17440
rect 30728 17376 30744 17440
rect 30808 17376 30824 17440
rect 30888 17376 30904 17440
rect 30968 17376 30974 17440
rect 30658 17375 30974 17376
rect 4660 16896 4976 16897
rect 4660 16832 4666 16896
rect 4730 16832 4746 16896
rect 4810 16832 4826 16896
rect 4890 16832 4906 16896
rect 4970 16832 4976 16896
rect 4660 16831 4976 16832
rect 12088 16896 12404 16897
rect 12088 16832 12094 16896
rect 12158 16832 12174 16896
rect 12238 16832 12254 16896
rect 12318 16832 12334 16896
rect 12398 16832 12404 16896
rect 12088 16831 12404 16832
rect 19516 16896 19832 16897
rect 19516 16832 19522 16896
rect 19586 16832 19602 16896
rect 19666 16832 19682 16896
rect 19746 16832 19762 16896
rect 19826 16832 19832 16896
rect 19516 16831 19832 16832
rect 26944 16896 27260 16897
rect 26944 16832 26950 16896
rect 27014 16832 27030 16896
rect 27094 16832 27110 16896
rect 27174 16832 27190 16896
rect 27254 16832 27260 16896
rect 26944 16831 27260 16832
rect 8374 16352 8690 16353
rect 8374 16288 8380 16352
rect 8444 16288 8460 16352
rect 8524 16288 8540 16352
rect 8604 16288 8620 16352
rect 8684 16288 8690 16352
rect 8374 16287 8690 16288
rect 15802 16352 16118 16353
rect 15802 16288 15808 16352
rect 15872 16288 15888 16352
rect 15952 16288 15968 16352
rect 16032 16288 16048 16352
rect 16112 16288 16118 16352
rect 15802 16287 16118 16288
rect 23230 16352 23546 16353
rect 23230 16288 23236 16352
rect 23300 16288 23316 16352
rect 23380 16288 23396 16352
rect 23460 16288 23476 16352
rect 23540 16288 23546 16352
rect 23230 16287 23546 16288
rect 30658 16352 30974 16353
rect 30658 16288 30664 16352
rect 30728 16288 30744 16352
rect 30808 16288 30824 16352
rect 30888 16288 30904 16352
rect 30968 16288 30974 16352
rect 30658 16287 30974 16288
rect 4660 15808 4976 15809
rect 4660 15744 4666 15808
rect 4730 15744 4746 15808
rect 4810 15744 4826 15808
rect 4890 15744 4906 15808
rect 4970 15744 4976 15808
rect 4660 15743 4976 15744
rect 12088 15808 12404 15809
rect 12088 15744 12094 15808
rect 12158 15744 12174 15808
rect 12238 15744 12254 15808
rect 12318 15744 12334 15808
rect 12398 15744 12404 15808
rect 12088 15743 12404 15744
rect 19516 15808 19832 15809
rect 19516 15744 19522 15808
rect 19586 15744 19602 15808
rect 19666 15744 19682 15808
rect 19746 15744 19762 15808
rect 19826 15744 19832 15808
rect 19516 15743 19832 15744
rect 26944 15808 27260 15809
rect 26944 15744 26950 15808
rect 27014 15744 27030 15808
rect 27094 15744 27110 15808
rect 27174 15744 27190 15808
rect 27254 15744 27260 15808
rect 26944 15743 27260 15744
rect 8374 15264 8690 15265
rect 8374 15200 8380 15264
rect 8444 15200 8460 15264
rect 8524 15200 8540 15264
rect 8604 15200 8620 15264
rect 8684 15200 8690 15264
rect 8374 15199 8690 15200
rect 15802 15264 16118 15265
rect 15802 15200 15808 15264
rect 15872 15200 15888 15264
rect 15952 15200 15968 15264
rect 16032 15200 16048 15264
rect 16112 15200 16118 15264
rect 15802 15199 16118 15200
rect 23230 15264 23546 15265
rect 23230 15200 23236 15264
rect 23300 15200 23316 15264
rect 23380 15200 23396 15264
rect 23460 15200 23476 15264
rect 23540 15200 23546 15264
rect 23230 15199 23546 15200
rect 30658 15264 30974 15265
rect 30658 15200 30664 15264
rect 30728 15200 30744 15264
rect 30808 15200 30824 15264
rect 30888 15200 30904 15264
rect 30968 15200 30974 15264
rect 30658 15199 30974 15200
rect 4660 14720 4976 14721
rect 4660 14656 4666 14720
rect 4730 14656 4746 14720
rect 4810 14656 4826 14720
rect 4890 14656 4906 14720
rect 4970 14656 4976 14720
rect 4660 14655 4976 14656
rect 12088 14720 12404 14721
rect 12088 14656 12094 14720
rect 12158 14656 12174 14720
rect 12238 14656 12254 14720
rect 12318 14656 12334 14720
rect 12398 14656 12404 14720
rect 12088 14655 12404 14656
rect 19516 14720 19832 14721
rect 19516 14656 19522 14720
rect 19586 14656 19602 14720
rect 19666 14656 19682 14720
rect 19746 14656 19762 14720
rect 19826 14656 19832 14720
rect 19516 14655 19832 14656
rect 26944 14720 27260 14721
rect 26944 14656 26950 14720
rect 27014 14656 27030 14720
rect 27094 14656 27110 14720
rect 27174 14656 27190 14720
rect 27254 14656 27260 14720
rect 26944 14655 27260 14656
rect 8374 14176 8690 14177
rect 8374 14112 8380 14176
rect 8444 14112 8460 14176
rect 8524 14112 8540 14176
rect 8604 14112 8620 14176
rect 8684 14112 8690 14176
rect 8374 14111 8690 14112
rect 15802 14176 16118 14177
rect 15802 14112 15808 14176
rect 15872 14112 15888 14176
rect 15952 14112 15968 14176
rect 16032 14112 16048 14176
rect 16112 14112 16118 14176
rect 15802 14111 16118 14112
rect 23230 14176 23546 14177
rect 23230 14112 23236 14176
rect 23300 14112 23316 14176
rect 23380 14112 23396 14176
rect 23460 14112 23476 14176
rect 23540 14112 23546 14176
rect 23230 14111 23546 14112
rect 30658 14176 30974 14177
rect 30658 14112 30664 14176
rect 30728 14112 30744 14176
rect 30808 14112 30824 14176
rect 30888 14112 30904 14176
rect 30968 14112 30974 14176
rect 30658 14111 30974 14112
rect 31017 13970 31083 13973
rect 31200 13970 32000 14000
rect 31017 13968 32000 13970
rect 31017 13912 31022 13968
rect 31078 13912 32000 13968
rect 31017 13910 32000 13912
rect 31017 13907 31083 13910
rect 31200 13880 32000 13910
rect 4660 13632 4976 13633
rect 4660 13568 4666 13632
rect 4730 13568 4746 13632
rect 4810 13568 4826 13632
rect 4890 13568 4906 13632
rect 4970 13568 4976 13632
rect 4660 13567 4976 13568
rect 12088 13632 12404 13633
rect 12088 13568 12094 13632
rect 12158 13568 12174 13632
rect 12238 13568 12254 13632
rect 12318 13568 12334 13632
rect 12398 13568 12404 13632
rect 12088 13567 12404 13568
rect 19516 13632 19832 13633
rect 19516 13568 19522 13632
rect 19586 13568 19602 13632
rect 19666 13568 19682 13632
rect 19746 13568 19762 13632
rect 19826 13568 19832 13632
rect 19516 13567 19832 13568
rect 26944 13632 27260 13633
rect 26944 13568 26950 13632
rect 27014 13568 27030 13632
rect 27094 13568 27110 13632
rect 27174 13568 27190 13632
rect 27254 13568 27260 13632
rect 26944 13567 27260 13568
rect 8374 13088 8690 13089
rect 8374 13024 8380 13088
rect 8444 13024 8460 13088
rect 8524 13024 8540 13088
rect 8604 13024 8620 13088
rect 8684 13024 8690 13088
rect 8374 13023 8690 13024
rect 15802 13088 16118 13089
rect 15802 13024 15808 13088
rect 15872 13024 15888 13088
rect 15952 13024 15968 13088
rect 16032 13024 16048 13088
rect 16112 13024 16118 13088
rect 15802 13023 16118 13024
rect 23230 13088 23546 13089
rect 23230 13024 23236 13088
rect 23300 13024 23316 13088
rect 23380 13024 23396 13088
rect 23460 13024 23476 13088
rect 23540 13024 23546 13088
rect 23230 13023 23546 13024
rect 30658 13088 30974 13089
rect 30658 13024 30664 13088
rect 30728 13024 30744 13088
rect 30808 13024 30824 13088
rect 30888 13024 30904 13088
rect 30968 13024 30974 13088
rect 30658 13023 30974 13024
rect 4660 12544 4976 12545
rect 4660 12480 4666 12544
rect 4730 12480 4746 12544
rect 4810 12480 4826 12544
rect 4890 12480 4906 12544
rect 4970 12480 4976 12544
rect 4660 12479 4976 12480
rect 12088 12544 12404 12545
rect 12088 12480 12094 12544
rect 12158 12480 12174 12544
rect 12238 12480 12254 12544
rect 12318 12480 12334 12544
rect 12398 12480 12404 12544
rect 12088 12479 12404 12480
rect 19516 12544 19832 12545
rect 19516 12480 19522 12544
rect 19586 12480 19602 12544
rect 19666 12480 19682 12544
rect 19746 12480 19762 12544
rect 19826 12480 19832 12544
rect 19516 12479 19832 12480
rect 26944 12544 27260 12545
rect 26944 12480 26950 12544
rect 27014 12480 27030 12544
rect 27094 12480 27110 12544
rect 27174 12480 27190 12544
rect 27254 12480 27260 12544
rect 26944 12479 27260 12480
rect 8374 12000 8690 12001
rect 8374 11936 8380 12000
rect 8444 11936 8460 12000
rect 8524 11936 8540 12000
rect 8604 11936 8620 12000
rect 8684 11936 8690 12000
rect 8374 11935 8690 11936
rect 15802 12000 16118 12001
rect 15802 11936 15808 12000
rect 15872 11936 15888 12000
rect 15952 11936 15968 12000
rect 16032 11936 16048 12000
rect 16112 11936 16118 12000
rect 15802 11935 16118 11936
rect 23230 12000 23546 12001
rect 23230 11936 23236 12000
rect 23300 11936 23316 12000
rect 23380 11936 23396 12000
rect 23460 11936 23476 12000
rect 23540 11936 23546 12000
rect 23230 11935 23546 11936
rect 30658 12000 30974 12001
rect 30658 11936 30664 12000
rect 30728 11936 30744 12000
rect 30808 11936 30824 12000
rect 30888 11936 30904 12000
rect 30968 11936 30974 12000
rect 30658 11935 30974 11936
rect 4660 11456 4976 11457
rect 4660 11392 4666 11456
rect 4730 11392 4746 11456
rect 4810 11392 4826 11456
rect 4890 11392 4906 11456
rect 4970 11392 4976 11456
rect 4660 11391 4976 11392
rect 12088 11456 12404 11457
rect 12088 11392 12094 11456
rect 12158 11392 12174 11456
rect 12238 11392 12254 11456
rect 12318 11392 12334 11456
rect 12398 11392 12404 11456
rect 12088 11391 12404 11392
rect 19516 11456 19832 11457
rect 19516 11392 19522 11456
rect 19586 11392 19602 11456
rect 19666 11392 19682 11456
rect 19746 11392 19762 11456
rect 19826 11392 19832 11456
rect 19516 11391 19832 11392
rect 26944 11456 27260 11457
rect 26944 11392 26950 11456
rect 27014 11392 27030 11456
rect 27094 11392 27110 11456
rect 27174 11392 27190 11456
rect 27254 11392 27260 11456
rect 26944 11391 27260 11392
rect 8374 10912 8690 10913
rect 8374 10848 8380 10912
rect 8444 10848 8460 10912
rect 8524 10848 8540 10912
rect 8604 10848 8620 10912
rect 8684 10848 8690 10912
rect 8374 10847 8690 10848
rect 15802 10912 16118 10913
rect 15802 10848 15808 10912
rect 15872 10848 15888 10912
rect 15952 10848 15968 10912
rect 16032 10848 16048 10912
rect 16112 10848 16118 10912
rect 15802 10847 16118 10848
rect 23230 10912 23546 10913
rect 23230 10848 23236 10912
rect 23300 10848 23316 10912
rect 23380 10848 23396 10912
rect 23460 10848 23476 10912
rect 23540 10848 23546 10912
rect 23230 10847 23546 10848
rect 30658 10912 30974 10913
rect 30658 10848 30664 10912
rect 30728 10848 30744 10912
rect 30808 10848 30824 10912
rect 30888 10848 30904 10912
rect 30968 10848 30974 10912
rect 30658 10847 30974 10848
rect 4660 10368 4976 10369
rect 4660 10304 4666 10368
rect 4730 10304 4746 10368
rect 4810 10304 4826 10368
rect 4890 10304 4906 10368
rect 4970 10304 4976 10368
rect 4660 10303 4976 10304
rect 12088 10368 12404 10369
rect 12088 10304 12094 10368
rect 12158 10304 12174 10368
rect 12238 10304 12254 10368
rect 12318 10304 12334 10368
rect 12398 10304 12404 10368
rect 12088 10303 12404 10304
rect 19516 10368 19832 10369
rect 19516 10304 19522 10368
rect 19586 10304 19602 10368
rect 19666 10304 19682 10368
rect 19746 10304 19762 10368
rect 19826 10304 19832 10368
rect 19516 10303 19832 10304
rect 26944 10368 27260 10369
rect 26944 10304 26950 10368
rect 27014 10304 27030 10368
rect 27094 10304 27110 10368
rect 27174 10304 27190 10368
rect 27254 10304 27260 10368
rect 26944 10303 27260 10304
rect 31017 10026 31083 10029
rect 31200 10026 32000 10056
rect 31017 10024 32000 10026
rect 31017 9968 31022 10024
rect 31078 9968 32000 10024
rect 31017 9966 32000 9968
rect 31017 9963 31083 9966
rect 31200 9936 32000 9966
rect 8374 9824 8690 9825
rect 8374 9760 8380 9824
rect 8444 9760 8460 9824
rect 8524 9760 8540 9824
rect 8604 9760 8620 9824
rect 8684 9760 8690 9824
rect 8374 9759 8690 9760
rect 15802 9824 16118 9825
rect 15802 9760 15808 9824
rect 15872 9760 15888 9824
rect 15952 9760 15968 9824
rect 16032 9760 16048 9824
rect 16112 9760 16118 9824
rect 15802 9759 16118 9760
rect 23230 9824 23546 9825
rect 23230 9760 23236 9824
rect 23300 9760 23316 9824
rect 23380 9760 23396 9824
rect 23460 9760 23476 9824
rect 23540 9760 23546 9824
rect 23230 9759 23546 9760
rect 30658 9824 30974 9825
rect 30658 9760 30664 9824
rect 30728 9760 30744 9824
rect 30808 9760 30824 9824
rect 30888 9760 30904 9824
rect 30968 9760 30974 9824
rect 30658 9759 30974 9760
rect 4660 9280 4976 9281
rect 4660 9216 4666 9280
rect 4730 9216 4746 9280
rect 4810 9216 4826 9280
rect 4890 9216 4906 9280
rect 4970 9216 4976 9280
rect 4660 9215 4976 9216
rect 12088 9280 12404 9281
rect 12088 9216 12094 9280
rect 12158 9216 12174 9280
rect 12238 9216 12254 9280
rect 12318 9216 12334 9280
rect 12398 9216 12404 9280
rect 12088 9215 12404 9216
rect 19516 9280 19832 9281
rect 19516 9216 19522 9280
rect 19586 9216 19602 9280
rect 19666 9216 19682 9280
rect 19746 9216 19762 9280
rect 19826 9216 19832 9280
rect 19516 9215 19832 9216
rect 26944 9280 27260 9281
rect 26944 9216 26950 9280
rect 27014 9216 27030 9280
rect 27094 9216 27110 9280
rect 27174 9216 27190 9280
rect 27254 9216 27260 9280
rect 26944 9215 27260 9216
rect 8374 8736 8690 8737
rect 8374 8672 8380 8736
rect 8444 8672 8460 8736
rect 8524 8672 8540 8736
rect 8604 8672 8620 8736
rect 8684 8672 8690 8736
rect 8374 8671 8690 8672
rect 15802 8736 16118 8737
rect 15802 8672 15808 8736
rect 15872 8672 15888 8736
rect 15952 8672 15968 8736
rect 16032 8672 16048 8736
rect 16112 8672 16118 8736
rect 15802 8671 16118 8672
rect 23230 8736 23546 8737
rect 23230 8672 23236 8736
rect 23300 8672 23316 8736
rect 23380 8672 23396 8736
rect 23460 8672 23476 8736
rect 23540 8672 23546 8736
rect 23230 8671 23546 8672
rect 30658 8736 30974 8737
rect 30658 8672 30664 8736
rect 30728 8672 30744 8736
rect 30808 8672 30824 8736
rect 30888 8672 30904 8736
rect 30968 8672 30974 8736
rect 30658 8671 30974 8672
rect 4660 8192 4976 8193
rect 4660 8128 4666 8192
rect 4730 8128 4746 8192
rect 4810 8128 4826 8192
rect 4890 8128 4906 8192
rect 4970 8128 4976 8192
rect 4660 8127 4976 8128
rect 12088 8192 12404 8193
rect 12088 8128 12094 8192
rect 12158 8128 12174 8192
rect 12238 8128 12254 8192
rect 12318 8128 12334 8192
rect 12398 8128 12404 8192
rect 12088 8127 12404 8128
rect 19516 8192 19832 8193
rect 19516 8128 19522 8192
rect 19586 8128 19602 8192
rect 19666 8128 19682 8192
rect 19746 8128 19762 8192
rect 19826 8128 19832 8192
rect 19516 8127 19832 8128
rect 26944 8192 27260 8193
rect 26944 8128 26950 8192
rect 27014 8128 27030 8192
rect 27094 8128 27110 8192
rect 27174 8128 27190 8192
rect 27254 8128 27260 8192
rect 26944 8127 27260 8128
rect 8374 7648 8690 7649
rect 8374 7584 8380 7648
rect 8444 7584 8460 7648
rect 8524 7584 8540 7648
rect 8604 7584 8620 7648
rect 8684 7584 8690 7648
rect 8374 7583 8690 7584
rect 15802 7648 16118 7649
rect 15802 7584 15808 7648
rect 15872 7584 15888 7648
rect 15952 7584 15968 7648
rect 16032 7584 16048 7648
rect 16112 7584 16118 7648
rect 15802 7583 16118 7584
rect 23230 7648 23546 7649
rect 23230 7584 23236 7648
rect 23300 7584 23316 7648
rect 23380 7584 23396 7648
rect 23460 7584 23476 7648
rect 23540 7584 23546 7648
rect 23230 7583 23546 7584
rect 30658 7648 30974 7649
rect 30658 7584 30664 7648
rect 30728 7584 30744 7648
rect 30808 7584 30824 7648
rect 30888 7584 30904 7648
rect 30968 7584 30974 7648
rect 30658 7583 30974 7584
rect 4660 7104 4976 7105
rect 4660 7040 4666 7104
rect 4730 7040 4746 7104
rect 4810 7040 4826 7104
rect 4890 7040 4906 7104
rect 4970 7040 4976 7104
rect 4660 7039 4976 7040
rect 12088 7104 12404 7105
rect 12088 7040 12094 7104
rect 12158 7040 12174 7104
rect 12238 7040 12254 7104
rect 12318 7040 12334 7104
rect 12398 7040 12404 7104
rect 12088 7039 12404 7040
rect 19516 7104 19832 7105
rect 19516 7040 19522 7104
rect 19586 7040 19602 7104
rect 19666 7040 19682 7104
rect 19746 7040 19762 7104
rect 19826 7040 19832 7104
rect 19516 7039 19832 7040
rect 26944 7104 27260 7105
rect 26944 7040 26950 7104
rect 27014 7040 27030 7104
rect 27094 7040 27110 7104
rect 27174 7040 27190 7104
rect 27254 7040 27260 7104
rect 26944 7039 27260 7040
rect 8374 6560 8690 6561
rect 8374 6496 8380 6560
rect 8444 6496 8460 6560
rect 8524 6496 8540 6560
rect 8604 6496 8620 6560
rect 8684 6496 8690 6560
rect 8374 6495 8690 6496
rect 15802 6560 16118 6561
rect 15802 6496 15808 6560
rect 15872 6496 15888 6560
rect 15952 6496 15968 6560
rect 16032 6496 16048 6560
rect 16112 6496 16118 6560
rect 15802 6495 16118 6496
rect 23230 6560 23546 6561
rect 23230 6496 23236 6560
rect 23300 6496 23316 6560
rect 23380 6496 23396 6560
rect 23460 6496 23476 6560
rect 23540 6496 23546 6560
rect 23230 6495 23546 6496
rect 30658 6560 30974 6561
rect 30658 6496 30664 6560
rect 30728 6496 30744 6560
rect 30808 6496 30824 6560
rect 30888 6496 30904 6560
rect 30968 6496 30974 6560
rect 30658 6495 30974 6496
rect 31017 6082 31083 6085
rect 31200 6082 32000 6112
rect 31017 6080 32000 6082
rect 31017 6024 31022 6080
rect 31078 6024 32000 6080
rect 31017 6022 32000 6024
rect 31017 6019 31083 6022
rect 4660 6016 4976 6017
rect 4660 5952 4666 6016
rect 4730 5952 4746 6016
rect 4810 5952 4826 6016
rect 4890 5952 4906 6016
rect 4970 5952 4976 6016
rect 4660 5951 4976 5952
rect 12088 6016 12404 6017
rect 12088 5952 12094 6016
rect 12158 5952 12174 6016
rect 12238 5952 12254 6016
rect 12318 5952 12334 6016
rect 12398 5952 12404 6016
rect 12088 5951 12404 5952
rect 19516 6016 19832 6017
rect 19516 5952 19522 6016
rect 19586 5952 19602 6016
rect 19666 5952 19682 6016
rect 19746 5952 19762 6016
rect 19826 5952 19832 6016
rect 19516 5951 19832 5952
rect 26944 6016 27260 6017
rect 26944 5952 26950 6016
rect 27014 5952 27030 6016
rect 27094 5952 27110 6016
rect 27174 5952 27190 6016
rect 27254 5952 27260 6016
rect 31200 5992 32000 6022
rect 26944 5951 27260 5952
rect 8374 5472 8690 5473
rect 8374 5408 8380 5472
rect 8444 5408 8460 5472
rect 8524 5408 8540 5472
rect 8604 5408 8620 5472
rect 8684 5408 8690 5472
rect 8374 5407 8690 5408
rect 15802 5472 16118 5473
rect 15802 5408 15808 5472
rect 15872 5408 15888 5472
rect 15952 5408 15968 5472
rect 16032 5408 16048 5472
rect 16112 5408 16118 5472
rect 15802 5407 16118 5408
rect 23230 5472 23546 5473
rect 23230 5408 23236 5472
rect 23300 5408 23316 5472
rect 23380 5408 23396 5472
rect 23460 5408 23476 5472
rect 23540 5408 23546 5472
rect 23230 5407 23546 5408
rect 30658 5472 30974 5473
rect 30658 5408 30664 5472
rect 30728 5408 30744 5472
rect 30808 5408 30824 5472
rect 30888 5408 30904 5472
rect 30968 5408 30974 5472
rect 30658 5407 30974 5408
rect 4660 4928 4976 4929
rect 4660 4864 4666 4928
rect 4730 4864 4746 4928
rect 4810 4864 4826 4928
rect 4890 4864 4906 4928
rect 4970 4864 4976 4928
rect 4660 4863 4976 4864
rect 12088 4928 12404 4929
rect 12088 4864 12094 4928
rect 12158 4864 12174 4928
rect 12238 4864 12254 4928
rect 12318 4864 12334 4928
rect 12398 4864 12404 4928
rect 12088 4863 12404 4864
rect 19516 4928 19832 4929
rect 19516 4864 19522 4928
rect 19586 4864 19602 4928
rect 19666 4864 19682 4928
rect 19746 4864 19762 4928
rect 19826 4864 19832 4928
rect 19516 4863 19832 4864
rect 26944 4928 27260 4929
rect 26944 4864 26950 4928
rect 27014 4864 27030 4928
rect 27094 4864 27110 4928
rect 27174 4864 27190 4928
rect 27254 4864 27260 4928
rect 26944 4863 27260 4864
rect 8374 4384 8690 4385
rect 8374 4320 8380 4384
rect 8444 4320 8460 4384
rect 8524 4320 8540 4384
rect 8604 4320 8620 4384
rect 8684 4320 8690 4384
rect 8374 4319 8690 4320
rect 15802 4384 16118 4385
rect 15802 4320 15808 4384
rect 15872 4320 15888 4384
rect 15952 4320 15968 4384
rect 16032 4320 16048 4384
rect 16112 4320 16118 4384
rect 15802 4319 16118 4320
rect 23230 4384 23546 4385
rect 23230 4320 23236 4384
rect 23300 4320 23316 4384
rect 23380 4320 23396 4384
rect 23460 4320 23476 4384
rect 23540 4320 23546 4384
rect 23230 4319 23546 4320
rect 30658 4384 30974 4385
rect 30658 4320 30664 4384
rect 30728 4320 30744 4384
rect 30808 4320 30824 4384
rect 30888 4320 30904 4384
rect 30968 4320 30974 4384
rect 30658 4319 30974 4320
rect 4660 3840 4976 3841
rect 4660 3776 4666 3840
rect 4730 3776 4746 3840
rect 4810 3776 4826 3840
rect 4890 3776 4906 3840
rect 4970 3776 4976 3840
rect 4660 3775 4976 3776
rect 12088 3840 12404 3841
rect 12088 3776 12094 3840
rect 12158 3776 12174 3840
rect 12238 3776 12254 3840
rect 12318 3776 12334 3840
rect 12398 3776 12404 3840
rect 12088 3775 12404 3776
rect 19516 3840 19832 3841
rect 19516 3776 19522 3840
rect 19586 3776 19602 3840
rect 19666 3776 19682 3840
rect 19746 3776 19762 3840
rect 19826 3776 19832 3840
rect 19516 3775 19832 3776
rect 26944 3840 27260 3841
rect 26944 3776 26950 3840
rect 27014 3776 27030 3840
rect 27094 3776 27110 3840
rect 27174 3776 27190 3840
rect 27254 3776 27260 3840
rect 26944 3775 27260 3776
rect 8374 3296 8690 3297
rect 8374 3232 8380 3296
rect 8444 3232 8460 3296
rect 8524 3232 8540 3296
rect 8604 3232 8620 3296
rect 8684 3232 8690 3296
rect 8374 3231 8690 3232
rect 15802 3296 16118 3297
rect 15802 3232 15808 3296
rect 15872 3232 15888 3296
rect 15952 3232 15968 3296
rect 16032 3232 16048 3296
rect 16112 3232 16118 3296
rect 15802 3231 16118 3232
rect 23230 3296 23546 3297
rect 23230 3232 23236 3296
rect 23300 3232 23316 3296
rect 23380 3232 23396 3296
rect 23460 3232 23476 3296
rect 23540 3232 23546 3296
rect 23230 3231 23546 3232
rect 30658 3296 30974 3297
rect 30658 3232 30664 3296
rect 30728 3232 30744 3296
rect 30808 3232 30824 3296
rect 30888 3232 30904 3296
rect 30968 3232 30974 3296
rect 30658 3231 30974 3232
rect 4660 2752 4976 2753
rect 4660 2688 4666 2752
rect 4730 2688 4746 2752
rect 4810 2688 4826 2752
rect 4890 2688 4906 2752
rect 4970 2688 4976 2752
rect 4660 2687 4976 2688
rect 12088 2752 12404 2753
rect 12088 2688 12094 2752
rect 12158 2688 12174 2752
rect 12238 2688 12254 2752
rect 12318 2688 12334 2752
rect 12398 2688 12404 2752
rect 12088 2687 12404 2688
rect 19516 2752 19832 2753
rect 19516 2688 19522 2752
rect 19586 2688 19602 2752
rect 19666 2688 19682 2752
rect 19746 2688 19762 2752
rect 19826 2688 19832 2752
rect 19516 2687 19832 2688
rect 26944 2752 27260 2753
rect 26944 2688 26950 2752
rect 27014 2688 27030 2752
rect 27094 2688 27110 2752
rect 27174 2688 27190 2752
rect 27254 2688 27260 2752
rect 26944 2687 27260 2688
rect 8374 2208 8690 2209
rect 8374 2144 8380 2208
rect 8444 2144 8460 2208
rect 8524 2144 8540 2208
rect 8604 2144 8620 2208
rect 8684 2144 8690 2208
rect 8374 2143 8690 2144
rect 15802 2208 16118 2209
rect 15802 2144 15808 2208
rect 15872 2144 15888 2208
rect 15952 2144 15968 2208
rect 16032 2144 16048 2208
rect 16112 2144 16118 2208
rect 15802 2143 16118 2144
rect 23230 2208 23546 2209
rect 23230 2144 23236 2208
rect 23300 2144 23316 2208
rect 23380 2144 23396 2208
rect 23460 2144 23476 2208
rect 23540 2144 23546 2208
rect 23230 2143 23546 2144
rect 30658 2208 30974 2209
rect 30658 2144 30664 2208
rect 30728 2144 30744 2208
rect 30808 2144 30824 2208
rect 30888 2144 30904 2208
rect 30968 2144 30974 2208
rect 30658 2143 30974 2144
rect 31200 2138 32000 2168
rect 31158 2048 32000 2138
rect 31017 2002 31083 2005
rect 31158 2002 31218 2048
rect 31017 2000 31218 2002
rect 31017 1944 31022 2000
rect 31078 1944 31218 2000
rect 31017 1942 31218 1944
rect 31017 1939 31083 1942
<< via3 >>
rect 8380 29404 8444 29408
rect 8380 29348 8384 29404
rect 8384 29348 8440 29404
rect 8440 29348 8444 29404
rect 8380 29344 8444 29348
rect 8460 29404 8524 29408
rect 8460 29348 8464 29404
rect 8464 29348 8520 29404
rect 8520 29348 8524 29404
rect 8460 29344 8524 29348
rect 8540 29404 8604 29408
rect 8540 29348 8544 29404
rect 8544 29348 8600 29404
rect 8600 29348 8604 29404
rect 8540 29344 8604 29348
rect 8620 29404 8684 29408
rect 8620 29348 8624 29404
rect 8624 29348 8680 29404
rect 8680 29348 8684 29404
rect 8620 29344 8684 29348
rect 15808 29404 15872 29408
rect 15808 29348 15812 29404
rect 15812 29348 15868 29404
rect 15868 29348 15872 29404
rect 15808 29344 15872 29348
rect 15888 29404 15952 29408
rect 15888 29348 15892 29404
rect 15892 29348 15948 29404
rect 15948 29348 15952 29404
rect 15888 29344 15952 29348
rect 15968 29404 16032 29408
rect 15968 29348 15972 29404
rect 15972 29348 16028 29404
rect 16028 29348 16032 29404
rect 15968 29344 16032 29348
rect 16048 29404 16112 29408
rect 16048 29348 16052 29404
rect 16052 29348 16108 29404
rect 16108 29348 16112 29404
rect 16048 29344 16112 29348
rect 23236 29404 23300 29408
rect 23236 29348 23240 29404
rect 23240 29348 23296 29404
rect 23296 29348 23300 29404
rect 23236 29344 23300 29348
rect 23316 29404 23380 29408
rect 23316 29348 23320 29404
rect 23320 29348 23376 29404
rect 23376 29348 23380 29404
rect 23316 29344 23380 29348
rect 23396 29404 23460 29408
rect 23396 29348 23400 29404
rect 23400 29348 23456 29404
rect 23456 29348 23460 29404
rect 23396 29344 23460 29348
rect 23476 29404 23540 29408
rect 23476 29348 23480 29404
rect 23480 29348 23536 29404
rect 23536 29348 23540 29404
rect 23476 29344 23540 29348
rect 30664 29404 30728 29408
rect 30664 29348 30668 29404
rect 30668 29348 30724 29404
rect 30724 29348 30728 29404
rect 30664 29344 30728 29348
rect 30744 29404 30808 29408
rect 30744 29348 30748 29404
rect 30748 29348 30804 29404
rect 30804 29348 30808 29404
rect 30744 29344 30808 29348
rect 30824 29404 30888 29408
rect 30824 29348 30828 29404
rect 30828 29348 30884 29404
rect 30884 29348 30888 29404
rect 30824 29344 30888 29348
rect 30904 29404 30968 29408
rect 30904 29348 30908 29404
rect 30908 29348 30964 29404
rect 30964 29348 30968 29404
rect 30904 29344 30968 29348
rect 4666 28860 4730 28864
rect 4666 28804 4670 28860
rect 4670 28804 4726 28860
rect 4726 28804 4730 28860
rect 4666 28800 4730 28804
rect 4746 28860 4810 28864
rect 4746 28804 4750 28860
rect 4750 28804 4806 28860
rect 4806 28804 4810 28860
rect 4746 28800 4810 28804
rect 4826 28860 4890 28864
rect 4826 28804 4830 28860
rect 4830 28804 4886 28860
rect 4886 28804 4890 28860
rect 4826 28800 4890 28804
rect 4906 28860 4970 28864
rect 4906 28804 4910 28860
rect 4910 28804 4966 28860
rect 4966 28804 4970 28860
rect 4906 28800 4970 28804
rect 12094 28860 12158 28864
rect 12094 28804 12098 28860
rect 12098 28804 12154 28860
rect 12154 28804 12158 28860
rect 12094 28800 12158 28804
rect 12174 28860 12238 28864
rect 12174 28804 12178 28860
rect 12178 28804 12234 28860
rect 12234 28804 12238 28860
rect 12174 28800 12238 28804
rect 12254 28860 12318 28864
rect 12254 28804 12258 28860
rect 12258 28804 12314 28860
rect 12314 28804 12318 28860
rect 12254 28800 12318 28804
rect 12334 28860 12398 28864
rect 12334 28804 12338 28860
rect 12338 28804 12394 28860
rect 12394 28804 12398 28860
rect 12334 28800 12398 28804
rect 19522 28860 19586 28864
rect 19522 28804 19526 28860
rect 19526 28804 19582 28860
rect 19582 28804 19586 28860
rect 19522 28800 19586 28804
rect 19602 28860 19666 28864
rect 19602 28804 19606 28860
rect 19606 28804 19662 28860
rect 19662 28804 19666 28860
rect 19602 28800 19666 28804
rect 19682 28860 19746 28864
rect 19682 28804 19686 28860
rect 19686 28804 19742 28860
rect 19742 28804 19746 28860
rect 19682 28800 19746 28804
rect 19762 28860 19826 28864
rect 19762 28804 19766 28860
rect 19766 28804 19822 28860
rect 19822 28804 19826 28860
rect 19762 28800 19826 28804
rect 26950 28860 27014 28864
rect 26950 28804 26954 28860
rect 26954 28804 27010 28860
rect 27010 28804 27014 28860
rect 26950 28800 27014 28804
rect 27030 28860 27094 28864
rect 27030 28804 27034 28860
rect 27034 28804 27090 28860
rect 27090 28804 27094 28860
rect 27030 28800 27094 28804
rect 27110 28860 27174 28864
rect 27110 28804 27114 28860
rect 27114 28804 27170 28860
rect 27170 28804 27174 28860
rect 27110 28800 27174 28804
rect 27190 28860 27254 28864
rect 27190 28804 27194 28860
rect 27194 28804 27250 28860
rect 27250 28804 27254 28860
rect 27190 28800 27254 28804
rect 8380 28316 8444 28320
rect 8380 28260 8384 28316
rect 8384 28260 8440 28316
rect 8440 28260 8444 28316
rect 8380 28256 8444 28260
rect 8460 28316 8524 28320
rect 8460 28260 8464 28316
rect 8464 28260 8520 28316
rect 8520 28260 8524 28316
rect 8460 28256 8524 28260
rect 8540 28316 8604 28320
rect 8540 28260 8544 28316
rect 8544 28260 8600 28316
rect 8600 28260 8604 28316
rect 8540 28256 8604 28260
rect 8620 28316 8684 28320
rect 8620 28260 8624 28316
rect 8624 28260 8680 28316
rect 8680 28260 8684 28316
rect 8620 28256 8684 28260
rect 15808 28316 15872 28320
rect 15808 28260 15812 28316
rect 15812 28260 15868 28316
rect 15868 28260 15872 28316
rect 15808 28256 15872 28260
rect 15888 28316 15952 28320
rect 15888 28260 15892 28316
rect 15892 28260 15948 28316
rect 15948 28260 15952 28316
rect 15888 28256 15952 28260
rect 15968 28316 16032 28320
rect 15968 28260 15972 28316
rect 15972 28260 16028 28316
rect 16028 28260 16032 28316
rect 15968 28256 16032 28260
rect 16048 28316 16112 28320
rect 16048 28260 16052 28316
rect 16052 28260 16108 28316
rect 16108 28260 16112 28316
rect 16048 28256 16112 28260
rect 23236 28316 23300 28320
rect 23236 28260 23240 28316
rect 23240 28260 23296 28316
rect 23296 28260 23300 28316
rect 23236 28256 23300 28260
rect 23316 28316 23380 28320
rect 23316 28260 23320 28316
rect 23320 28260 23376 28316
rect 23376 28260 23380 28316
rect 23316 28256 23380 28260
rect 23396 28316 23460 28320
rect 23396 28260 23400 28316
rect 23400 28260 23456 28316
rect 23456 28260 23460 28316
rect 23396 28256 23460 28260
rect 23476 28316 23540 28320
rect 23476 28260 23480 28316
rect 23480 28260 23536 28316
rect 23536 28260 23540 28316
rect 23476 28256 23540 28260
rect 30664 28316 30728 28320
rect 30664 28260 30668 28316
rect 30668 28260 30724 28316
rect 30724 28260 30728 28316
rect 30664 28256 30728 28260
rect 30744 28316 30808 28320
rect 30744 28260 30748 28316
rect 30748 28260 30804 28316
rect 30804 28260 30808 28316
rect 30744 28256 30808 28260
rect 30824 28316 30888 28320
rect 30824 28260 30828 28316
rect 30828 28260 30884 28316
rect 30884 28260 30888 28316
rect 30824 28256 30888 28260
rect 30904 28316 30968 28320
rect 30904 28260 30908 28316
rect 30908 28260 30964 28316
rect 30964 28260 30968 28316
rect 30904 28256 30968 28260
rect 4666 27772 4730 27776
rect 4666 27716 4670 27772
rect 4670 27716 4726 27772
rect 4726 27716 4730 27772
rect 4666 27712 4730 27716
rect 4746 27772 4810 27776
rect 4746 27716 4750 27772
rect 4750 27716 4806 27772
rect 4806 27716 4810 27772
rect 4746 27712 4810 27716
rect 4826 27772 4890 27776
rect 4826 27716 4830 27772
rect 4830 27716 4886 27772
rect 4886 27716 4890 27772
rect 4826 27712 4890 27716
rect 4906 27772 4970 27776
rect 4906 27716 4910 27772
rect 4910 27716 4966 27772
rect 4966 27716 4970 27772
rect 4906 27712 4970 27716
rect 12094 27772 12158 27776
rect 12094 27716 12098 27772
rect 12098 27716 12154 27772
rect 12154 27716 12158 27772
rect 12094 27712 12158 27716
rect 12174 27772 12238 27776
rect 12174 27716 12178 27772
rect 12178 27716 12234 27772
rect 12234 27716 12238 27772
rect 12174 27712 12238 27716
rect 12254 27772 12318 27776
rect 12254 27716 12258 27772
rect 12258 27716 12314 27772
rect 12314 27716 12318 27772
rect 12254 27712 12318 27716
rect 12334 27772 12398 27776
rect 12334 27716 12338 27772
rect 12338 27716 12394 27772
rect 12394 27716 12398 27772
rect 12334 27712 12398 27716
rect 19522 27772 19586 27776
rect 19522 27716 19526 27772
rect 19526 27716 19582 27772
rect 19582 27716 19586 27772
rect 19522 27712 19586 27716
rect 19602 27772 19666 27776
rect 19602 27716 19606 27772
rect 19606 27716 19662 27772
rect 19662 27716 19666 27772
rect 19602 27712 19666 27716
rect 19682 27772 19746 27776
rect 19682 27716 19686 27772
rect 19686 27716 19742 27772
rect 19742 27716 19746 27772
rect 19682 27712 19746 27716
rect 19762 27772 19826 27776
rect 19762 27716 19766 27772
rect 19766 27716 19822 27772
rect 19822 27716 19826 27772
rect 19762 27712 19826 27716
rect 26950 27772 27014 27776
rect 26950 27716 26954 27772
rect 26954 27716 27010 27772
rect 27010 27716 27014 27772
rect 26950 27712 27014 27716
rect 27030 27772 27094 27776
rect 27030 27716 27034 27772
rect 27034 27716 27090 27772
rect 27090 27716 27094 27772
rect 27030 27712 27094 27716
rect 27110 27772 27174 27776
rect 27110 27716 27114 27772
rect 27114 27716 27170 27772
rect 27170 27716 27174 27772
rect 27110 27712 27174 27716
rect 27190 27772 27254 27776
rect 27190 27716 27194 27772
rect 27194 27716 27250 27772
rect 27250 27716 27254 27772
rect 27190 27712 27254 27716
rect 8380 27228 8444 27232
rect 8380 27172 8384 27228
rect 8384 27172 8440 27228
rect 8440 27172 8444 27228
rect 8380 27168 8444 27172
rect 8460 27228 8524 27232
rect 8460 27172 8464 27228
rect 8464 27172 8520 27228
rect 8520 27172 8524 27228
rect 8460 27168 8524 27172
rect 8540 27228 8604 27232
rect 8540 27172 8544 27228
rect 8544 27172 8600 27228
rect 8600 27172 8604 27228
rect 8540 27168 8604 27172
rect 8620 27228 8684 27232
rect 8620 27172 8624 27228
rect 8624 27172 8680 27228
rect 8680 27172 8684 27228
rect 8620 27168 8684 27172
rect 15808 27228 15872 27232
rect 15808 27172 15812 27228
rect 15812 27172 15868 27228
rect 15868 27172 15872 27228
rect 15808 27168 15872 27172
rect 15888 27228 15952 27232
rect 15888 27172 15892 27228
rect 15892 27172 15948 27228
rect 15948 27172 15952 27228
rect 15888 27168 15952 27172
rect 15968 27228 16032 27232
rect 15968 27172 15972 27228
rect 15972 27172 16028 27228
rect 16028 27172 16032 27228
rect 15968 27168 16032 27172
rect 16048 27228 16112 27232
rect 16048 27172 16052 27228
rect 16052 27172 16108 27228
rect 16108 27172 16112 27228
rect 16048 27168 16112 27172
rect 23236 27228 23300 27232
rect 23236 27172 23240 27228
rect 23240 27172 23296 27228
rect 23296 27172 23300 27228
rect 23236 27168 23300 27172
rect 23316 27228 23380 27232
rect 23316 27172 23320 27228
rect 23320 27172 23376 27228
rect 23376 27172 23380 27228
rect 23316 27168 23380 27172
rect 23396 27228 23460 27232
rect 23396 27172 23400 27228
rect 23400 27172 23456 27228
rect 23456 27172 23460 27228
rect 23396 27168 23460 27172
rect 23476 27228 23540 27232
rect 23476 27172 23480 27228
rect 23480 27172 23536 27228
rect 23536 27172 23540 27228
rect 23476 27168 23540 27172
rect 30664 27228 30728 27232
rect 30664 27172 30668 27228
rect 30668 27172 30724 27228
rect 30724 27172 30728 27228
rect 30664 27168 30728 27172
rect 30744 27228 30808 27232
rect 30744 27172 30748 27228
rect 30748 27172 30804 27228
rect 30804 27172 30808 27228
rect 30744 27168 30808 27172
rect 30824 27228 30888 27232
rect 30824 27172 30828 27228
rect 30828 27172 30884 27228
rect 30884 27172 30888 27228
rect 30824 27168 30888 27172
rect 30904 27228 30968 27232
rect 30904 27172 30908 27228
rect 30908 27172 30964 27228
rect 30964 27172 30968 27228
rect 30904 27168 30968 27172
rect 4666 26684 4730 26688
rect 4666 26628 4670 26684
rect 4670 26628 4726 26684
rect 4726 26628 4730 26684
rect 4666 26624 4730 26628
rect 4746 26684 4810 26688
rect 4746 26628 4750 26684
rect 4750 26628 4806 26684
rect 4806 26628 4810 26684
rect 4746 26624 4810 26628
rect 4826 26684 4890 26688
rect 4826 26628 4830 26684
rect 4830 26628 4886 26684
rect 4886 26628 4890 26684
rect 4826 26624 4890 26628
rect 4906 26684 4970 26688
rect 4906 26628 4910 26684
rect 4910 26628 4966 26684
rect 4966 26628 4970 26684
rect 4906 26624 4970 26628
rect 12094 26684 12158 26688
rect 12094 26628 12098 26684
rect 12098 26628 12154 26684
rect 12154 26628 12158 26684
rect 12094 26624 12158 26628
rect 12174 26684 12238 26688
rect 12174 26628 12178 26684
rect 12178 26628 12234 26684
rect 12234 26628 12238 26684
rect 12174 26624 12238 26628
rect 12254 26684 12318 26688
rect 12254 26628 12258 26684
rect 12258 26628 12314 26684
rect 12314 26628 12318 26684
rect 12254 26624 12318 26628
rect 12334 26684 12398 26688
rect 12334 26628 12338 26684
rect 12338 26628 12394 26684
rect 12394 26628 12398 26684
rect 12334 26624 12398 26628
rect 19522 26684 19586 26688
rect 19522 26628 19526 26684
rect 19526 26628 19582 26684
rect 19582 26628 19586 26684
rect 19522 26624 19586 26628
rect 19602 26684 19666 26688
rect 19602 26628 19606 26684
rect 19606 26628 19662 26684
rect 19662 26628 19666 26684
rect 19602 26624 19666 26628
rect 19682 26684 19746 26688
rect 19682 26628 19686 26684
rect 19686 26628 19742 26684
rect 19742 26628 19746 26684
rect 19682 26624 19746 26628
rect 19762 26684 19826 26688
rect 19762 26628 19766 26684
rect 19766 26628 19822 26684
rect 19822 26628 19826 26684
rect 19762 26624 19826 26628
rect 26950 26684 27014 26688
rect 26950 26628 26954 26684
rect 26954 26628 27010 26684
rect 27010 26628 27014 26684
rect 26950 26624 27014 26628
rect 27030 26684 27094 26688
rect 27030 26628 27034 26684
rect 27034 26628 27090 26684
rect 27090 26628 27094 26684
rect 27030 26624 27094 26628
rect 27110 26684 27174 26688
rect 27110 26628 27114 26684
rect 27114 26628 27170 26684
rect 27170 26628 27174 26684
rect 27110 26624 27174 26628
rect 27190 26684 27254 26688
rect 27190 26628 27194 26684
rect 27194 26628 27250 26684
rect 27250 26628 27254 26684
rect 27190 26624 27254 26628
rect 8380 26140 8444 26144
rect 8380 26084 8384 26140
rect 8384 26084 8440 26140
rect 8440 26084 8444 26140
rect 8380 26080 8444 26084
rect 8460 26140 8524 26144
rect 8460 26084 8464 26140
rect 8464 26084 8520 26140
rect 8520 26084 8524 26140
rect 8460 26080 8524 26084
rect 8540 26140 8604 26144
rect 8540 26084 8544 26140
rect 8544 26084 8600 26140
rect 8600 26084 8604 26140
rect 8540 26080 8604 26084
rect 8620 26140 8684 26144
rect 8620 26084 8624 26140
rect 8624 26084 8680 26140
rect 8680 26084 8684 26140
rect 8620 26080 8684 26084
rect 15808 26140 15872 26144
rect 15808 26084 15812 26140
rect 15812 26084 15868 26140
rect 15868 26084 15872 26140
rect 15808 26080 15872 26084
rect 15888 26140 15952 26144
rect 15888 26084 15892 26140
rect 15892 26084 15948 26140
rect 15948 26084 15952 26140
rect 15888 26080 15952 26084
rect 15968 26140 16032 26144
rect 15968 26084 15972 26140
rect 15972 26084 16028 26140
rect 16028 26084 16032 26140
rect 15968 26080 16032 26084
rect 16048 26140 16112 26144
rect 16048 26084 16052 26140
rect 16052 26084 16108 26140
rect 16108 26084 16112 26140
rect 16048 26080 16112 26084
rect 23236 26140 23300 26144
rect 23236 26084 23240 26140
rect 23240 26084 23296 26140
rect 23296 26084 23300 26140
rect 23236 26080 23300 26084
rect 23316 26140 23380 26144
rect 23316 26084 23320 26140
rect 23320 26084 23376 26140
rect 23376 26084 23380 26140
rect 23316 26080 23380 26084
rect 23396 26140 23460 26144
rect 23396 26084 23400 26140
rect 23400 26084 23456 26140
rect 23456 26084 23460 26140
rect 23396 26080 23460 26084
rect 23476 26140 23540 26144
rect 23476 26084 23480 26140
rect 23480 26084 23536 26140
rect 23536 26084 23540 26140
rect 23476 26080 23540 26084
rect 30664 26140 30728 26144
rect 30664 26084 30668 26140
rect 30668 26084 30724 26140
rect 30724 26084 30728 26140
rect 30664 26080 30728 26084
rect 30744 26140 30808 26144
rect 30744 26084 30748 26140
rect 30748 26084 30804 26140
rect 30804 26084 30808 26140
rect 30744 26080 30808 26084
rect 30824 26140 30888 26144
rect 30824 26084 30828 26140
rect 30828 26084 30884 26140
rect 30884 26084 30888 26140
rect 30824 26080 30888 26084
rect 30904 26140 30968 26144
rect 30904 26084 30908 26140
rect 30908 26084 30964 26140
rect 30964 26084 30968 26140
rect 30904 26080 30968 26084
rect 4666 25596 4730 25600
rect 4666 25540 4670 25596
rect 4670 25540 4726 25596
rect 4726 25540 4730 25596
rect 4666 25536 4730 25540
rect 4746 25596 4810 25600
rect 4746 25540 4750 25596
rect 4750 25540 4806 25596
rect 4806 25540 4810 25596
rect 4746 25536 4810 25540
rect 4826 25596 4890 25600
rect 4826 25540 4830 25596
rect 4830 25540 4886 25596
rect 4886 25540 4890 25596
rect 4826 25536 4890 25540
rect 4906 25596 4970 25600
rect 4906 25540 4910 25596
rect 4910 25540 4966 25596
rect 4966 25540 4970 25596
rect 4906 25536 4970 25540
rect 12094 25596 12158 25600
rect 12094 25540 12098 25596
rect 12098 25540 12154 25596
rect 12154 25540 12158 25596
rect 12094 25536 12158 25540
rect 12174 25596 12238 25600
rect 12174 25540 12178 25596
rect 12178 25540 12234 25596
rect 12234 25540 12238 25596
rect 12174 25536 12238 25540
rect 12254 25596 12318 25600
rect 12254 25540 12258 25596
rect 12258 25540 12314 25596
rect 12314 25540 12318 25596
rect 12254 25536 12318 25540
rect 12334 25596 12398 25600
rect 12334 25540 12338 25596
rect 12338 25540 12394 25596
rect 12394 25540 12398 25596
rect 12334 25536 12398 25540
rect 19522 25596 19586 25600
rect 19522 25540 19526 25596
rect 19526 25540 19582 25596
rect 19582 25540 19586 25596
rect 19522 25536 19586 25540
rect 19602 25596 19666 25600
rect 19602 25540 19606 25596
rect 19606 25540 19662 25596
rect 19662 25540 19666 25596
rect 19602 25536 19666 25540
rect 19682 25596 19746 25600
rect 19682 25540 19686 25596
rect 19686 25540 19742 25596
rect 19742 25540 19746 25596
rect 19682 25536 19746 25540
rect 19762 25596 19826 25600
rect 19762 25540 19766 25596
rect 19766 25540 19822 25596
rect 19822 25540 19826 25596
rect 19762 25536 19826 25540
rect 26950 25596 27014 25600
rect 26950 25540 26954 25596
rect 26954 25540 27010 25596
rect 27010 25540 27014 25596
rect 26950 25536 27014 25540
rect 27030 25596 27094 25600
rect 27030 25540 27034 25596
rect 27034 25540 27090 25596
rect 27090 25540 27094 25596
rect 27030 25536 27094 25540
rect 27110 25596 27174 25600
rect 27110 25540 27114 25596
rect 27114 25540 27170 25596
rect 27170 25540 27174 25596
rect 27110 25536 27174 25540
rect 27190 25596 27254 25600
rect 27190 25540 27194 25596
rect 27194 25540 27250 25596
rect 27250 25540 27254 25596
rect 27190 25536 27254 25540
rect 8380 25052 8444 25056
rect 8380 24996 8384 25052
rect 8384 24996 8440 25052
rect 8440 24996 8444 25052
rect 8380 24992 8444 24996
rect 8460 25052 8524 25056
rect 8460 24996 8464 25052
rect 8464 24996 8520 25052
rect 8520 24996 8524 25052
rect 8460 24992 8524 24996
rect 8540 25052 8604 25056
rect 8540 24996 8544 25052
rect 8544 24996 8600 25052
rect 8600 24996 8604 25052
rect 8540 24992 8604 24996
rect 8620 25052 8684 25056
rect 8620 24996 8624 25052
rect 8624 24996 8680 25052
rect 8680 24996 8684 25052
rect 8620 24992 8684 24996
rect 15808 25052 15872 25056
rect 15808 24996 15812 25052
rect 15812 24996 15868 25052
rect 15868 24996 15872 25052
rect 15808 24992 15872 24996
rect 15888 25052 15952 25056
rect 15888 24996 15892 25052
rect 15892 24996 15948 25052
rect 15948 24996 15952 25052
rect 15888 24992 15952 24996
rect 15968 25052 16032 25056
rect 15968 24996 15972 25052
rect 15972 24996 16028 25052
rect 16028 24996 16032 25052
rect 15968 24992 16032 24996
rect 16048 25052 16112 25056
rect 16048 24996 16052 25052
rect 16052 24996 16108 25052
rect 16108 24996 16112 25052
rect 16048 24992 16112 24996
rect 23236 25052 23300 25056
rect 23236 24996 23240 25052
rect 23240 24996 23296 25052
rect 23296 24996 23300 25052
rect 23236 24992 23300 24996
rect 23316 25052 23380 25056
rect 23316 24996 23320 25052
rect 23320 24996 23376 25052
rect 23376 24996 23380 25052
rect 23316 24992 23380 24996
rect 23396 25052 23460 25056
rect 23396 24996 23400 25052
rect 23400 24996 23456 25052
rect 23456 24996 23460 25052
rect 23396 24992 23460 24996
rect 23476 25052 23540 25056
rect 23476 24996 23480 25052
rect 23480 24996 23536 25052
rect 23536 24996 23540 25052
rect 23476 24992 23540 24996
rect 30664 25052 30728 25056
rect 30664 24996 30668 25052
rect 30668 24996 30724 25052
rect 30724 24996 30728 25052
rect 30664 24992 30728 24996
rect 30744 25052 30808 25056
rect 30744 24996 30748 25052
rect 30748 24996 30804 25052
rect 30804 24996 30808 25052
rect 30744 24992 30808 24996
rect 30824 25052 30888 25056
rect 30824 24996 30828 25052
rect 30828 24996 30884 25052
rect 30884 24996 30888 25052
rect 30824 24992 30888 24996
rect 30904 25052 30968 25056
rect 30904 24996 30908 25052
rect 30908 24996 30964 25052
rect 30964 24996 30968 25052
rect 30904 24992 30968 24996
rect 4666 24508 4730 24512
rect 4666 24452 4670 24508
rect 4670 24452 4726 24508
rect 4726 24452 4730 24508
rect 4666 24448 4730 24452
rect 4746 24508 4810 24512
rect 4746 24452 4750 24508
rect 4750 24452 4806 24508
rect 4806 24452 4810 24508
rect 4746 24448 4810 24452
rect 4826 24508 4890 24512
rect 4826 24452 4830 24508
rect 4830 24452 4886 24508
rect 4886 24452 4890 24508
rect 4826 24448 4890 24452
rect 4906 24508 4970 24512
rect 4906 24452 4910 24508
rect 4910 24452 4966 24508
rect 4966 24452 4970 24508
rect 4906 24448 4970 24452
rect 12094 24508 12158 24512
rect 12094 24452 12098 24508
rect 12098 24452 12154 24508
rect 12154 24452 12158 24508
rect 12094 24448 12158 24452
rect 12174 24508 12238 24512
rect 12174 24452 12178 24508
rect 12178 24452 12234 24508
rect 12234 24452 12238 24508
rect 12174 24448 12238 24452
rect 12254 24508 12318 24512
rect 12254 24452 12258 24508
rect 12258 24452 12314 24508
rect 12314 24452 12318 24508
rect 12254 24448 12318 24452
rect 12334 24508 12398 24512
rect 12334 24452 12338 24508
rect 12338 24452 12394 24508
rect 12394 24452 12398 24508
rect 12334 24448 12398 24452
rect 19522 24508 19586 24512
rect 19522 24452 19526 24508
rect 19526 24452 19582 24508
rect 19582 24452 19586 24508
rect 19522 24448 19586 24452
rect 19602 24508 19666 24512
rect 19602 24452 19606 24508
rect 19606 24452 19662 24508
rect 19662 24452 19666 24508
rect 19602 24448 19666 24452
rect 19682 24508 19746 24512
rect 19682 24452 19686 24508
rect 19686 24452 19742 24508
rect 19742 24452 19746 24508
rect 19682 24448 19746 24452
rect 19762 24508 19826 24512
rect 19762 24452 19766 24508
rect 19766 24452 19822 24508
rect 19822 24452 19826 24508
rect 19762 24448 19826 24452
rect 26950 24508 27014 24512
rect 26950 24452 26954 24508
rect 26954 24452 27010 24508
rect 27010 24452 27014 24508
rect 26950 24448 27014 24452
rect 27030 24508 27094 24512
rect 27030 24452 27034 24508
rect 27034 24452 27090 24508
rect 27090 24452 27094 24508
rect 27030 24448 27094 24452
rect 27110 24508 27174 24512
rect 27110 24452 27114 24508
rect 27114 24452 27170 24508
rect 27170 24452 27174 24508
rect 27110 24448 27174 24452
rect 27190 24508 27254 24512
rect 27190 24452 27194 24508
rect 27194 24452 27250 24508
rect 27250 24452 27254 24508
rect 27190 24448 27254 24452
rect 8380 23964 8444 23968
rect 8380 23908 8384 23964
rect 8384 23908 8440 23964
rect 8440 23908 8444 23964
rect 8380 23904 8444 23908
rect 8460 23964 8524 23968
rect 8460 23908 8464 23964
rect 8464 23908 8520 23964
rect 8520 23908 8524 23964
rect 8460 23904 8524 23908
rect 8540 23964 8604 23968
rect 8540 23908 8544 23964
rect 8544 23908 8600 23964
rect 8600 23908 8604 23964
rect 8540 23904 8604 23908
rect 8620 23964 8684 23968
rect 8620 23908 8624 23964
rect 8624 23908 8680 23964
rect 8680 23908 8684 23964
rect 8620 23904 8684 23908
rect 15808 23964 15872 23968
rect 15808 23908 15812 23964
rect 15812 23908 15868 23964
rect 15868 23908 15872 23964
rect 15808 23904 15872 23908
rect 15888 23964 15952 23968
rect 15888 23908 15892 23964
rect 15892 23908 15948 23964
rect 15948 23908 15952 23964
rect 15888 23904 15952 23908
rect 15968 23964 16032 23968
rect 15968 23908 15972 23964
rect 15972 23908 16028 23964
rect 16028 23908 16032 23964
rect 15968 23904 16032 23908
rect 16048 23964 16112 23968
rect 16048 23908 16052 23964
rect 16052 23908 16108 23964
rect 16108 23908 16112 23964
rect 16048 23904 16112 23908
rect 23236 23964 23300 23968
rect 23236 23908 23240 23964
rect 23240 23908 23296 23964
rect 23296 23908 23300 23964
rect 23236 23904 23300 23908
rect 23316 23964 23380 23968
rect 23316 23908 23320 23964
rect 23320 23908 23376 23964
rect 23376 23908 23380 23964
rect 23316 23904 23380 23908
rect 23396 23964 23460 23968
rect 23396 23908 23400 23964
rect 23400 23908 23456 23964
rect 23456 23908 23460 23964
rect 23396 23904 23460 23908
rect 23476 23964 23540 23968
rect 23476 23908 23480 23964
rect 23480 23908 23536 23964
rect 23536 23908 23540 23964
rect 23476 23904 23540 23908
rect 30664 23964 30728 23968
rect 30664 23908 30668 23964
rect 30668 23908 30724 23964
rect 30724 23908 30728 23964
rect 30664 23904 30728 23908
rect 30744 23964 30808 23968
rect 30744 23908 30748 23964
rect 30748 23908 30804 23964
rect 30804 23908 30808 23964
rect 30744 23904 30808 23908
rect 30824 23964 30888 23968
rect 30824 23908 30828 23964
rect 30828 23908 30884 23964
rect 30884 23908 30888 23964
rect 30824 23904 30888 23908
rect 30904 23964 30968 23968
rect 30904 23908 30908 23964
rect 30908 23908 30964 23964
rect 30964 23908 30968 23964
rect 30904 23904 30968 23908
rect 4666 23420 4730 23424
rect 4666 23364 4670 23420
rect 4670 23364 4726 23420
rect 4726 23364 4730 23420
rect 4666 23360 4730 23364
rect 4746 23420 4810 23424
rect 4746 23364 4750 23420
rect 4750 23364 4806 23420
rect 4806 23364 4810 23420
rect 4746 23360 4810 23364
rect 4826 23420 4890 23424
rect 4826 23364 4830 23420
rect 4830 23364 4886 23420
rect 4886 23364 4890 23420
rect 4826 23360 4890 23364
rect 4906 23420 4970 23424
rect 4906 23364 4910 23420
rect 4910 23364 4966 23420
rect 4966 23364 4970 23420
rect 4906 23360 4970 23364
rect 12094 23420 12158 23424
rect 12094 23364 12098 23420
rect 12098 23364 12154 23420
rect 12154 23364 12158 23420
rect 12094 23360 12158 23364
rect 12174 23420 12238 23424
rect 12174 23364 12178 23420
rect 12178 23364 12234 23420
rect 12234 23364 12238 23420
rect 12174 23360 12238 23364
rect 12254 23420 12318 23424
rect 12254 23364 12258 23420
rect 12258 23364 12314 23420
rect 12314 23364 12318 23420
rect 12254 23360 12318 23364
rect 12334 23420 12398 23424
rect 12334 23364 12338 23420
rect 12338 23364 12394 23420
rect 12394 23364 12398 23420
rect 12334 23360 12398 23364
rect 19522 23420 19586 23424
rect 19522 23364 19526 23420
rect 19526 23364 19582 23420
rect 19582 23364 19586 23420
rect 19522 23360 19586 23364
rect 19602 23420 19666 23424
rect 19602 23364 19606 23420
rect 19606 23364 19662 23420
rect 19662 23364 19666 23420
rect 19602 23360 19666 23364
rect 19682 23420 19746 23424
rect 19682 23364 19686 23420
rect 19686 23364 19742 23420
rect 19742 23364 19746 23420
rect 19682 23360 19746 23364
rect 19762 23420 19826 23424
rect 19762 23364 19766 23420
rect 19766 23364 19822 23420
rect 19822 23364 19826 23420
rect 19762 23360 19826 23364
rect 26950 23420 27014 23424
rect 26950 23364 26954 23420
rect 26954 23364 27010 23420
rect 27010 23364 27014 23420
rect 26950 23360 27014 23364
rect 27030 23420 27094 23424
rect 27030 23364 27034 23420
rect 27034 23364 27090 23420
rect 27090 23364 27094 23420
rect 27030 23360 27094 23364
rect 27110 23420 27174 23424
rect 27110 23364 27114 23420
rect 27114 23364 27170 23420
rect 27170 23364 27174 23420
rect 27110 23360 27174 23364
rect 27190 23420 27254 23424
rect 27190 23364 27194 23420
rect 27194 23364 27250 23420
rect 27250 23364 27254 23420
rect 27190 23360 27254 23364
rect 8380 22876 8444 22880
rect 8380 22820 8384 22876
rect 8384 22820 8440 22876
rect 8440 22820 8444 22876
rect 8380 22816 8444 22820
rect 8460 22876 8524 22880
rect 8460 22820 8464 22876
rect 8464 22820 8520 22876
rect 8520 22820 8524 22876
rect 8460 22816 8524 22820
rect 8540 22876 8604 22880
rect 8540 22820 8544 22876
rect 8544 22820 8600 22876
rect 8600 22820 8604 22876
rect 8540 22816 8604 22820
rect 8620 22876 8684 22880
rect 8620 22820 8624 22876
rect 8624 22820 8680 22876
rect 8680 22820 8684 22876
rect 8620 22816 8684 22820
rect 15808 22876 15872 22880
rect 15808 22820 15812 22876
rect 15812 22820 15868 22876
rect 15868 22820 15872 22876
rect 15808 22816 15872 22820
rect 15888 22876 15952 22880
rect 15888 22820 15892 22876
rect 15892 22820 15948 22876
rect 15948 22820 15952 22876
rect 15888 22816 15952 22820
rect 15968 22876 16032 22880
rect 15968 22820 15972 22876
rect 15972 22820 16028 22876
rect 16028 22820 16032 22876
rect 15968 22816 16032 22820
rect 16048 22876 16112 22880
rect 16048 22820 16052 22876
rect 16052 22820 16108 22876
rect 16108 22820 16112 22876
rect 16048 22816 16112 22820
rect 23236 22876 23300 22880
rect 23236 22820 23240 22876
rect 23240 22820 23296 22876
rect 23296 22820 23300 22876
rect 23236 22816 23300 22820
rect 23316 22876 23380 22880
rect 23316 22820 23320 22876
rect 23320 22820 23376 22876
rect 23376 22820 23380 22876
rect 23316 22816 23380 22820
rect 23396 22876 23460 22880
rect 23396 22820 23400 22876
rect 23400 22820 23456 22876
rect 23456 22820 23460 22876
rect 23396 22816 23460 22820
rect 23476 22876 23540 22880
rect 23476 22820 23480 22876
rect 23480 22820 23536 22876
rect 23536 22820 23540 22876
rect 23476 22816 23540 22820
rect 30664 22876 30728 22880
rect 30664 22820 30668 22876
rect 30668 22820 30724 22876
rect 30724 22820 30728 22876
rect 30664 22816 30728 22820
rect 30744 22876 30808 22880
rect 30744 22820 30748 22876
rect 30748 22820 30804 22876
rect 30804 22820 30808 22876
rect 30744 22816 30808 22820
rect 30824 22876 30888 22880
rect 30824 22820 30828 22876
rect 30828 22820 30884 22876
rect 30884 22820 30888 22876
rect 30824 22816 30888 22820
rect 30904 22876 30968 22880
rect 30904 22820 30908 22876
rect 30908 22820 30964 22876
rect 30964 22820 30968 22876
rect 30904 22816 30968 22820
rect 4666 22332 4730 22336
rect 4666 22276 4670 22332
rect 4670 22276 4726 22332
rect 4726 22276 4730 22332
rect 4666 22272 4730 22276
rect 4746 22332 4810 22336
rect 4746 22276 4750 22332
rect 4750 22276 4806 22332
rect 4806 22276 4810 22332
rect 4746 22272 4810 22276
rect 4826 22332 4890 22336
rect 4826 22276 4830 22332
rect 4830 22276 4886 22332
rect 4886 22276 4890 22332
rect 4826 22272 4890 22276
rect 4906 22332 4970 22336
rect 4906 22276 4910 22332
rect 4910 22276 4966 22332
rect 4966 22276 4970 22332
rect 4906 22272 4970 22276
rect 12094 22332 12158 22336
rect 12094 22276 12098 22332
rect 12098 22276 12154 22332
rect 12154 22276 12158 22332
rect 12094 22272 12158 22276
rect 12174 22332 12238 22336
rect 12174 22276 12178 22332
rect 12178 22276 12234 22332
rect 12234 22276 12238 22332
rect 12174 22272 12238 22276
rect 12254 22332 12318 22336
rect 12254 22276 12258 22332
rect 12258 22276 12314 22332
rect 12314 22276 12318 22332
rect 12254 22272 12318 22276
rect 12334 22332 12398 22336
rect 12334 22276 12338 22332
rect 12338 22276 12394 22332
rect 12394 22276 12398 22332
rect 12334 22272 12398 22276
rect 19522 22332 19586 22336
rect 19522 22276 19526 22332
rect 19526 22276 19582 22332
rect 19582 22276 19586 22332
rect 19522 22272 19586 22276
rect 19602 22332 19666 22336
rect 19602 22276 19606 22332
rect 19606 22276 19662 22332
rect 19662 22276 19666 22332
rect 19602 22272 19666 22276
rect 19682 22332 19746 22336
rect 19682 22276 19686 22332
rect 19686 22276 19742 22332
rect 19742 22276 19746 22332
rect 19682 22272 19746 22276
rect 19762 22332 19826 22336
rect 19762 22276 19766 22332
rect 19766 22276 19822 22332
rect 19822 22276 19826 22332
rect 19762 22272 19826 22276
rect 26950 22332 27014 22336
rect 26950 22276 26954 22332
rect 26954 22276 27010 22332
rect 27010 22276 27014 22332
rect 26950 22272 27014 22276
rect 27030 22332 27094 22336
rect 27030 22276 27034 22332
rect 27034 22276 27090 22332
rect 27090 22276 27094 22332
rect 27030 22272 27094 22276
rect 27110 22332 27174 22336
rect 27110 22276 27114 22332
rect 27114 22276 27170 22332
rect 27170 22276 27174 22332
rect 27110 22272 27174 22276
rect 27190 22332 27254 22336
rect 27190 22276 27194 22332
rect 27194 22276 27250 22332
rect 27250 22276 27254 22332
rect 27190 22272 27254 22276
rect 8380 21788 8444 21792
rect 8380 21732 8384 21788
rect 8384 21732 8440 21788
rect 8440 21732 8444 21788
rect 8380 21728 8444 21732
rect 8460 21788 8524 21792
rect 8460 21732 8464 21788
rect 8464 21732 8520 21788
rect 8520 21732 8524 21788
rect 8460 21728 8524 21732
rect 8540 21788 8604 21792
rect 8540 21732 8544 21788
rect 8544 21732 8600 21788
rect 8600 21732 8604 21788
rect 8540 21728 8604 21732
rect 8620 21788 8684 21792
rect 8620 21732 8624 21788
rect 8624 21732 8680 21788
rect 8680 21732 8684 21788
rect 8620 21728 8684 21732
rect 15808 21788 15872 21792
rect 15808 21732 15812 21788
rect 15812 21732 15868 21788
rect 15868 21732 15872 21788
rect 15808 21728 15872 21732
rect 15888 21788 15952 21792
rect 15888 21732 15892 21788
rect 15892 21732 15948 21788
rect 15948 21732 15952 21788
rect 15888 21728 15952 21732
rect 15968 21788 16032 21792
rect 15968 21732 15972 21788
rect 15972 21732 16028 21788
rect 16028 21732 16032 21788
rect 15968 21728 16032 21732
rect 16048 21788 16112 21792
rect 16048 21732 16052 21788
rect 16052 21732 16108 21788
rect 16108 21732 16112 21788
rect 16048 21728 16112 21732
rect 23236 21788 23300 21792
rect 23236 21732 23240 21788
rect 23240 21732 23296 21788
rect 23296 21732 23300 21788
rect 23236 21728 23300 21732
rect 23316 21788 23380 21792
rect 23316 21732 23320 21788
rect 23320 21732 23376 21788
rect 23376 21732 23380 21788
rect 23316 21728 23380 21732
rect 23396 21788 23460 21792
rect 23396 21732 23400 21788
rect 23400 21732 23456 21788
rect 23456 21732 23460 21788
rect 23396 21728 23460 21732
rect 23476 21788 23540 21792
rect 23476 21732 23480 21788
rect 23480 21732 23536 21788
rect 23536 21732 23540 21788
rect 23476 21728 23540 21732
rect 30664 21788 30728 21792
rect 30664 21732 30668 21788
rect 30668 21732 30724 21788
rect 30724 21732 30728 21788
rect 30664 21728 30728 21732
rect 30744 21788 30808 21792
rect 30744 21732 30748 21788
rect 30748 21732 30804 21788
rect 30804 21732 30808 21788
rect 30744 21728 30808 21732
rect 30824 21788 30888 21792
rect 30824 21732 30828 21788
rect 30828 21732 30884 21788
rect 30884 21732 30888 21788
rect 30824 21728 30888 21732
rect 30904 21788 30968 21792
rect 30904 21732 30908 21788
rect 30908 21732 30964 21788
rect 30964 21732 30968 21788
rect 30904 21728 30968 21732
rect 4666 21244 4730 21248
rect 4666 21188 4670 21244
rect 4670 21188 4726 21244
rect 4726 21188 4730 21244
rect 4666 21184 4730 21188
rect 4746 21244 4810 21248
rect 4746 21188 4750 21244
rect 4750 21188 4806 21244
rect 4806 21188 4810 21244
rect 4746 21184 4810 21188
rect 4826 21244 4890 21248
rect 4826 21188 4830 21244
rect 4830 21188 4886 21244
rect 4886 21188 4890 21244
rect 4826 21184 4890 21188
rect 4906 21244 4970 21248
rect 4906 21188 4910 21244
rect 4910 21188 4966 21244
rect 4966 21188 4970 21244
rect 4906 21184 4970 21188
rect 12094 21244 12158 21248
rect 12094 21188 12098 21244
rect 12098 21188 12154 21244
rect 12154 21188 12158 21244
rect 12094 21184 12158 21188
rect 12174 21244 12238 21248
rect 12174 21188 12178 21244
rect 12178 21188 12234 21244
rect 12234 21188 12238 21244
rect 12174 21184 12238 21188
rect 12254 21244 12318 21248
rect 12254 21188 12258 21244
rect 12258 21188 12314 21244
rect 12314 21188 12318 21244
rect 12254 21184 12318 21188
rect 12334 21244 12398 21248
rect 12334 21188 12338 21244
rect 12338 21188 12394 21244
rect 12394 21188 12398 21244
rect 12334 21184 12398 21188
rect 19522 21244 19586 21248
rect 19522 21188 19526 21244
rect 19526 21188 19582 21244
rect 19582 21188 19586 21244
rect 19522 21184 19586 21188
rect 19602 21244 19666 21248
rect 19602 21188 19606 21244
rect 19606 21188 19662 21244
rect 19662 21188 19666 21244
rect 19602 21184 19666 21188
rect 19682 21244 19746 21248
rect 19682 21188 19686 21244
rect 19686 21188 19742 21244
rect 19742 21188 19746 21244
rect 19682 21184 19746 21188
rect 19762 21244 19826 21248
rect 19762 21188 19766 21244
rect 19766 21188 19822 21244
rect 19822 21188 19826 21244
rect 19762 21184 19826 21188
rect 26950 21244 27014 21248
rect 26950 21188 26954 21244
rect 26954 21188 27010 21244
rect 27010 21188 27014 21244
rect 26950 21184 27014 21188
rect 27030 21244 27094 21248
rect 27030 21188 27034 21244
rect 27034 21188 27090 21244
rect 27090 21188 27094 21244
rect 27030 21184 27094 21188
rect 27110 21244 27174 21248
rect 27110 21188 27114 21244
rect 27114 21188 27170 21244
rect 27170 21188 27174 21244
rect 27110 21184 27174 21188
rect 27190 21244 27254 21248
rect 27190 21188 27194 21244
rect 27194 21188 27250 21244
rect 27250 21188 27254 21244
rect 27190 21184 27254 21188
rect 8380 20700 8444 20704
rect 8380 20644 8384 20700
rect 8384 20644 8440 20700
rect 8440 20644 8444 20700
rect 8380 20640 8444 20644
rect 8460 20700 8524 20704
rect 8460 20644 8464 20700
rect 8464 20644 8520 20700
rect 8520 20644 8524 20700
rect 8460 20640 8524 20644
rect 8540 20700 8604 20704
rect 8540 20644 8544 20700
rect 8544 20644 8600 20700
rect 8600 20644 8604 20700
rect 8540 20640 8604 20644
rect 8620 20700 8684 20704
rect 8620 20644 8624 20700
rect 8624 20644 8680 20700
rect 8680 20644 8684 20700
rect 8620 20640 8684 20644
rect 15808 20700 15872 20704
rect 15808 20644 15812 20700
rect 15812 20644 15868 20700
rect 15868 20644 15872 20700
rect 15808 20640 15872 20644
rect 15888 20700 15952 20704
rect 15888 20644 15892 20700
rect 15892 20644 15948 20700
rect 15948 20644 15952 20700
rect 15888 20640 15952 20644
rect 15968 20700 16032 20704
rect 15968 20644 15972 20700
rect 15972 20644 16028 20700
rect 16028 20644 16032 20700
rect 15968 20640 16032 20644
rect 16048 20700 16112 20704
rect 16048 20644 16052 20700
rect 16052 20644 16108 20700
rect 16108 20644 16112 20700
rect 16048 20640 16112 20644
rect 23236 20700 23300 20704
rect 23236 20644 23240 20700
rect 23240 20644 23296 20700
rect 23296 20644 23300 20700
rect 23236 20640 23300 20644
rect 23316 20700 23380 20704
rect 23316 20644 23320 20700
rect 23320 20644 23376 20700
rect 23376 20644 23380 20700
rect 23316 20640 23380 20644
rect 23396 20700 23460 20704
rect 23396 20644 23400 20700
rect 23400 20644 23456 20700
rect 23456 20644 23460 20700
rect 23396 20640 23460 20644
rect 23476 20700 23540 20704
rect 23476 20644 23480 20700
rect 23480 20644 23536 20700
rect 23536 20644 23540 20700
rect 23476 20640 23540 20644
rect 30664 20700 30728 20704
rect 30664 20644 30668 20700
rect 30668 20644 30724 20700
rect 30724 20644 30728 20700
rect 30664 20640 30728 20644
rect 30744 20700 30808 20704
rect 30744 20644 30748 20700
rect 30748 20644 30804 20700
rect 30804 20644 30808 20700
rect 30744 20640 30808 20644
rect 30824 20700 30888 20704
rect 30824 20644 30828 20700
rect 30828 20644 30884 20700
rect 30884 20644 30888 20700
rect 30824 20640 30888 20644
rect 30904 20700 30968 20704
rect 30904 20644 30908 20700
rect 30908 20644 30964 20700
rect 30964 20644 30968 20700
rect 30904 20640 30968 20644
rect 4666 20156 4730 20160
rect 4666 20100 4670 20156
rect 4670 20100 4726 20156
rect 4726 20100 4730 20156
rect 4666 20096 4730 20100
rect 4746 20156 4810 20160
rect 4746 20100 4750 20156
rect 4750 20100 4806 20156
rect 4806 20100 4810 20156
rect 4746 20096 4810 20100
rect 4826 20156 4890 20160
rect 4826 20100 4830 20156
rect 4830 20100 4886 20156
rect 4886 20100 4890 20156
rect 4826 20096 4890 20100
rect 4906 20156 4970 20160
rect 4906 20100 4910 20156
rect 4910 20100 4966 20156
rect 4966 20100 4970 20156
rect 4906 20096 4970 20100
rect 12094 20156 12158 20160
rect 12094 20100 12098 20156
rect 12098 20100 12154 20156
rect 12154 20100 12158 20156
rect 12094 20096 12158 20100
rect 12174 20156 12238 20160
rect 12174 20100 12178 20156
rect 12178 20100 12234 20156
rect 12234 20100 12238 20156
rect 12174 20096 12238 20100
rect 12254 20156 12318 20160
rect 12254 20100 12258 20156
rect 12258 20100 12314 20156
rect 12314 20100 12318 20156
rect 12254 20096 12318 20100
rect 12334 20156 12398 20160
rect 12334 20100 12338 20156
rect 12338 20100 12394 20156
rect 12394 20100 12398 20156
rect 12334 20096 12398 20100
rect 19522 20156 19586 20160
rect 19522 20100 19526 20156
rect 19526 20100 19582 20156
rect 19582 20100 19586 20156
rect 19522 20096 19586 20100
rect 19602 20156 19666 20160
rect 19602 20100 19606 20156
rect 19606 20100 19662 20156
rect 19662 20100 19666 20156
rect 19602 20096 19666 20100
rect 19682 20156 19746 20160
rect 19682 20100 19686 20156
rect 19686 20100 19742 20156
rect 19742 20100 19746 20156
rect 19682 20096 19746 20100
rect 19762 20156 19826 20160
rect 19762 20100 19766 20156
rect 19766 20100 19822 20156
rect 19822 20100 19826 20156
rect 19762 20096 19826 20100
rect 26950 20156 27014 20160
rect 26950 20100 26954 20156
rect 26954 20100 27010 20156
rect 27010 20100 27014 20156
rect 26950 20096 27014 20100
rect 27030 20156 27094 20160
rect 27030 20100 27034 20156
rect 27034 20100 27090 20156
rect 27090 20100 27094 20156
rect 27030 20096 27094 20100
rect 27110 20156 27174 20160
rect 27110 20100 27114 20156
rect 27114 20100 27170 20156
rect 27170 20100 27174 20156
rect 27110 20096 27174 20100
rect 27190 20156 27254 20160
rect 27190 20100 27194 20156
rect 27194 20100 27250 20156
rect 27250 20100 27254 20156
rect 27190 20096 27254 20100
rect 8380 19612 8444 19616
rect 8380 19556 8384 19612
rect 8384 19556 8440 19612
rect 8440 19556 8444 19612
rect 8380 19552 8444 19556
rect 8460 19612 8524 19616
rect 8460 19556 8464 19612
rect 8464 19556 8520 19612
rect 8520 19556 8524 19612
rect 8460 19552 8524 19556
rect 8540 19612 8604 19616
rect 8540 19556 8544 19612
rect 8544 19556 8600 19612
rect 8600 19556 8604 19612
rect 8540 19552 8604 19556
rect 8620 19612 8684 19616
rect 8620 19556 8624 19612
rect 8624 19556 8680 19612
rect 8680 19556 8684 19612
rect 8620 19552 8684 19556
rect 15808 19612 15872 19616
rect 15808 19556 15812 19612
rect 15812 19556 15868 19612
rect 15868 19556 15872 19612
rect 15808 19552 15872 19556
rect 15888 19612 15952 19616
rect 15888 19556 15892 19612
rect 15892 19556 15948 19612
rect 15948 19556 15952 19612
rect 15888 19552 15952 19556
rect 15968 19612 16032 19616
rect 15968 19556 15972 19612
rect 15972 19556 16028 19612
rect 16028 19556 16032 19612
rect 15968 19552 16032 19556
rect 16048 19612 16112 19616
rect 16048 19556 16052 19612
rect 16052 19556 16108 19612
rect 16108 19556 16112 19612
rect 16048 19552 16112 19556
rect 23236 19612 23300 19616
rect 23236 19556 23240 19612
rect 23240 19556 23296 19612
rect 23296 19556 23300 19612
rect 23236 19552 23300 19556
rect 23316 19612 23380 19616
rect 23316 19556 23320 19612
rect 23320 19556 23376 19612
rect 23376 19556 23380 19612
rect 23316 19552 23380 19556
rect 23396 19612 23460 19616
rect 23396 19556 23400 19612
rect 23400 19556 23456 19612
rect 23456 19556 23460 19612
rect 23396 19552 23460 19556
rect 23476 19612 23540 19616
rect 23476 19556 23480 19612
rect 23480 19556 23536 19612
rect 23536 19556 23540 19612
rect 23476 19552 23540 19556
rect 30664 19612 30728 19616
rect 30664 19556 30668 19612
rect 30668 19556 30724 19612
rect 30724 19556 30728 19612
rect 30664 19552 30728 19556
rect 30744 19612 30808 19616
rect 30744 19556 30748 19612
rect 30748 19556 30804 19612
rect 30804 19556 30808 19612
rect 30744 19552 30808 19556
rect 30824 19612 30888 19616
rect 30824 19556 30828 19612
rect 30828 19556 30884 19612
rect 30884 19556 30888 19612
rect 30824 19552 30888 19556
rect 30904 19612 30968 19616
rect 30904 19556 30908 19612
rect 30908 19556 30964 19612
rect 30964 19556 30968 19612
rect 30904 19552 30968 19556
rect 4666 19068 4730 19072
rect 4666 19012 4670 19068
rect 4670 19012 4726 19068
rect 4726 19012 4730 19068
rect 4666 19008 4730 19012
rect 4746 19068 4810 19072
rect 4746 19012 4750 19068
rect 4750 19012 4806 19068
rect 4806 19012 4810 19068
rect 4746 19008 4810 19012
rect 4826 19068 4890 19072
rect 4826 19012 4830 19068
rect 4830 19012 4886 19068
rect 4886 19012 4890 19068
rect 4826 19008 4890 19012
rect 4906 19068 4970 19072
rect 4906 19012 4910 19068
rect 4910 19012 4966 19068
rect 4966 19012 4970 19068
rect 4906 19008 4970 19012
rect 12094 19068 12158 19072
rect 12094 19012 12098 19068
rect 12098 19012 12154 19068
rect 12154 19012 12158 19068
rect 12094 19008 12158 19012
rect 12174 19068 12238 19072
rect 12174 19012 12178 19068
rect 12178 19012 12234 19068
rect 12234 19012 12238 19068
rect 12174 19008 12238 19012
rect 12254 19068 12318 19072
rect 12254 19012 12258 19068
rect 12258 19012 12314 19068
rect 12314 19012 12318 19068
rect 12254 19008 12318 19012
rect 12334 19068 12398 19072
rect 12334 19012 12338 19068
rect 12338 19012 12394 19068
rect 12394 19012 12398 19068
rect 12334 19008 12398 19012
rect 19522 19068 19586 19072
rect 19522 19012 19526 19068
rect 19526 19012 19582 19068
rect 19582 19012 19586 19068
rect 19522 19008 19586 19012
rect 19602 19068 19666 19072
rect 19602 19012 19606 19068
rect 19606 19012 19662 19068
rect 19662 19012 19666 19068
rect 19602 19008 19666 19012
rect 19682 19068 19746 19072
rect 19682 19012 19686 19068
rect 19686 19012 19742 19068
rect 19742 19012 19746 19068
rect 19682 19008 19746 19012
rect 19762 19068 19826 19072
rect 19762 19012 19766 19068
rect 19766 19012 19822 19068
rect 19822 19012 19826 19068
rect 19762 19008 19826 19012
rect 26950 19068 27014 19072
rect 26950 19012 26954 19068
rect 26954 19012 27010 19068
rect 27010 19012 27014 19068
rect 26950 19008 27014 19012
rect 27030 19068 27094 19072
rect 27030 19012 27034 19068
rect 27034 19012 27090 19068
rect 27090 19012 27094 19068
rect 27030 19008 27094 19012
rect 27110 19068 27174 19072
rect 27110 19012 27114 19068
rect 27114 19012 27170 19068
rect 27170 19012 27174 19068
rect 27110 19008 27174 19012
rect 27190 19068 27254 19072
rect 27190 19012 27194 19068
rect 27194 19012 27250 19068
rect 27250 19012 27254 19068
rect 27190 19008 27254 19012
rect 8380 18524 8444 18528
rect 8380 18468 8384 18524
rect 8384 18468 8440 18524
rect 8440 18468 8444 18524
rect 8380 18464 8444 18468
rect 8460 18524 8524 18528
rect 8460 18468 8464 18524
rect 8464 18468 8520 18524
rect 8520 18468 8524 18524
rect 8460 18464 8524 18468
rect 8540 18524 8604 18528
rect 8540 18468 8544 18524
rect 8544 18468 8600 18524
rect 8600 18468 8604 18524
rect 8540 18464 8604 18468
rect 8620 18524 8684 18528
rect 8620 18468 8624 18524
rect 8624 18468 8680 18524
rect 8680 18468 8684 18524
rect 8620 18464 8684 18468
rect 15808 18524 15872 18528
rect 15808 18468 15812 18524
rect 15812 18468 15868 18524
rect 15868 18468 15872 18524
rect 15808 18464 15872 18468
rect 15888 18524 15952 18528
rect 15888 18468 15892 18524
rect 15892 18468 15948 18524
rect 15948 18468 15952 18524
rect 15888 18464 15952 18468
rect 15968 18524 16032 18528
rect 15968 18468 15972 18524
rect 15972 18468 16028 18524
rect 16028 18468 16032 18524
rect 15968 18464 16032 18468
rect 16048 18524 16112 18528
rect 16048 18468 16052 18524
rect 16052 18468 16108 18524
rect 16108 18468 16112 18524
rect 16048 18464 16112 18468
rect 23236 18524 23300 18528
rect 23236 18468 23240 18524
rect 23240 18468 23296 18524
rect 23296 18468 23300 18524
rect 23236 18464 23300 18468
rect 23316 18524 23380 18528
rect 23316 18468 23320 18524
rect 23320 18468 23376 18524
rect 23376 18468 23380 18524
rect 23316 18464 23380 18468
rect 23396 18524 23460 18528
rect 23396 18468 23400 18524
rect 23400 18468 23456 18524
rect 23456 18468 23460 18524
rect 23396 18464 23460 18468
rect 23476 18524 23540 18528
rect 23476 18468 23480 18524
rect 23480 18468 23536 18524
rect 23536 18468 23540 18524
rect 23476 18464 23540 18468
rect 30664 18524 30728 18528
rect 30664 18468 30668 18524
rect 30668 18468 30724 18524
rect 30724 18468 30728 18524
rect 30664 18464 30728 18468
rect 30744 18524 30808 18528
rect 30744 18468 30748 18524
rect 30748 18468 30804 18524
rect 30804 18468 30808 18524
rect 30744 18464 30808 18468
rect 30824 18524 30888 18528
rect 30824 18468 30828 18524
rect 30828 18468 30884 18524
rect 30884 18468 30888 18524
rect 30824 18464 30888 18468
rect 30904 18524 30968 18528
rect 30904 18468 30908 18524
rect 30908 18468 30964 18524
rect 30964 18468 30968 18524
rect 30904 18464 30968 18468
rect 4666 17980 4730 17984
rect 4666 17924 4670 17980
rect 4670 17924 4726 17980
rect 4726 17924 4730 17980
rect 4666 17920 4730 17924
rect 4746 17980 4810 17984
rect 4746 17924 4750 17980
rect 4750 17924 4806 17980
rect 4806 17924 4810 17980
rect 4746 17920 4810 17924
rect 4826 17980 4890 17984
rect 4826 17924 4830 17980
rect 4830 17924 4886 17980
rect 4886 17924 4890 17980
rect 4826 17920 4890 17924
rect 4906 17980 4970 17984
rect 4906 17924 4910 17980
rect 4910 17924 4966 17980
rect 4966 17924 4970 17980
rect 4906 17920 4970 17924
rect 12094 17980 12158 17984
rect 12094 17924 12098 17980
rect 12098 17924 12154 17980
rect 12154 17924 12158 17980
rect 12094 17920 12158 17924
rect 12174 17980 12238 17984
rect 12174 17924 12178 17980
rect 12178 17924 12234 17980
rect 12234 17924 12238 17980
rect 12174 17920 12238 17924
rect 12254 17980 12318 17984
rect 12254 17924 12258 17980
rect 12258 17924 12314 17980
rect 12314 17924 12318 17980
rect 12254 17920 12318 17924
rect 12334 17980 12398 17984
rect 12334 17924 12338 17980
rect 12338 17924 12394 17980
rect 12394 17924 12398 17980
rect 12334 17920 12398 17924
rect 19522 17980 19586 17984
rect 19522 17924 19526 17980
rect 19526 17924 19582 17980
rect 19582 17924 19586 17980
rect 19522 17920 19586 17924
rect 19602 17980 19666 17984
rect 19602 17924 19606 17980
rect 19606 17924 19662 17980
rect 19662 17924 19666 17980
rect 19602 17920 19666 17924
rect 19682 17980 19746 17984
rect 19682 17924 19686 17980
rect 19686 17924 19742 17980
rect 19742 17924 19746 17980
rect 19682 17920 19746 17924
rect 19762 17980 19826 17984
rect 19762 17924 19766 17980
rect 19766 17924 19822 17980
rect 19822 17924 19826 17980
rect 19762 17920 19826 17924
rect 26950 17980 27014 17984
rect 26950 17924 26954 17980
rect 26954 17924 27010 17980
rect 27010 17924 27014 17980
rect 26950 17920 27014 17924
rect 27030 17980 27094 17984
rect 27030 17924 27034 17980
rect 27034 17924 27090 17980
rect 27090 17924 27094 17980
rect 27030 17920 27094 17924
rect 27110 17980 27174 17984
rect 27110 17924 27114 17980
rect 27114 17924 27170 17980
rect 27170 17924 27174 17980
rect 27110 17920 27174 17924
rect 27190 17980 27254 17984
rect 27190 17924 27194 17980
rect 27194 17924 27250 17980
rect 27250 17924 27254 17980
rect 27190 17920 27254 17924
rect 8380 17436 8444 17440
rect 8380 17380 8384 17436
rect 8384 17380 8440 17436
rect 8440 17380 8444 17436
rect 8380 17376 8444 17380
rect 8460 17436 8524 17440
rect 8460 17380 8464 17436
rect 8464 17380 8520 17436
rect 8520 17380 8524 17436
rect 8460 17376 8524 17380
rect 8540 17436 8604 17440
rect 8540 17380 8544 17436
rect 8544 17380 8600 17436
rect 8600 17380 8604 17436
rect 8540 17376 8604 17380
rect 8620 17436 8684 17440
rect 8620 17380 8624 17436
rect 8624 17380 8680 17436
rect 8680 17380 8684 17436
rect 8620 17376 8684 17380
rect 15808 17436 15872 17440
rect 15808 17380 15812 17436
rect 15812 17380 15868 17436
rect 15868 17380 15872 17436
rect 15808 17376 15872 17380
rect 15888 17436 15952 17440
rect 15888 17380 15892 17436
rect 15892 17380 15948 17436
rect 15948 17380 15952 17436
rect 15888 17376 15952 17380
rect 15968 17436 16032 17440
rect 15968 17380 15972 17436
rect 15972 17380 16028 17436
rect 16028 17380 16032 17436
rect 15968 17376 16032 17380
rect 16048 17436 16112 17440
rect 16048 17380 16052 17436
rect 16052 17380 16108 17436
rect 16108 17380 16112 17436
rect 16048 17376 16112 17380
rect 23236 17436 23300 17440
rect 23236 17380 23240 17436
rect 23240 17380 23296 17436
rect 23296 17380 23300 17436
rect 23236 17376 23300 17380
rect 23316 17436 23380 17440
rect 23316 17380 23320 17436
rect 23320 17380 23376 17436
rect 23376 17380 23380 17436
rect 23316 17376 23380 17380
rect 23396 17436 23460 17440
rect 23396 17380 23400 17436
rect 23400 17380 23456 17436
rect 23456 17380 23460 17436
rect 23396 17376 23460 17380
rect 23476 17436 23540 17440
rect 23476 17380 23480 17436
rect 23480 17380 23536 17436
rect 23536 17380 23540 17436
rect 23476 17376 23540 17380
rect 30664 17436 30728 17440
rect 30664 17380 30668 17436
rect 30668 17380 30724 17436
rect 30724 17380 30728 17436
rect 30664 17376 30728 17380
rect 30744 17436 30808 17440
rect 30744 17380 30748 17436
rect 30748 17380 30804 17436
rect 30804 17380 30808 17436
rect 30744 17376 30808 17380
rect 30824 17436 30888 17440
rect 30824 17380 30828 17436
rect 30828 17380 30884 17436
rect 30884 17380 30888 17436
rect 30824 17376 30888 17380
rect 30904 17436 30968 17440
rect 30904 17380 30908 17436
rect 30908 17380 30964 17436
rect 30964 17380 30968 17436
rect 30904 17376 30968 17380
rect 4666 16892 4730 16896
rect 4666 16836 4670 16892
rect 4670 16836 4726 16892
rect 4726 16836 4730 16892
rect 4666 16832 4730 16836
rect 4746 16892 4810 16896
rect 4746 16836 4750 16892
rect 4750 16836 4806 16892
rect 4806 16836 4810 16892
rect 4746 16832 4810 16836
rect 4826 16892 4890 16896
rect 4826 16836 4830 16892
rect 4830 16836 4886 16892
rect 4886 16836 4890 16892
rect 4826 16832 4890 16836
rect 4906 16892 4970 16896
rect 4906 16836 4910 16892
rect 4910 16836 4966 16892
rect 4966 16836 4970 16892
rect 4906 16832 4970 16836
rect 12094 16892 12158 16896
rect 12094 16836 12098 16892
rect 12098 16836 12154 16892
rect 12154 16836 12158 16892
rect 12094 16832 12158 16836
rect 12174 16892 12238 16896
rect 12174 16836 12178 16892
rect 12178 16836 12234 16892
rect 12234 16836 12238 16892
rect 12174 16832 12238 16836
rect 12254 16892 12318 16896
rect 12254 16836 12258 16892
rect 12258 16836 12314 16892
rect 12314 16836 12318 16892
rect 12254 16832 12318 16836
rect 12334 16892 12398 16896
rect 12334 16836 12338 16892
rect 12338 16836 12394 16892
rect 12394 16836 12398 16892
rect 12334 16832 12398 16836
rect 19522 16892 19586 16896
rect 19522 16836 19526 16892
rect 19526 16836 19582 16892
rect 19582 16836 19586 16892
rect 19522 16832 19586 16836
rect 19602 16892 19666 16896
rect 19602 16836 19606 16892
rect 19606 16836 19662 16892
rect 19662 16836 19666 16892
rect 19602 16832 19666 16836
rect 19682 16892 19746 16896
rect 19682 16836 19686 16892
rect 19686 16836 19742 16892
rect 19742 16836 19746 16892
rect 19682 16832 19746 16836
rect 19762 16892 19826 16896
rect 19762 16836 19766 16892
rect 19766 16836 19822 16892
rect 19822 16836 19826 16892
rect 19762 16832 19826 16836
rect 26950 16892 27014 16896
rect 26950 16836 26954 16892
rect 26954 16836 27010 16892
rect 27010 16836 27014 16892
rect 26950 16832 27014 16836
rect 27030 16892 27094 16896
rect 27030 16836 27034 16892
rect 27034 16836 27090 16892
rect 27090 16836 27094 16892
rect 27030 16832 27094 16836
rect 27110 16892 27174 16896
rect 27110 16836 27114 16892
rect 27114 16836 27170 16892
rect 27170 16836 27174 16892
rect 27110 16832 27174 16836
rect 27190 16892 27254 16896
rect 27190 16836 27194 16892
rect 27194 16836 27250 16892
rect 27250 16836 27254 16892
rect 27190 16832 27254 16836
rect 8380 16348 8444 16352
rect 8380 16292 8384 16348
rect 8384 16292 8440 16348
rect 8440 16292 8444 16348
rect 8380 16288 8444 16292
rect 8460 16348 8524 16352
rect 8460 16292 8464 16348
rect 8464 16292 8520 16348
rect 8520 16292 8524 16348
rect 8460 16288 8524 16292
rect 8540 16348 8604 16352
rect 8540 16292 8544 16348
rect 8544 16292 8600 16348
rect 8600 16292 8604 16348
rect 8540 16288 8604 16292
rect 8620 16348 8684 16352
rect 8620 16292 8624 16348
rect 8624 16292 8680 16348
rect 8680 16292 8684 16348
rect 8620 16288 8684 16292
rect 15808 16348 15872 16352
rect 15808 16292 15812 16348
rect 15812 16292 15868 16348
rect 15868 16292 15872 16348
rect 15808 16288 15872 16292
rect 15888 16348 15952 16352
rect 15888 16292 15892 16348
rect 15892 16292 15948 16348
rect 15948 16292 15952 16348
rect 15888 16288 15952 16292
rect 15968 16348 16032 16352
rect 15968 16292 15972 16348
rect 15972 16292 16028 16348
rect 16028 16292 16032 16348
rect 15968 16288 16032 16292
rect 16048 16348 16112 16352
rect 16048 16292 16052 16348
rect 16052 16292 16108 16348
rect 16108 16292 16112 16348
rect 16048 16288 16112 16292
rect 23236 16348 23300 16352
rect 23236 16292 23240 16348
rect 23240 16292 23296 16348
rect 23296 16292 23300 16348
rect 23236 16288 23300 16292
rect 23316 16348 23380 16352
rect 23316 16292 23320 16348
rect 23320 16292 23376 16348
rect 23376 16292 23380 16348
rect 23316 16288 23380 16292
rect 23396 16348 23460 16352
rect 23396 16292 23400 16348
rect 23400 16292 23456 16348
rect 23456 16292 23460 16348
rect 23396 16288 23460 16292
rect 23476 16348 23540 16352
rect 23476 16292 23480 16348
rect 23480 16292 23536 16348
rect 23536 16292 23540 16348
rect 23476 16288 23540 16292
rect 30664 16348 30728 16352
rect 30664 16292 30668 16348
rect 30668 16292 30724 16348
rect 30724 16292 30728 16348
rect 30664 16288 30728 16292
rect 30744 16348 30808 16352
rect 30744 16292 30748 16348
rect 30748 16292 30804 16348
rect 30804 16292 30808 16348
rect 30744 16288 30808 16292
rect 30824 16348 30888 16352
rect 30824 16292 30828 16348
rect 30828 16292 30884 16348
rect 30884 16292 30888 16348
rect 30824 16288 30888 16292
rect 30904 16348 30968 16352
rect 30904 16292 30908 16348
rect 30908 16292 30964 16348
rect 30964 16292 30968 16348
rect 30904 16288 30968 16292
rect 4666 15804 4730 15808
rect 4666 15748 4670 15804
rect 4670 15748 4726 15804
rect 4726 15748 4730 15804
rect 4666 15744 4730 15748
rect 4746 15804 4810 15808
rect 4746 15748 4750 15804
rect 4750 15748 4806 15804
rect 4806 15748 4810 15804
rect 4746 15744 4810 15748
rect 4826 15804 4890 15808
rect 4826 15748 4830 15804
rect 4830 15748 4886 15804
rect 4886 15748 4890 15804
rect 4826 15744 4890 15748
rect 4906 15804 4970 15808
rect 4906 15748 4910 15804
rect 4910 15748 4966 15804
rect 4966 15748 4970 15804
rect 4906 15744 4970 15748
rect 12094 15804 12158 15808
rect 12094 15748 12098 15804
rect 12098 15748 12154 15804
rect 12154 15748 12158 15804
rect 12094 15744 12158 15748
rect 12174 15804 12238 15808
rect 12174 15748 12178 15804
rect 12178 15748 12234 15804
rect 12234 15748 12238 15804
rect 12174 15744 12238 15748
rect 12254 15804 12318 15808
rect 12254 15748 12258 15804
rect 12258 15748 12314 15804
rect 12314 15748 12318 15804
rect 12254 15744 12318 15748
rect 12334 15804 12398 15808
rect 12334 15748 12338 15804
rect 12338 15748 12394 15804
rect 12394 15748 12398 15804
rect 12334 15744 12398 15748
rect 19522 15804 19586 15808
rect 19522 15748 19526 15804
rect 19526 15748 19582 15804
rect 19582 15748 19586 15804
rect 19522 15744 19586 15748
rect 19602 15804 19666 15808
rect 19602 15748 19606 15804
rect 19606 15748 19662 15804
rect 19662 15748 19666 15804
rect 19602 15744 19666 15748
rect 19682 15804 19746 15808
rect 19682 15748 19686 15804
rect 19686 15748 19742 15804
rect 19742 15748 19746 15804
rect 19682 15744 19746 15748
rect 19762 15804 19826 15808
rect 19762 15748 19766 15804
rect 19766 15748 19822 15804
rect 19822 15748 19826 15804
rect 19762 15744 19826 15748
rect 26950 15804 27014 15808
rect 26950 15748 26954 15804
rect 26954 15748 27010 15804
rect 27010 15748 27014 15804
rect 26950 15744 27014 15748
rect 27030 15804 27094 15808
rect 27030 15748 27034 15804
rect 27034 15748 27090 15804
rect 27090 15748 27094 15804
rect 27030 15744 27094 15748
rect 27110 15804 27174 15808
rect 27110 15748 27114 15804
rect 27114 15748 27170 15804
rect 27170 15748 27174 15804
rect 27110 15744 27174 15748
rect 27190 15804 27254 15808
rect 27190 15748 27194 15804
rect 27194 15748 27250 15804
rect 27250 15748 27254 15804
rect 27190 15744 27254 15748
rect 8380 15260 8444 15264
rect 8380 15204 8384 15260
rect 8384 15204 8440 15260
rect 8440 15204 8444 15260
rect 8380 15200 8444 15204
rect 8460 15260 8524 15264
rect 8460 15204 8464 15260
rect 8464 15204 8520 15260
rect 8520 15204 8524 15260
rect 8460 15200 8524 15204
rect 8540 15260 8604 15264
rect 8540 15204 8544 15260
rect 8544 15204 8600 15260
rect 8600 15204 8604 15260
rect 8540 15200 8604 15204
rect 8620 15260 8684 15264
rect 8620 15204 8624 15260
rect 8624 15204 8680 15260
rect 8680 15204 8684 15260
rect 8620 15200 8684 15204
rect 15808 15260 15872 15264
rect 15808 15204 15812 15260
rect 15812 15204 15868 15260
rect 15868 15204 15872 15260
rect 15808 15200 15872 15204
rect 15888 15260 15952 15264
rect 15888 15204 15892 15260
rect 15892 15204 15948 15260
rect 15948 15204 15952 15260
rect 15888 15200 15952 15204
rect 15968 15260 16032 15264
rect 15968 15204 15972 15260
rect 15972 15204 16028 15260
rect 16028 15204 16032 15260
rect 15968 15200 16032 15204
rect 16048 15260 16112 15264
rect 16048 15204 16052 15260
rect 16052 15204 16108 15260
rect 16108 15204 16112 15260
rect 16048 15200 16112 15204
rect 23236 15260 23300 15264
rect 23236 15204 23240 15260
rect 23240 15204 23296 15260
rect 23296 15204 23300 15260
rect 23236 15200 23300 15204
rect 23316 15260 23380 15264
rect 23316 15204 23320 15260
rect 23320 15204 23376 15260
rect 23376 15204 23380 15260
rect 23316 15200 23380 15204
rect 23396 15260 23460 15264
rect 23396 15204 23400 15260
rect 23400 15204 23456 15260
rect 23456 15204 23460 15260
rect 23396 15200 23460 15204
rect 23476 15260 23540 15264
rect 23476 15204 23480 15260
rect 23480 15204 23536 15260
rect 23536 15204 23540 15260
rect 23476 15200 23540 15204
rect 30664 15260 30728 15264
rect 30664 15204 30668 15260
rect 30668 15204 30724 15260
rect 30724 15204 30728 15260
rect 30664 15200 30728 15204
rect 30744 15260 30808 15264
rect 30744 15204 30748 15260
rect 30748 15204 30804 15260
rect 30804 15204 30808 15260
rect 30744 15200 30808 15204
rect 30824 15260 30888 15264
rect 30824 15204 30828 15260
rect 30828 15204 30884 15260
rect 30884 15204 30888 15260
rect 30824 15200 30888 15204
rect 30904 15260 30968 15264
rect 30904 15204 30908 15260
rect 30908 15204 30964 15260
rect 30964 15204 30968 15260
rect 30904 15200 30968 15204
rect 4666 14716 4730 14720
rect 4666 14660 4670 14716
rect 4670 14660 4726 14716
rect 4726 14660 4730 14716
rect 4666 14656 4730 14660
rect 4746 14716 4810 14720
rect 4746 14660 4750 14716
rect 4750 14660 4806 14716
rect 4806 14660 4810 14716
rect 4746 14656 4810 14660
rect 4826 14716 4890 14720
rect 4826 14660 4830 14716
rect 4830 14660 4886 14716
rect 4886 14660 4890 14716
rect 4826 14656 4890 14660
rect 4906 14716 4970 14720
rect 4906 14660 4910 14716
rect 4910 14660 4966 14716
rect 4966 14660 4970 14716
rect 4906 14656 4970 14660
rect 12094 14716 12158 14720
rect 12094 14660 12098 14716
rect 12098 14660 12154 14716
rect 12154 14660 12158 14716
rect 12094 14656 12158 14660
rect 12174 14716 12238 14720
rect 12174 14660 12178 14716
rect 12178 14660 12234 14716
rect 12234 14660 12238 14716
rect 12174 14656 12238 14660
rect 12254 14716 12318 14720
rect 12254 14660 12258 14716
rect 12258 14660 12314 14716
rect 12314 14660 12318 14716
rect 12254 14656 12318 14660
rect 12334 14716 12398 14720
rect 12334 14660 12338 14716
rect 12338 14660 12394 14716
rect 12394 14660 12398 14716
rect 12334 14656 12398 14660
rect 19522 14716 19586 14720
rect 19522 14660 19526 14716
rect 19526 14660 19582 14716
rect 19582 14660 19586 14716
rect 19522 14656 19586 14660
rect 19602 14716 19666 14720
rect 19602 14660 19606 14716
rect 19606 14660 19662 14716
rect 19662 14660 19666 14716
rect 19602 14656 19666 14660
rect 19682 14716 19746 14720
rect 19682 14660 19686 14716
rect 19686 14660 19742 14716
rect 19742 14660 19746 14716
rect 19682 14656 19746 14660
rect 19762 14716 19826 14720
rect 19762 14660 19766 14716
rect 19766 14660 19822 14716
rect 19822 14660 19826 14716
rect 19762 14656 19826 14660
rect 26950 14716 27014 14720
rect 26950 14660 26954 14716
rect 26954 14660 27010 14716
rect 27010 14660 27014 14716
rect 26950 14656 27014 14660
rect 27030 14716 27094 14720
rect 27030 14660 27034 14716
rect 27034 14660 27090 14716
rect 27090 14660 27094 14716
rect 27030 14656 27094 14660
rect 27110 14716 27174 14720
rect 27110 14660 27114 14716
rect 27114 14660 27170 14716
rect 27170 14660 27174 14716
rect 27110 14656 27174 14660
rect 27190 14716 27254 14720
rect 27190 14660 27194 14716
rect 27194 14660 27250 14716
rect 27250 14660 27254 14716
rect 27190 14656 27254 14660
rect 8380 14172 8444 14176
rect 8380 14116 8384 14172
rect 8384 14116 8440 14172
rect 8440 14116 8444 14172
rect 8380 14112 8444 14116
rect 8460 14172 8524 14176
rect 8460 14116 8464 14172
rect 8464 14116 8520 14172
rect 8520 14116 8524 14172
rect 8460 14112 8524 14116
rect 8540 14172 8604 14176
rect 8540 14116 8544 14172
rect 8544 14116 8600 14172
rect 8600 14116 8604 14172
rect 8540 14112 8604 14116
rect 8620 14172 8684 14176
rect 8620 14116 8624 14172
rect 8624 14116 8680 14172
rect 8680 14116 8684 14172
rect 8620 14112 8684 14116
rect 15808 14172 15872 14176
rect 15808 14116 15812 14172
rect 15812 14116 15868 14172
rect 15868 14116 15872 14172
rect 15808 14112 15872 14116
rect 15888 14172 15952 14176
rect 15888 14116 15892 14172
rect 15892 14116 15948 14172
rect 15948 14116 15952 14172
rect 15888 14112 15952 14116
rect 15968 14172 16032 14176
rect 15968 14116 15972 14172
rect 15972 14116 16028 14172
rect 16028 14116 16032 14172
rect 15968 14112 16032 14116
rect 16048 14172 16112 14176
rect 16048 14116 16052 14172
rect 16052 14116 16108 14172
rect 16108 14116 16112 14172
rect 16048 14112 16112 14116
rect 23236 14172 23300 14176
rect 23236 14116 23240 14172
rect 23240 14116 23296 14172
rect 23296 14116 23300 14172
rect 23236 14112 23300 14116
rect 23316 14172 23380 14176
rect 23316 14116 23320 14172
rect 23320 14116 23376 14172
rect 23376 14116 23380 14172
rect 23316 14112 23380 14116
rect 23396 14172 23460 14176
rect 23396 14116 23400 14172
rect 23400 14116 23456 14172
rect 23456 14116 23460 14172
rect 23396 14112 23460 14116
rect 23476 14172 23540 14176
rect 23476 14116 23480 14172
rect 23480 14116 23536 14172
rect 23536 14116 23540 14172
rect 23476 14112 23540 14116
rect 30664 14172 30728 14176
rect 30664 14116 30668 14172
rect 30668 14116 30724 14172
rect 30724 14116 30728 14172
rect 30664 14112 30728 14116
rect 30744 14172 30808 14176
rect 30744 14116 30748 14172
rect 30748 14116 30804 14172
rect 30804 14116 30808 14172
rect 30744 14112 30808 14116
rect 30824 14172 30888 14176
rect 30824 14116 30828 14172
rect 30828 14116 30884 14172
rect 30884 14116 30888 14172
rect 30824 14112 30888 14116
rect 30904 14172 30968 14176
rect 30904 14116 30908 14172
rect 30908 14116 30964 14172
rect 30964 14116 30968 14172
rect 30904 14112 30968 14116
rect 4666 13628 4730 13632
rect 4666 13572 4670 13628
rect 4670 13572 4726 13628
rect 4726 13572 4730 13628
rect 4666 13568 4730 13572
rect 4746 13628 4810 13632
rect 4746 13572 4750 13628
rect 4750 13572 4806 13628
rect 4806 13572 4810 13628
rect 4746 13568 4810 13572
rect 4826 13628 4890 13632
rect 4826 13572 4830 13628
rect 4830 13572 4886 13628
rect 4886 13572 4890 13628
rect 4826 13568 4890 13572
rect 4906 13628 4970 13632
rect 4906 13572 4910 13628
rect 4910 13572 4966 13628
rect 4966 13572 4970 13628
rect 4906 13568 4970 13572
rect 12094 13628 12158 13632
rect 12094 13572 12098 13628
rect 12098 13572 12154 13628
rect 12154 13572 12158 13628
rect 12094 13568 12158 13572
rect 12174 13628 12238 13632
rect 12174 13572 12178 13628
rect 12178 13572 12234 13628
rect 12234 13572 12238 13628
rect 12174 13568 12238 13572
rect 12254 13628 12318 13632
rect 12254 13572 12258 13628
rect 12258 13572 12314 13628
rect 12314 13572 12318 13628
rect 12254 13568 12318 13572
rect 12334 13628 12398 13632
rect 12334 13572 12338 13628
rect 12338 13572 12394 13628
rect 12394 13572 12398 13628
rect 12334 13568 12398 13572
rect 19522 13628 19586 13632
rect 19522 13572 19526 13628
rect 19526 13572 19582 13628
rect 19582 13572 19586 13628
rect 19522 13568 19586 13572
rect 19602 13628 19666 13632
rect 19602 13572 19606 13628
rect 19606 13572 19662 13628
rect 19662 13572 19666 13628
rect 19602 13568 19666 13572
rect 19682 13628 19746 13632
rect 19682 13572 19686 13628
rect 19686 13572 19742 13628
rect 19742 13572 19746 13628
rect 19682 13568 19746 13572
rect 19762 13628 19826 13632
rect 19762 13572 19766 13628
rect 19766 13572 19822 13628
rect 19822 13572 19826 13628
rect 19762 13568 19826 13572
rect 26950 13628 27014 13632
rect 26950 13572 26954 13628
rect 26954 13572 27010 13628
rect 27010 13572 27014 13628
rect 26950 13568 27014 13572
rect 27030 13628 27094 13632
rect 27030 13572 27034 13628
rect 27034 13572 27090 13628
rect 27090 13572 27094 13628
rect 27030 13568 27094 13572
rect 27110 13628 27174 13632
rect 27110 13572 27114 13628
rect 27114 13572 27170 13628
rect 27170 13572 27174 13628
rect 27110 13568 27174 13572
rect 27190 13628 27254 13632
rect 27190 13572 27194 13628
rect 27194 13572 27250 13628
rect 27250 13572 27254 13628
rect 27190 13568 27254 13572
rect 8380 13084 8444 13088
rect 8380 13028 8384 13084
rect 8384 13028 8440 13084
rect 8440 13028 8444 13084
rect 8380 13024 8444 13028
rect 8460 13084 8524 13088
rect 8460 13028 8464 13084
rect 8464 13028 8520 13084
rect 8520 13028 8524 13084
rect 8460 13024 8524 13028
rect 8540 13084 8604 13088
rect 8540 13028 8544 13084
rect 8544 13028 8600 13084
rect 8600 13028 8604 13084
rect 8540 13024 8604 13028
rect 8620 13084 8684 13088
rect 8620 13028 8624 13084
rect 8624 13028 8680 13084
rect 8680 13028 8684 13084
rect 8620 13024 8684 13028
rect 15808 13084 15872 13088
rect 15808 13028 15812 13084
rect 15812 13028 15868 13084
rect 15868 13028 15872 13084
rect 15808 13024 15872 13028
rect 15888 13084 15952 13088
rect 15888 13028 15892 13084
rect 15892 13028 15948 13084
rect 15948 13028 15952 13084
rect 15888 13024 15952 13028
rect 15968 13084 16032 13088
rect 15968 13028 15972 13084
rect 15972 13028 16028 13084
rect 16028 13028 16032 13084
rect 15968 13024 16032 13028
rect 16048 13084 16112 13088
rect 16048 13028 16052 13084
rect 16052 13028 16108 13084
rect 16108 13028 16112 13084
rect 16048 13024 16112 13028
rect 23236 13084 23300 13088
rect 23236 13028 23240 13084
rect 23240 13028 23296 13084
rect 23296 13028 23300 13084
rect 23236 13024 23300 13028
rect 23316 13084 23380 13088
rect 23316 13028 23320 13084
rect 23320 13028 23376 13084
rect 23376 13028 23380 13084
rect 23316 13024 23380 13028
rect 23396 13084 23460 13088
rect 23396 13028 23400 13084
rect 23400 13028 23456 13084
rect 23456 13028 23460 13084
rect 23396 13024 23460 13028
rect 23476 13084 23540 13088
rect 23476 13028 23480 13084
rect 23480 13028 23536 13084
rect 23536 13028 23540 13084
rect 23476 13024 23540 13028
rect 30664 13084 30728 13088
rect 30664 13028 30668 13084
rect 30668 13028 30724 13084
rect 30724 13028 30728 13084
rect 30664 13024 30728 13028
rect 30744 13084 30808 13088
rect 30744 13028 30748 13084
rect 30748 13028 30804 13084
rect 30804 13028 30808 13084
rect 30744 13024 30808 13028
rect 30824 13084 30888 13088
rect 30824 13028 30828 13084
rect 30828 13028 30884 13084
rect 30884 13028 30888 13084
rect 30824 13024 30888 13028
rect 30904 13084 30968 13088
rect 30904 13028 30908 13084
rect 30908 13028 30964 13084
rect 30964 13028 30968 13084
rect 30904 13024 30968 13028
rect 4666 12540 4730 12544
rect 4666 12484 4670 12540
rect 4670 12484 4726 12540
rect 4726 12484 4730 12540
rect 4666 12480 4730 12484
rect 4746 12540 4810 12544
rect 4746 12484 4750 12540
rect 4750 12484 4806 12540
rect 4806 12484 4810 12540
rect 4746 12480 4810 12484
rect 4826 12540 4890 12544
rect 4826 12484 4830 12540
rect 4830 12484 4886 12540
rect 4886 12484 4890 12540
rect 4826 12480 4890 12484
rect 4906 12540 4970 12544
rect 4906 12484 4910 12540
rect 4910 12484 4966 12540
rect 4966 12484 4970 12540
rect 4906 12480 4970 12484
rect 12094 12540 12158 12544
rect 12094 12484 12098 12540
rect 12098 12484 12154 12540
rect 12154 12484 12158 12540
rect 12094 12480 12158 12484
rect 12174 12540 12238 12544
rect 12174 12484 12178 12540
rect 12178 12484 12234 12540
rect 12234 12484 12238 12540
rect 12174 12480 12238 12484
rect 12254 12540 12318 12544
rect 12254 12484 12258 12540
rect 12258 12484 12314 12540
rect 12314 12484 12318 12540
rect 12254 12480 12318 12484
rect 12334 12540 12398 12544
rect 12334 12484 12338 12540
rect 12338 12484 12394 12540
rect 12394 12484 12398 12540
rect 12334 12480 12398 12484
rect 19522 12540 19586 12544
rect 19522 12484 19526 12540
rect 19526 12484 19582 12540
rect 19582 12484 19586 12540
rect 19522 12480 19586 12484
rect 19602 12540 19666 12544
rect 19602 12484 19606 12540
rect 19606 12484 19662 12540
rect 19662 12484 19666 12540
rect 19602 12480 19666 12484
rect 19682 12540 19746 12544
rect 19682 12484 19686 12540
rect 19686 12484 19742 12540
rect 19742 12484 19746 12540
rect 19682 12480 19746 12484
rect 19762 12540 19826 12544
rect 19762 12484 19766 12540
rect 19766 12484 19822 12540
rect 19822 12484 19826 12540
rect 19762 12480 19826 12484
rect 26950 12540 27014 12544
rect 26950 12484 26954 12540
rect 26954 12484 27010 12540
rect 27010 12484 27014 12540
rect 26950 12480 27014 12484
rect 27030 12540 27094 12544
rect 27030 12484 27034 12540
rect 27034 12484 27090 12540
rect 27090 12484 27094 12540
rect 27030 12480 27094 12484
rect 27110 12540 27174 12544
rect 27110 12484 27114 12540
rect 27114 12484 27170 12540
rect 27170 12484 27174 12540
rect 27110 12480 27174 12484
rect 27190 12540 27254 12544
rect 27190 12484 27194 12540
rect 27194 12484 27250 12540
rect 27250 12484 27254 12540
rect 27190 12480 27254 12484
rect 8380 11996 8444 12000
rect 8380 11940 8384 11996
rect 8384 11940 8440 11996
rect 8440 11940 8444 11996
rect 8380 11936 8444 11940
rect 8460 11996 8524 12000
rect 8460 11940 8464 11996
rect 8464 11940 8520 11996
rect 8520 11940 8524 11996
rect 8460 11936 8524 11940
rect 8540 11996 8604 12000
rect 8540 11940 8544 11996
rect 8544 11940 8600 11996
rect 8600 11940 8604 11996
rect 8540 11936 8604 11940
rect 8620 11996 8684 12000
rect 8620 11940 8624 11996
rect 8624 11940 8680 11996
rect 8680 11940 8684 11996
rect 8620 11936 8684 11940
rect 15808 11996 15872 12000
rect 15808 11940 15812 11996
rect 15812 11940 15868 11996
rect 15868 11940 15872 11996
rect 15808 11936 15872 11940
rect 15888 11996 15952 12000
rect 15888 11940 15892 11996
rect 15892 11940 15948 11996
rect 15948 11940 15952 11996
rect 15888 11936 15952 11940
rect 15968 11996 16032 12000
rect 15968 11940 15972 11996
rect 15972 11940 16028 11996
rect 16028 11940 16032 11996
rect 15968 11936 16032 11940
rect 16048 11996 16112 12000
rect 16048 11940 16052 11996
rect 16052 11940 16108 11996
rect 16108 11940 16112 11996
rect 16048 11936 16112 11940
rect 23236 11996 23300 12000
rect 23236 11940 23240 11996
rect 23240 11940 23296 11996
rect 23296 11940 23300 11996
rect 23236 11936 23300 11940
rect 23316 11996 23380 12000
rect 23316 11940 23320 11996
rect 23320 11940 23376 11996
rect 23376 11940 23380 11996
rect 23316 11936 23380 11940
rect 23396 11996 23460 12000
rect 23396 11940 23400 11996
rect 23400 11940 23456 11996
rect 23456 11940 23460 11996
rect 23396 11936 23460 11940
rect 23476 11996 23540 12000
rect 23476 11940 23480 11996
rect 23480 11940 23536 11996
rect 23536 11940 23540 11996
rect 23476 11936 23540 11940
rect 30664 11996 30728 12000
rect 30664 11940 30668 11996
rect 30668 11940 30724 11996
rect 30724 11940 30728 11996
rect 30664 11936 30728 11940
rect 30744 11996 30808 12000
rect 30744 11940 30748 11996
rect 30748 11940 30804 11996
rect 30804 11940 30808 11996
rect 30744 11936 30808 11940
rect 30824 11996 30888 12000
rect 30824 11940 30828 11996
rect 30828 11940 30884 11996
rect 30884 11940 30888 11996
rect 30824 11936 30888 11940
rect 30904 11996 30968 12000
rect 30904 11940 30908 11996
rect 30908 11940 30964 11996
rect 30964 11940 30968 11996
rect 30904 11936 30968 11940
rect 4666 11452 4730 11456
rect 4666 11396 4670 11452
rect 4670 11396 4726 11452
rect 4726 11396 4730 11452
rect 4666 11392 4730 11396
rect 4746 11452 4810 11456
rect 4746 11396 4750 11452
rect 4750 11396 4806 11452
rect 4806 11396 4810 11452
rect 4746 11392 4810 11396
rect 4826 11452 4890 11456
rect 4826 11396 4830 11452
rect 4830 11396 4886 11452
rect 4886 11396 4890 11452
rect 4826 11392 4890 11396
rect 4906 11452 4970 11456
rect 4906 11396 4910 11452
rect 4910 11396 4966 11452
rect 4966 11396 4970 11452
rect 4906 11392 4970 11396
rect 12094 11452 12158 11456
rect 12094 11396 12098 11452
rect 12098 11396 12154 11452
rect 12154 11396 12158 11452
rect 12094 11392 12158 11396
rect 12174 11452 12238 11456
rect 12174 11396 12178 11452
rect 12178 11396 12234 11452
rect 12234 11396 12238 11452
rect 12174 11392 12238 11396
rect 12254 11452 12318 11456
rect 12254 11396 12258 11452
rect 12258 11396 12314 11452
rect 12314 11396 12318 11452
rect 12254 11392 12318 11396
rect 12334 11452 12398 11456
rect 12334 11396 12338 11452
rect 12338 11396 12394 11452
rect 12394 11396 12398 11452
rect 12334 11392 12398 11396
rect 19522 11452 19586 11456
rect 19522 11396 19526 11452
rect 19526 11396 19582 11452
rect 19582 11396 19586 11452
rect 19522 11392 19586 11396
rect 19602 11452 19666 11456
rect 19602 11396 19606 11452
rect 19606 11396 19662 11452
rect 19662 11396 19666 11452
rect 19602 11392 19666 11396
rect 19682 11452 19746 11456
rect 19682 11396 19686 11452
rect 19686 11396 19742 11452
rect 19742 11396 19746 11452
rect 19682 11392 19746 11396
rect 19762 11452 19826 11456
rect 19762 11396 19766 11452
rect 19766 11396 19822 11452
rect 19822 11396 19826 11452
rect 19762 11392 19826 11396
rect 26950 11452 27014 11456
rect 26950 11396 26954 11452
rect 26954 11396 27010 11452
rect 27010 11396 27014 11452
rect 26950 11392 27014 11396
rect 27030 11452 27094 11456
rect 27030 11396 27034 11452
rect 27034 11396 27090 11452
rect 27090 11396 27094 11452
rect 27030 11392 27094 11396
rect 27110 11452 27174 11456
rect 27110 11396 27114 11452
rect 27114 11396 27170 11452
rect 27170 11396 27174 11452
rect 27110 11392 27174 11396
rect 27190 11452 27254 11456
rect 27190 11396 27194 11452
rect 27194 11396 27250 11452
rect 27250 11396 27254 11452
rect 27190 11392 27254 11396
rect 8380 10908 8444 10912
rect 8380 10852 8384 10908
rect 8384 10852 8440 10908
rect 8440 10852 8444 10908
rect 8380 10848 8444 10852
rect 8460 10908 8524 10912
rect 8460 10852 8464 10908
rect 8464 10852 8520 10908
rect 8520 10852 8524 10908
rect 8460 10848 8524 10852
rect 8540 10908 8604 10912
rect 8540 10852 8544 10908
rect 8544 10852 8600 10908
rect 8600 10852 8604 10908
rect 8540 10848 8604 10852
rect 8620 10908 8684 10912
rect 8620 10852 8624 10908
rect 8624 10852 8680 10908
rect 8680 10852 8684 10908
rect 8620 10848 8684 10852
rect 15808 10908 15872 10912
rect 15808 10852 15812 10908
rect 15812 10852 15868 10908
rect 15868 10852 15872 10908
rect 15808 10848 15872 10852
rect 15888 10908 15952 10912
rect 15888 10852 15892 10908
rect 15892 10852 15948 10908
rect 15948 10852 15952 10908
rect 15888 10848 15952 10852
rect 15968 10908 16032 10912
rect 15968 10852 15972 10908
rect 15972 10852 16028 10908
rect 16028 10852 16032 10908
rect 15968 10848 16032 10852
rect 16048 10908 16112 10912
rect 16048 10852 16052 10908
rect 16052 10852 16108 10908
rect 16108 10852 16112 10908
rect 16048 10848 16112 10852
rect 23236 10908 23300 10912
rect 23236 10852 23240 10908
rect 23240 10852 23296 10908
rect 23296 10852 23300 10908
rect 23236 10848 23300 10852
rect 23316 10908 23380 10912
rect 23316 10852 23320 10908
rect 23320 10852 23376 10908
rect 23376 10852 23380 10908
rect 23316 10848 23380 10852
rect 23396 10908 23460 10912
rect 23396 10852 23400 10908
rect 23400 10852 23456 10908
rect 23456 10852 23460 10908
rect 23396 10848 23460 10852
rect 23476 10908 23540 10912
rect 23476 10852 23480 10908
rect 23480 10852 23536 10908
rect 23536 10852 23540 10908
rect 23476 10848 23540 10852
rect 30664 10908 30728 10912
rect 30664 10852 30668 10908
rect 30668 10852 30724 10908
rect 30724 10852 30728 10908
rect 30664 10848 30728 10852
rect 30744 10908 30808 10912
rect 30744 10852 30748 10908
rect 30748 10852 30804 10908
rect 30804 10852 30808 10908
rect 30744 10848 30808 10852
rect 30824 10908 30888 10912
rect 30824 10852 30828 10908
rect 30828 10852 30884 10908
rect 30884 10852 30888 10908
rect 30824 10848 30888 10852
rect 30904 10908 30968 10912
rect 30904 10852 30908 10908
rect 30908 10852 30964 10908
rect 30964 10852 30968 10908
rect 30904 10848 30968 10852
rect 4666 10364 4730 10368
rect 4666 10308 4670 10364
rect 4670 10308 4726 10364
rect 4726 10308 4730 10364
rect 4666 10304 4730 10308
rect 4746 10364 4810 10368
rect 4746 10308 4750 10364
rect 4750 10308 4806 10364
rect 4806 10308 4810 10364
rect 4746 10304 4810 10308
rect 4826 10364 4890 10368
rect 4826 10308 4830 10364
rect 4830 10308 4886 10364
rect 4886 10308 4890 10364
rect 4826 10304 4890 10308
rect 4906 10364 4970 10368
rect 4906 10308 4910 10364
rect 4910 10308 4966 10364
rect 4966 10308 4970 10364
rect 4906 10304 4970 10308
rect 12094 10364 12158 10368
rect 12094 10308 12098 10364
rect 12098 10308 12154 10364
rect 12154 10308 12158 10364
rect 12094 10304 12158 10308
rect 12174 10364 12238 10368
rect 12174 10308 12178 10364
rect 12178 10308 12234 10364
rect 12234 10308 12238 10364
rect 12174 10304 12238 10308
rect 12254 10364 12318 10368
rect 12254 10308 12258 10364
rect 12258 10308 12314 10364
rect 12314 10308 12318 10364
rect 12254 10304 12318 10308
rect 12334 10364 12398 10368
rect 12334 10308 12338 10364
rect 12338 10308 12394 10364
rect 12394 10308 12398 10364
rect 12334 10304 12398 10308
rect 19522 10364 19586 10368
rect 19522 10308 19526 10364
rect 19526 10308 19582 10364
rect 19582 10308 19586 10364
rect 19522 10304 19586 10308
rect 19602 10364 19666 10368
rect 19602 10308 19606 10364
rect 19606 10308 19662 10364
rect 19662 10308 19666 10364
rect 19602 10304 19666 10308
rect 19682 10364 19746 10368
rect 19682 10308 19686 10364
rect 19686 10308 19742 10364
rect 19742 10308 19746 10364
rect 19682 10304 19746 10308
rect 19762 10364 19826 10368
rect 19762 10308 19766 10364
rect 19766 10308 19822 10364
rect 19822 10308 19826 10364
rect 19762 10304 19826 10308
rect 26950 10364 27014 10368
rect 26950 10308 26954 10364
rect 26954 10308 27010 10364
rect 27010 10308 27014 10364
rect 26950 10304 27014 10308
rect 27030 10364 27094 10368
rect 27030 10308 27034 10364
rect 27034 10308 27090 10364
rect 27090 10308 27094 10364
rect 27030 10304 27094 10308
rect 27110 10364 27174 10368
rect 27110 10308 27114 10364
rect 27114 10308 27170 10364
rect 27170 10308 27174 10364
rect 27110 10304 27174 10308
rect 27190 10364 27254 10368
rect 27190 10308 27194 10364
rect 27194 10308 27250 10364
rect 27250 10308 27254 10364
rect 27190 10304 27254 10308
rect 8380 9820 8444 9824
rect 8380 9764 8384 9820
rect 8384 9764 8440 9820
rect 8440 9764 8444 9820
rect 8380 9760 8444 9764
rect 8460 9820 8524 9824
rect 8460 9764 8464 9820
rect 8464 9764 8520 9820
rect 8520 9764 8524 9820
rect 8460 9760 8524 9764
rect 8540 9820 8604 9824
rect 8540 9764 8544 9820
rect 8544 9764 8600 9820
rect 8600 9764 8604 9820
rect 8540 9760 8604 9764
rect 8620 9820 8684 9824
rect 8620 9764 8624 9820
rect 8624 9764 8680 9820
rect 8680 9764 8684 9820
rect 8620 9760 8684 9764
rect 15808 9820 15872 9824
rect 15808 9764 15812 9820
rect 15812 9764 15868 9820
rect 15868 9764 15872 9820
rect 15808 9760 15872 9764
rect 15888 9820 15952 9824
rect 15888 9764 15892 9820
rect 15892 9764 15948 9820
rect 15948 9764 15952 9820
rect 15888 9760 15952 9764
rect 15968 9820 16032 9824
rect 15968 9764 15972 9820
rect 15972 9764 16028 9820
rect 16028 9764 16032 9820
rect 15968 9760 16032 9764
rect 16048 9820 16112 9824
rect 16048 9764 16052 9820
rect 16052 9764 16108 9820
rect 16108 9764 16112 9820
rect 16048 9760 16112 9764
rect 23236 9820 23300 9824
rect 23236 9764 23240 9820
rect 23240 9764 23296 9820
rect 23296 9764 23300 9820
rect 23236 9760 23300 9764
rect 23316 9820 23380 9824
rect 23316 9764 23320 9820
rect 23320 9764 23376 9820
rect 23376 9764 23380 9820
rect 23316 9760 23380 9764
rect 23396 9820 23460 9824
rect 23396 9764 23400 9820
rect 23400 9764 23456 9820
rect 23456 9764 23460 9820
rect 23396 9760 23460 9764
rect 23476 9820 23540 9824
rect 23476 9764 23480 9820
rect 23480 9764 23536 9820
rect 23536 9764 23540 9820
rect 23476 9760 23540 9764
rect 30664 9820 30728 9824
rect 30664 9764 30668 9820
rect 30668 9764 30724 9820
rect 30724 9764 30728 9820
rect 30664 9760 30728 9764
rect 30744 9820 30808 9824
rect 30744 9764 30748 9820
rect 30748 9764 30804 9820
rect 30804 9764 30808 9820
rect 30744 9760 30808 9764
rect 30824 9820 30888 9824
rect 30824 9764 30828 9820
rect 30828 9764 30884 9820
rect 30884 9764 30888 9820
rect 30824 9760 30888 9764
rect 30904 9820 30968 9824
rect 30904 9764 30908 9820
rect 30908 9764 30964 9820
rect 30964 9764 30968 9820
rect 30904 9760 30968 9764
rect 4666 9276 4730 9280
rect 4666 9220 4670 9276
rect 4670 9220 4726 9276
rect 4726 9220 4730 9276
rect 4666 9216 4730 9220
rect 4746 9276 4810 9280
rect 4746 9220 4750 9276
rect 4750 9220 4806 9276
rect 4806 9220 4810 9276
rect 4746 9216 4810 9220
rect 4826 9276 4890 9280
rect 4826 9220 4830 9276
rect 4830 9220 4886 9276
rect 4886 9220 4890 9276
rect 4826 9216 4890 9220
rect 4906 9276 4970 9280
rect 4906 9220 4910 9276
rect 4910 9220 4966 9276
rect 4966 9220 4970 9276
rect 4906 9216 4970 9220
rect 12094 9276 12158 9280
rect 12094 9220 12098 9276
rect 12098 9220 12154 9276
rect 12154 9220 12158 9276
rect 12094 9216 12158 9220
rect 12174 9276 12238 9280
rect 12174 9220 12178 9276
rect 12178 9220 12234 9276
rect 12234 9220 12238 9276
rect 12174 9216 12238 9220
rect 12254 9276 12318 9280
rect 12254 9220 12258 9276
rect 12258 9220 12314 9276
rect 12314 9220 12318 9276
rect 12254 9216 12318 9220
rect 12334 9276 12398 9280
rect 12334 9220 12338 9276
rect 12338 9220 12394 9276
rect 12394 9220 12398 9276
rect 12334 9216 12398 9220
rect 19522 9276 19586 9280
rect 19522 9220 19526 9276
rect 19526 9220 19582 9276
rect 19582 9220 19586 9276
rect 19522 9216 19586 9220
rect 19602 9276 19666 9280
rect 19602 9220 19606 9276
rect 19606 9220 19662 9276
rect 19662 9220 19666 9276
rect 19602 9216 19666 9220
rect 19682 9276 19746 9280
rect 19682 9220 19686 9276
rect 19686 9220 19742 9276
rect 19742 9220 19746 9276
rect 19682 9216 19746 9220
rect 19762 9276 19826 9280
rect 19762 9220 19766 9276
rect 19766 9220 19822 9276
rect 19822 9220 19826 9276
rect 19762 9216 19826 9220
rect 26950 9276 27014 9280
rect 26950 9220 26954 9276
rect 26954 9220 27010 9276
rect 27010 9220 27014 9276
rect 26950 9216 27014 9220
rect 27030 9276 27094 9280
rect 27030 9220 27034 9276
rect 27034 9220 27090 9276
rect 27090 9220 27094 9276
rect 27030 9216 27094 9220
rect 27110 9276 27174 9280
rect 27110 9220 27114 9276
rect 27114 9220 27170 9276
rect 27170 9220 27174 9276
rect 27110 9216 27174 9220
rect 27190 9276 27254 9280
rect 27190 9220 27194 9276
rect 27194 9220 27250 9276
rect 27250 9220 27254 9276
rect 27190 9216 27254 9220
rect 8380 8732 8444 8736
rect 8380 8676 8384 8732
rect 8384 8676 8440 8732
rect 8440 8676 8444 8732
rect 8380 8672 8444 8676
rect 8460 8732 8524 8736
rect 8460 8676 8464 8732
rect 8464 8676 8520 8732
rect 8520 8676 8524 8732
rect 8460 8672 8524 8676
rect 8540 8732 8604 8736
rect 8540 8676 8544 8732
rect 8544 8676 8600 8732
rect 8600 8676 8604 8732
rect 8540 8672 8604 8676
rect 8620 8732 8684 8736
rect 8620 8676 8624 8732
rect 8624 8676 8680 8732
rect 8680 8676 8684 8732
rect 8620 8672 8684 8676
rect 15808 8732 15872 8736
rect 15808 8676 15812 8732
rect 15812 8676 15868 8732
rect 15868 8676 15872 8732
rect 15808 8672 15872 8676
rect 15888 8732 15952 8736
rect 15888 8676 15892 8732
rect 15892 8676 15948 8732
rect 15948 8676 15952 8732
rect 15888 8672 15952 8676
rect 15968 8732 16032 8736
rect 15968 8676 15972 8732
rect 15972 8676 16028 8732
rect 16028 8676 16032 8732
rect 15968 8672 16032 8676
rect 16048 8732 16112 8736
rect 16048 8676 16052 8732
rect 16052 8676 16108 8732
rect 16108 8676 16112 8732
rect 16048 8672 16112 8676
rect 23236 8732 23300 8736
rect 23236 8676 23240 8732
rect 23240 8676 23296 8732
rect 23296 8676 23300 8732
rect 23236 8672 23300 8676
rect 23316 8732 23380 8736
rect 23316 8676 23320 8732
rect 23320 8676 23376 8732
rect 23376 8676 23380 8732
rect 23316 8672 23380 8676
rect 23396 8732 23460 8736
rect 23396 8676 23400 8732
rect 23400 8676 23456 8732
rect 23456 8676 23460 8732
rect 23396 8672 23460 8676
rect 23476 8732 23540 8736
rect 23476 8676 23480 8732
rect 23480 8676 23536 8732
rect 23536 8676 23540 8732
rect 23476 8672 23540 8676
rect 30664 8732 30728 8736
rect 30664 8676 30668 8732
rect 30668 8676 30724 8732
rect 30724 8676 30728 8732
rect 30664 8672 30728 8676
rect 30744 8732 30808 8736
rect 30744 8676 30748 8732
rect 30748 8676 30804 8732
rect 30804 8676 30808 8732
rect 30744 8672 30808 8676
rect 30824 8732 30888 8736
rect 30824 8676 30828 8732
rect 30828 8676 30884 8732
rect 30884 8676 30888 8732
rect 30824 8672 30888 8676
rect 30904 8732 30968 8736
rect 30904 8676 30908 8732
rect 30908 8676 30964 8732
rect 30964 8676 30968 8732
rect 30904 8672 30968 8676
rect 4666 8188 4730 8192
rect 4666 8132 4670 8188
rect 4670 8132 4726 8188
rect 4726 8132 4730 8188
rect 4666 8128 4730 8132
rect 4746 8188 4810 8192
rect 4746 8132 4750 8188
rect 4750 8132 4806 8188
rect 4806 8132 4810 8188
rect 4746 8128 4810 8132
rect 4826 8188 4890 8192
rect 4826 8132 4830 8188
rect 4830 8132 4886 8188
rect 4886 8132 4890 8188
rect 4826 8128 4890 8132
rect 4906 8188 4970 8192
rect 4906 8132 4910 8188
rect 4910 8132 4966 8188
rect 4966 8132 4970 8188
rect 4906 8128 4970 8132
rect 12094 8188 12158 8192
rect 12094 8132 12098 8188
rect 12098 8132 12154 8188
rect 12154 8132 12158 8188
rect 12094 8128 12158 8132
rect 12174 8188 12238 8192
rect 12174 8132 12178 8188
rect 12178 8132 12234 8188
rect 12234 8132 12238 8188
rect 12174 8128 12238 8132
rect 12254 8188 12318 8192
rect 12254 8132 12258 8188
rect 12258 8132 12314 8188
rect 12314 8132 12318 8188
rect 12254 8128 12318 8132
rect 12334 8188 12398 8192
rect 12334 8132 12338 8188
rect 12338 8132 12394 8188
rect 12394 8132 12398 8188
rect 12334 8128 12398 8132
rect 19522 8188 19586 8192
rect 19522 8132 19526 8188
rect 19526 8132 19582 8188
rect 19582 8132 19586 8188
rect 19522 8128 19586 8132
rect 19602 8188 19666 8192
rect 19602 8132 19606 8188
rect 19606 8132 19662 8188
rect 19662 8132 19666 8188
rect 19602 8128 19666 8132
rect 19682 8188 19746 8192
rect 19682 8132 19686 8188
rect 19686 8132 19742 8188
rect 19742 8132 19746 8188
rect 19682 8128 19746 8132
rect 19762 8188 19826 8192
rect 19762 8132 19766 8188
rect 19766 8132 19822 8188
rect 19822 8132 19826 8188
rect 19762 8128 19826 8132
rect 26950 8188 27014 8192
rect 26950 8132 26954 8188
rect 26954 8132 27010 8188
rect 27010 8132 27014 8188
rect 26950 8128 27014 8132
rect 27030 8188 27094 8192
rect 27030 8132 27034 8188
rect 27034 8132 27090 8188
rect 27090 8132 27094 8188
rect 27030 8128 27094 8132
rect 27110 8188 27174 8192
rect 27110 8132 27114 8188
rect 27114 8132 27170 8188
rect 27170 8132 27174 8188
rect 27110 8128 27174 8132
rect 27190 8188 27254 8192
rect 27190 8132 27194 8188
rect 27194 8132 27250 8188
rect 27250 8132 27254 8188
rect 27190 8128 27254 8132
rect 8380 7644 8444 7648
rect 8380 7588 8384 7644
rect 8384 7588 8440 7644
rect 8440 7588 8444 7644
rect 8380 7584 8444 7588
rect 8460 7644 8524 7648
rect 8460 7588 8464 7644
rect 8464 7588 8520 7644
rect 8520 7588 8524 7644
rect 8460 7584 8524 7588
rect 8540 7644 8604 7648
rect 8540 7588 8544 7644
rect 8544 7588 8600 7644
rect 8600 7588 8604 7644
rect 8540 7584 8604 7588
rect 8620 7644 8684 7648
rect 8620 7588 8624 7644
rect 8624 7588 8680 7644
rect 8680 7588 8684 7644
rect 8620 7584 8684 7588
rect 15808 7644 15872 7648
rect 15808 7588 15812 7644
rect 15812 7588 15868 7644
rect 15868 7588 15872 7644
rect 15808 7584 15872 7588
rect 15888 7644 15952 7648
rect 15888 7588 15892 7644
rect 15892 7588 15948 7644
rect 15948 7588 15952 7644
rect 15888 7584 15952 7588
rect 15968 7644 16032 7648
rect 15968 7588 15972 7644
rect 15972 7588 16028 7644
rect 16028 7588 16032 7644
rect 15968 7584 16032 7588
rect 16048 7644 16112 7648
rect 16048 7588 16052 7644
rect 16052 7588 16108 7644
rect 16108 7588 16112 7644
rect 16048 7584 16112 7588
rect 23236 7644 23300 7648
rect 23236 7588 23240 7644
rect 23240 7588 23296 7644
rect 23296 7588 23300 7644
rect 23236 7584 23300 7588
rect 23316 7644 23380 7648
rect 23316 7588 23320 7644
rect 23320 7588 23376 7644
rect 23376 7588 23380 7644
rect 23316 7584 23380 7588
rect 23396 7644 23460 7648
rect 23396 7588 23400 7644
rect 23400 7588 23456 7644
rect 23456 7588 23460 7644
rect 23396 7584 23460 7588
rect 23476 7644 23540 7648
rect 23476 7588 23480 7644
rect 23480 7588 23536 7644
rect 23536 7588 23540 7644
rect 23476 7584 23540 7588
rect 30664 7644 30728 7648
rect 30664 7588 30668 7644
rect 30668 7588 30724 7644
rect 30724 7588 30728 7644
rect 30664 7584 30728 7588
rect 30744 7644 30808 7648
rect 30744 7588 30748 7644
rect 30748 7588 30804 7644
rect 30804 7588 30808 7644
rect 30744 7584 30808 7588
rect 30824 7644 30888 7648
rect 30824 7588 30828 7644
rect 30828 7588 30884 7644
rect 30884 7588 30888 7644
rect 30824 7584 30888 7588
rect 30904 7644 30968 7648
rect 30904 7588 30908 7644
rect 30908 7588 30964 7644
rect 30964 7588 30968 7644
rect 30904 7584 30968 7588
rect 4666 7100 4730 7104
rect 4666 7044 4670 7100
rect 4670 7044 4726 7100
rect 4726 7044 4730 7100
rect 4666 7040 4730 7044
rect 4746 7100 4810 7104
rect 4746 7044 4750 7100
rect 4750 7044 4806 7100
rect 4806 7044 4810 7100
rect 4746 7040 4810 7044
rect 4826 7100 4890 7104
rect 4826 7044 4830 7100
rect 4830 7044 4886 7100
rect 4886 7044 4890 7100
rect 4826 7040 4890 7044
rect 4906 7100 4970 7104
rect 4906 7044 4910 7100
rect 4910 7044 4966 7100
rect 4966 7044 4970 7100
rect 4906 7040 4970 7044
rect 12094 7100 12158 7104
rect 12094 7044 12098 7100
rect 12098 7044 12154 7100
rect 12154 7044 12158 7100
rect 12094 7040 12158 7044
rect 12174 7100 12238 7104
rect 12174 7044 12178 7100
rect 12178 7044 12234 7100
rect 12234 7044 12238 7100
rect 12174 7040 12238 7044
rect 12254 7100 12318 7104
rect 12254 7044 12258 7100
rect 12258 7044 12314 7100
rect 12314 7044 12318 7100
rect 12254 7040 12318 7044
rect 12334 7100 12398 7104
rect 12334 7044 12338 7100
rect 12338 7044 12394 7100
rect 12394 7044 12398 7100
rect 12334 7040 12398 7044
rect 19522 7100 19586 7104
rect 19522 7044 19526 7100
rect 19526 7044 19582 7100
rect 19582 7044 19586 7100
rect 19522 7040 19586 7044
rect 19602 7100 19666 7104
rect 19602 7044 19606 7100
rect 19606 7044 19662 7100
rect 19662 7044 19666 7100
rect 19602 7040 19666 7044
rect 19682 7100 19746 7104
rect 19682 7044 19686 7100
rect 19686 7044 19742 7100
rect 19742 7044 19746 7100
rect 19682 7040 19746 7044
rect 19762 7100 19826 7104
rect 19762 7044 19766 7100
rect 19766 7044 19822 7100
rect 19822 7044 19826 7100
rect 19762 7040 19826 7044
rect 26950 7100 27014 7104
rect 26950 7044 26954 7100
rect 26954 7044 27010 7100
rect 27010 7044 27014 7100
rect 26950 7040 27014 7044
rect 27030 7100 27094 7104
rect 27030 7044 27034 7100
rect 27034 7044 27090 7100
rect 27090 7044 27094 7100
rect 27030 7040 27094 7044
rect 27110 7100 27174 7104
rect 27110 7044 27114 7100
rect 27114 7044 27170 7100
rect 27170 7044 27174 7100
rect 27110 7040 27174 7044
rect 27190 7100 27254 7104
rect 27190 7044 27194 7100
rect 27194 7044 27250 7100
rect 27250 7044 27254 7100
rect 27190 7040 27254 7044
rect 8380 6556 8444 6560
rect 8380 6500 8384 6556
rect 8384 6500 8440 6556
rect 8440 6500 8444 6556
rect 8380 6496 8444 6500
rect 8460 6556 8524 6560
rect 8460 6500 8464 6556
rect 8464 6500 8520 6556
rect 8520 6500 8524 6556
rect 8460 6496 8524 6500
rect 8540 6556 8604 6560
rect 8540 6500 8544 6556
rect 8544 6500 8600 6556
rect 8600 6500 8604 6556
rect 8540 6496 8604 6500
rect 8620 6556 8684 6560
rect 8620 6500 8624 6556
rect 8624 6500 8680 6556
rect 8680 6500 8684 6556
rect 8620 6496 8684 6500
rect 15808 6556 15872 6560
rect 15808 6500 15812 6556
rect 15812 6500 15868 6556
rect 15868 6500 15872 6556
rect 15808 6496 15872 6500
rect 15888 6556 15952 6560
rect 15888 6500 15892 6556
rect 15892 6500 15948 6556
rect 15948 6500 15952 6556
rect 15888 6496 15952 6500
rect 15968 6556 16032 6560
rect 15968 6500 15972 6556
rect 15972 6500 16028 6556
rect 16028 6500 16032 6556
rect 15968 6496 16032 6500
rect 16048 6556 16112 6560
rect 16048 6500 16052 6556
rect 16052 6500 16108 6556
rect 16108 6500 16112 6556
rect 16048 6496 16112 6500
rect 23236 6556 23300 6560
rect 23236 6500 23240 6556
rect 23240 6500 23296 6556
rect 23296 6500 23300 6556
rect 23236 6496 23300 6500
rect 23316 6556 23380 6560
rect 23316 6500 23320 6556
rect 23320 6500 23376 6556
rect 23376 6500 23380 6556
rect 23316 6496 23380 6500
rect 23396 6556 23460 6560
rect 23396 6500 23400 6556
rect 23400 6500 23456 6556
rect 23456 6500 23460 6556
rect 23396 6496 23460 6500
rect 23476 6556 23540 6560
rect 23476 6500 23480 6556
rect 23480 6500 23536 6556
rect 23536 6500 23540 6556
rect 23476 6496 23540 6500
rect 30664 6556 30728 6560
rect 30664 6500 30668 6556
rect 30668 6500 30724 6556
rect 30724 6500 30728 6556
rect 30664 6496 30728 6500
rect 30744 6556 30808 6560
rect 30744 6500 30748 6556
rect 30748 6500 30804 6556
rect 30804 6500 30808 6556
rect 30744 6496 30808 6500
rect 30824 6556 30888 6560
rect 30824 6500 30828 6556
rect 30828 6500 30884 6556
rect 30884 6500 30888 6556
rect 30824 6496 30888 6500
rect 30904 6556 30968 6560
rect 30904 6500 30908 6556
rect 30908 6500 30964 6556
rect 30964 6500 30968 6556
rect 30904 6496 30968 6500
rect 4666 6012 4730 6016
rect 4666 5956 4670 6012
rect 4670 5956 4726 6012
rect 4726 5956 4730 6012
rect 4666 5952 4730 5956
rect 4746 6012 4810 6016
rect 4746 5956 4750 6012
rect 4750 5956 4806 6012
rect 4806 5956 4810 6012
rect 4746 5952 4810 5956
rect 4826 6012 4890 6016
rect 4826 5956 4830 6012
rect 4830 5956 4886 6012
rect 4886 5956 4890 6012
rect 4826 5952 4890 5956
rect 4906 6012 4970 6016
rect 4906 5956 4910 6012
rect 4910 5956 4966 6012
rect 4966 5956 4970 6012
rect 4906 5952 4970 5956
rect 12094 6012 12158 6016
rect 12094 5956 12098 6012
rect 12098 5956 12154 6012
rect 12154 5956 12158 6012
rect 12094 5952 12158 5956
rect 12174 6012 12238 6016
rect 12174 5956 12178 6012
rect 12178 5956 12234 6012
rect 12234 5956 12238 6012
rect 12174 5952 12238 5956
rect 12254 6012 12318 6016
rect 12254 5956 12258 6012
rect 12258 5956 12314 6012
rect 12314 5956 12318 6012
rect 12254 5952 12318 5956
rect 12334 6012 12398 6016
rect 12334 5956 12338 6012
rect 12338 5956 12394 6012
rect 12394 5956 12398 6012
rect 12334 5952 12398 5956
rect 19522 6012 19586 6016
rect 19522 5956 19526 6012
rect 19526 5956 19582 6012
rect 19582 5956 19586 6012
rect 19522 5952 19586 5956
rect 19602 6012 19666 6016
rect 19602 5956 19606 6012
rect 19606 5956 19662 6012
rect 19662 5956 19666 6012
rect 19602 5952 19666 5956
rect 19682 6012 19746 6016
rect 19682 5956 19686 6012
rect 19686 5956 19742 6012
rect 19742 5956 19746 6012
rect 19682 5952 19746 5956
rect 19762 6012 19826 6016
rect 19762 5956 19766 6012
rect 19766 5956 19822 6012
rect 19822 5956 19826 6012
rect 19762 5952 19826 5956
rect 26950 6012 27014 6016
rect 26950 5956 26954 6012
rect 26954 5956 27010 6012
rect 27010 5956 27014 6012
rect 26950 5952 27014 5956
rect 27030 6012 27094 6016
rect 27030 5956 27034 6012
rect 27034 5956 27090 6012
rect 27090 5956 27094 6012
rect 27030 5952 27094 5956
rect 27110 6012 27174 6016
rect 27110 5956 27114 6012
rect 27114 5956 27170 6012
rect 27170 5956 27174 6012
rect 27110 5952 27174 5956
rect 27190 6012 27254 6016
rect 27190 5956 27194 6012
rect 27194 5956 27250 6012
rect 27250 5956 27254 6012
rect 27190 5952 27254 5956
rect 8380 5468 8444 5472
rect 8380 5412 8384 5468
rect 8384 5412 8440 5468
rect 8440 5412 8444 5468
rect 8380 5408 8444 5412
rect 8460 5468 8524 5472
rect 8460 5412 8464 5468
rect 8464 5412 8520 5468
rect 8520 5412 8524 5468
rect 8460 5408 8524 5412
rect 8540 5468 8604 5472
rect 8540 5412 8544 5468
rect 8544 5412 8600 5468
rect 8600 5412 8604 5468
rect 8540 5408 8604 5412
rect 8620 5468 8684 5472
rect 8620 5412 8624 5468
rect 8624 5412 8680 5468
rect 8680 5412 8684 5468
rect 8620 5408 8684 5412
rect 15808 5468 15872 5472
rect 15808 5412 15812 5468
rect 15812 5412 15868 5468
rect 15868 5412 15872 5468
rect 15808 5408 15872 5412
rect 15888 5468 15952 5472
rect 15888 5412 15892 5468
rect 15892 5412 15948 5468
rect 15948 5412 15952 5468
rect 15888 5408 15952 5412
rect 15968 5468 16032 5472
rect 15968 5412 15972 5468
rect 15972 5412 16028 5468
rect 16028 5412 16032 5468
rect 15968 5408 16032 5412
rect 16048 5468 16112 5472
rect 16048 5412 16052 5468
rect 16052 5412 16108 5468
rect 16108 5412 16112 5468
rect 16048 5408 16112 5412
rect 23236 5468 23300 5472
rect 23236 5412 23240 5468
rect 23240 5412 23296 5468
rect 23296 5412 23300 5468
rect 23236 5408 23300 5412
rect 23316 5468 23380 5472
rect 23316 5412 23320 5468
rect 23320 5412 23376 5468
rect 23376 5412 23380 5468
rect 23316 5408 23380 5412
rect 23396 5468 23460 5472
rect 23396 5412 23400 5468
rect 23400 5412 23456 5468
rect 23456 5412 23460 5468
rect 23396 5408 23460 5412
rect 23476 5468 23540 5472
rect 23476 5412 23480 5468
rect 23480 5412 23536 5468
rect 23536 5412 23540 5468
rect 23476 5408 23540 5412
rect 30664 5468 30728 5472
rect 30664 5412 30668 5468
rect 30668 5412 30724 5468
rect 30724 5412 30728 5468
rect 30664 5408 30728 5412
rect 30744 5468 30808 5472
rect 30744 5412 30748 5468
rect 30748 5412 30804 5468
rect 30804 5412 30808 5468
rect 30744 5408 30808 5412
rect 30824 5468 30888 5472
rect 30824 5412 30828 5468
rect 30828 5412 30884 5468
rect 30884 5412 30888 5468
rect 30824 5408 30888 5412
rect 30904 5468 30968 5472
rect 30904 5412 30908 5468
rect 30908 5412 30964 5468
rect 30964 5412 30968 5468
rect 30904 5408 30968 5412
rect 4666 4924 4730 4928
rect 4666 4868 4670 4924
rect 4670 4868 4726 4924
rect 4726 4868 4730 4924
rect 4666 4864 4730 4868
rect 4746 4924 4810 4928
rect 4746 4868 4750 4924
rect 4750 4868 4806 4924
rect 4806 4868 4810 4924
rect 4746 4864 4810 4868
rect 4826 4924 4890 4928
rect 4826 4868 4830 4924
rect 4830 4868 4886 4924
rect 4886 4868 4890 4924
rect 4826 4864 4890 4868
rect 4906 4924 4970 4928
rect 4906 4868 4910 4924
rect 4910 4868 4966 4924
rect 4966 4868 4970 4924
rect 4906 4864 4970 4868
rect 12094 4924 12158 4928
rect 12094 4868 12098 4924
rect 12098 4868 12154 4924
rect 12154 4868 12158 4924
rect 12094 4864 12158 4868
rect 12174 4924 12238 4928
rect 12174 4868 12178 4924
rect 12178 4868 12234 4924
rect 12234 4868 12238 4924
rect 12174 4864 12238 4868
rect 12254 4924 12318 4928
rect 12254 4868 12258 4924
rect 12258 4868 12314 4924
rect 12314 4868 12318 4924
rect 12254 4864 12318 4868
rect 12334 4924 12398 4928
rect 12334 4868 12338 4924
rect 12338 4868 12394 4924
rect 12394 4868 12398 4924
rect 12334 4864 12398 4868
rect 19522 4924 19586 4928
rect 19522 4868 19526 4924
rect 19526 4868 19582 4924
rect 19582 4868 19586 4924
rect 19522 4864 19586 4868
rect 19602 4924 19666 4928
rect 19602 4868 19606 4924
rect 19606 4868 19662 4924
rect 19662 4868 19666 4924
rect 19602 4864 19666 4868
rect 19682 4924 19746 4928
rect 19682 4868 19686 4924
rect 19686 4868 19742 4924
rect 19742 4868 19746 4924
rect 19682 4864 19746 4868
rect 19762 4924 19826 4928
rect 19762 4868 19766 4924
rect 19766 4868 19822 4924
rect 19822 4868 19826 4924
rect 19762 4864 19826 4868
rect 26950 4924 27014 4928
rect 26950 4868 26954 4924
rect 26954 4868 27010 4924
rect 27010 4868 27014 4924
rect 26950 4864 27014 4868
rect 27030 4924 27094 4928
rect 27030 4868 27034 4924
rect 27034 4868 27090 4924
rect 27090 4868 27094 4924
rect 27030 4864 27094 4868
rect 27110 4924 27174 4928
rect 27110 4868 27114 4924
rect 27114 4868 27170 4924
rect 27170 4868 27174 4924
rect 27110 4864 27174 4868
rect 27190 4924 27254 4928
rect 27190 4868 27194 4924
rect 27194 4868 27250 4924
rect 27250 4868 27254 4924
rect 27190 4864 27254 4868
rect 8380 4380 8444 4384
rect 8380 4324 8384 4380
rect 8384 4324 8440 4380
rect 8440 4324 8444 4380
rect 8380 4320 8444 4324
rect 8460 4380 8524 4384
rect 8460 4324 8464 4380
rect 8464 4324 8520 4380
rect 8520 4324 8524 4380
rect 8460 4320 8524 4324
rect 8540 4380 8604 4384
rect 8540 4324 8544 4380
rect 8544 4324 8600 4380
rect 8600 4324 8604 4380
rect 8540 4320 8604 4324
rect 8620 4380 8684 4384
rect 8620 4324 8624 4380
rect 8624 4324 8680 4380
rect 8680 4324 8684 4380
rect 8620 4320 8684 4324
rect 15808 4380 15872 4384
rect 15808 4324 15812 4380
rect 15812 4324 15868 4380
rect 15868 4324 15872 4380
rect 15808 4320 15872 4324
rect 15888 4380 15952 4384
rect 15888 4324 15892 4380
rect 15892 4324 15948 4380
rect 15948 4324 15952 4380
rect 15888 4320 15952 4324
rect 15968 4380 16032 4384
rect 15968 4324 15972 4380
rect 15972 4324 16028 4380
rect 16028 4324 16032 4380
rect 15968 4320 16032 4324
rect 16048 4380 16112 4384
rect 16048 4324 16052 4380
rect 16052 4324 16108 4380
rect 16108 4324 16112 4380
rect 16048 4320 16112 4324
rect 23236 4380 23300 4384
rect 23236 4324 23240 4380
rect 23240 4324 23296 4380
rect 23296 4324 23300 4380
rect 23236 4320 23300 4324
rect 23316 4380 23380 4384
rect 23316 4324 23320 4380
rect 23320 4324 23376 4380
rect 23376 4324 23380 4380
rect 23316 4320 23380 4324
rect 23396 4380 23460 4384
rect 23396 4324 23400 4380
rect 23400 4324 23456 4380
rect 23456 4324 23460 4380
rect 23396 4320 23460 4324
rect 23476 4380 23540 4384
rect 23476 4324 23480 4380
rect 23480 4324 23536 4380
rect 23536 4324 23540 4380
rect 23476 4320 23540 4324
rect 30664 4380 30728 4384
rect 30664 4324 30668 4380
rect 30668 4324 30724 4380
rect 30724 4324 30728 4380
rect 30664 4320 30728 4324
rect 30744 4380 30808 4384
rect 30744 4324 30748 4380
rect 30748 4324 30804 4380
rect 30804 4324 30808 4380
rect 30744 4320 30808 4324
rect 30824 4380 30888 4384
rect 30824 4324 30828 4380
rect 30828 4324 30884 4380
rect 30884 4324 30888 4380
rect 30824 4320 30888 4324
rect 30904 4380 30968 4384
rect 30904 4324 30908 4380
rect 30908 4324 30964 4380
rect 30964 4324 30968 4380
rect 30904 4320 30968 4324
rect 4666 3836 4730 3840
rect 4666 3780 4670 3836
rect 4670 3780 4726 3836
rect 4726 3780 4730 3836
rect 4666 3776 4730 3780
rect 4746 3836 4810 3840
rect 4746 3780 4750 3836
rect 4750 3780 4806 3836
rect 4806 3780 4810 3836
rect 4746 3776 4810 3780
rect 4826 3836 4890 3840
rect 4826 3780 4830 3836
rect 4830 3780 4886 3836
rect 4886 3780 4890 3836
rect 4826 3776 4890 3780
rect 4906 3836 4970 3840
rect 4906 3780 4910 3836
rect 4910 3780 4966 3836
rect 4966 3780 4970 3836
rect 4906 3776 4970 3780
rect 12094 3836 12158 3840
rect 12094 3780 12098 3836
rect 12098 3780 12154 3836
rect 12154 3780 12158 3836
rect 12094 3776 12158 3780
rect 12174 3836 12238 3840
rect 12174 3780 12178 3836
rect 12178 3780 12234 3836
rect 12234 3780 12238 3836
rect 12174 3776 12238 3780
rect 12254 3836 12318 3840
rect 12254 3780 12258 3836
rect 12258 3780 12314 3836
rect 12314 3780 12318 3836
rect 12254 3776 12318 3780
rect 12334 3836 12398 3840
rect 12334 3780 12338 3836
rect 12338 3780 12394 3836
rect 12394 3780 12398 3836
rect 12334 3776 12398 3780
rect 19522 3836 19586 3840
rect 19522 3780 19526 3836
rect 19526 3780 19582 3836
rect 19582 3780 19586 3836
rect 19522 3776 19586 3780
rect 19602 3836 19666 3840
rect 19602 3780 19606 3836
rect 19606 3780 19662 3836
rect 19662 3780 19666 3836
rect 19602 3776 19666 3780
rect 19682 3836 19746 3840
rect 19682 3780 19686 3836
rect 19686 3780 19742 3836
rect 19742 3780 19746 3836
rect 19682 3776 19746 3780
rect 19762 3836 19826 3840
rect 19762 3780 19766 3836
rect 19766 3780 19822 3836
rect 19822 3780 19826 3836
rect 19762 3776 19826 3780
rect 26950 3836 27014 3840
rect 26950 3780 26954 3836
rect 26954 3780 27010 3836
rect 27010 3780 27014 3836
rect 26950 3776 27014 3780
rect 27030 3836 27094 3840
rect 27030 3780 27034 3836
rect 27034 3780 27090 3836
rect 27090 3780 27094 3836
rect 27030 3776 27094 3780
rect 27110 3836 27174 3840
rect 27110 3780 27114 3836
rect 27114 3780 27170 3836
rect 27170 3780 27174 3836
rect 27110 3776 27174 3780
rect 27190 3836 27254 3840
rect 27190 3780 27194 3836
rect 27194 3780 27250 3836
rect 27250 3780 27254 3836
rect 27190 3776 27254 3780
rect 8380 3292 8444 3296
rect 8380 3236 8384 3292
rect 8384 3236 8440 3292
rect 8440 3236 8444 3292
rect 8380 3232 8444 3236
rect 8460 3292 8524 3296
rect 8460 3236 8464 3292
rect 8464 3236 8520 3292
rect 8520 3236 8524 3292
rect 8460 3232 8524 3236
rect 8540 3292 8604 3296
rect 8540 3236 8544 3292
rect 8544 3236 8600 3292
rect 8600 3236 8604 3292
rect 8540 3232 8604 3236
rect 8620 3292 8684 3296
rect 8620 3236 8624 3292
rect 8624 3236 8680 3292
rect 8680 3236 8684 3292
rect 8620 3232 8684 3236
rect 15808 3292 15872 3296
rect 15808 3236 15812 3292
rect 15812 3236 15868 3292
rect 15868 3236 15872 3292
rect 15808 3232 15872 3236
rect 15888 3292 15952 3296
rect 15888 3236 15892 3292
rect 15892 3236 15948 3292
rect 15948 3236 15952 3292
rect 15888 3232 15952 3236
rect 15968 3292 16032 3296
rect 15968 3236 15972 3292
rect 15972 3236 16028 3292
rect 16028 3236 16032 3292
rect 15968 3232 16032 3236
rect 16048 3292 16112 3296
rect 16048 3236 16052 3292
rect 16052 3236 16108 3292
rect 16108 3236 16112 3292
rect 16048 3232 16112 3236
rect 23236 3292 23300 3296
rect 23236 3236 23240 3292
rect 23240 3236 23296 3292
rect 23296 3236 23300 3292
rect 23236 3232 23300 3236
rect 23316 3292 23380 3296
rect 23316 3236 23320 3292
rect 23320 3236 23376 3292
rect 23376 3236 23380 3292
rect 23316 3232 23380 3236
rect 23396 3292 23460 3296
rect 23396 3236 23400 3292
rect 23400 3236 23456 3292
rect 23456 3236 23460 3292
rect 23396 3232 23460 3236
rect 23476 3292 23540 3296
rect 23476 3236 23480 3292
rect 23480 3236 23536 3292
rect 23536 3236 23540 3292
rect 23476 3232 23540 3236
rect 30664 3292 30728 3296
rect 30664 3236 30668 3292
rect 30668 3236 30724 3292
rect 30724 3236 30728 3292
rect 30664 3232 30728 3236
rect 30744 3292 30808 3296
rect 30744 3236 30748 3292
rect 30748 3236 30804 3292
rect 30804 3236 30808 3292
rect 30744 3232 30808 3236
rect 30824 3292 30888 3296
rect 30824 3236 30828 3292
rect 30828 3236 30884 3292
rect 30884 3236 30888 3292
rect 30824 3232 30888 3236
rect 30904 3292 30968 3296
rect 30904 3236 30908 3292
rect 30908 3236 30964 3292
rect 30964 3236 30968 3292
rect 30904 3232 30968 3236
rect 4666 2748 4730 2752
rect 4666 2692 4670 2748
rect 4670 2692 4726 2748
rect 4726 2692 4730 2748
rect 4666 2688 4730 2692
rect 4746 2748 4810 2752
rect 4746 2692 4750 2748
rect 4750 2692 4806 2748
rect 4806 2692 4810 2748
rect 4746 2688 4810 2692
rect 4826 2748 4890 2752
rect 4826 2692 4830 2748
rect 4830 2692 4886 2748
rect 4886 2692 4890 2748
rect 4826 2688 4890 2692
rect 4906 2748 4970 2752
rect 4906 2692 4910 2748
rect 4910 2692 4966 2748
rect 4966 2692 4970 2748
rect 4906 2688 4970 2692
rect 12094 2748 12158 2752
rect 12094 2692 12098 2748
rect 12098 2692 12154 2748
rect 12154 2692 12158 2748
rect 12094 2688 12158 2692
rect 12174 2748 12238 2752
rect 12174 2692 12178 2748
rect 12178 2692 12234 2748
rect 12234 2692 12238 2748
rect 12174 2688 12238 2692
rect 12254 2748 12318 2752
rect 12254 2692 12258 2748
rect 12258 2692 12314 2748
rect 12314 2692 12318 2748
rect 12254 2688 12318 2692
rect 12334 2748 12398 2752
rect 12334 2692 12338 2748
rect 12338 2692 12394 2748
rect 12394 2692 12398 2748
rect 12334 2688 12398 2692
rect 19522 2748 19586 2752
rect 19522 2692 19526 2748
rect 19526 2692 19582 2748
rect 19582 2692 19586 2748
rect 19522 2688 19586 2692
rect 19602 2748 19666 2752
rect 19602 2692 19606 2748
rect 19606 2692 19662 2748
rect 19662 2692 19666 2748
rect 19602 2688 19666 2692
rect 19682 2748 19746 2752
rect 19682 2692 19686 2748
rect 19686 2692 19742 2748
rect 19742 2692 19746 2748
rect 19682 2688 19746 2692
rect 19762 2748 19826 2752
rect 19762 2692 19766 2748
rect 19766 2692 19822 2748
rect 19822 2692 19826 2748
rect 19762 2688 19826 2692
rect 26950 2748 27014 2752
rect 26950 2692 26954 2748
rect 26954 2692 27010 2748
rect 27010 2692 27014 2748
rect 26950 2688 27014 2692
rect 27030 2748 27094 2752
rect 27030 2692 27034 2748
rect 27034 2692 27090 2748
rect 27090 2692 27094 2748
rect 27030 2688 27094 2692
rect 27110 2748 27174 2752
rect 27110 2692 27114 2748
rect 27114 2692 27170 2748
rect 27170 2692 27174 2748
rect 27110 2688 27174 2692
rect 27190 2748 27254 2752
rect 27190 2692 27194 2748
rect 27194 2692 27250 2748
rect 27250 2692 27254 2748
rect 27190 2688 27254 2692
rect 8380 2204 8444 2208
rect 8380 2148 8384 2204
rect 8384 2148 8440 2204
rect 8440 2148 8444 2204
rect 8380 2144 8444 2148
rect 8460 2204 8524 2208
rect 8460 2148 8464 2204
rect 8464 2148 8520 2204
rect 8520 2148 8524 2204
rect 8460 2144 8524 2148
rect 8540 2204 8604 2208
rect 8540 2148 8544 2204
rect 8544 2148 8600 2204
rect 8600 2148 8604 2204
rect 8540 2144 8604 2148
rect 8620 2204 8684 2208
rect 8620 2148 8624 2204
rect 8624 2148 8680 2204
rect 8680 2148 8684 2204
rect 8620 2144 8684 2148
rect 15808 2204 15872 2208
rect 15808 2148 15812 2204
rect 15812 2148 15868 2204
rect 15868 2148 15872 2204
rect 15808 2144 15872 2148
rect 15888 2204 15952 2208
rect 15888 2148 15892 2204
rect 15892 2148 15948 2204
rect 15948 2148 15952 2204
rect 15888 2144 15952 2148
rect 15968 2204 16032 2208
rect 15968 2148 15972 2204
rect 15972 2148 16028 2204
rect 16028 2148 16032 2204
rect 15968 2144 16032 2148
rect 16048 2204 16112 2208
rect 16048 2148 16052 2204
rect 16052 2148 16108 2204
rect 16108 2148 16112 2204
rect 16048 2144 16112 2148
rect 23236 2204 23300 2208
rect 23236 2148 23240 2204
rect 23240 2148 23296 2204
rect 23296 2148 23300 2204
rect 23236 2144 23300 2148
rect 23316 2204 23380 2208
rect 23316 2148 23320 2204
rect 23320 2148 23376 2204
rect 23376 2148 23380 2204
rect 23316 2144 23380 2148
rect 23396 2204 23460 2208
rect 23396 2148 23400 2204
rect 23400 2148 23456 2204
rect 23456 2148 23460 2204
rect 23396 2144 23460 2148
rect 23476 2204 23540 2208
rect 23476 2148 23480 2204
rect 23480 2148 23536 2204
rect 23536 2148 23540 2204
rect 23476 2144 23540 2148
rect 30664 2204 30728 2208
rect 30664 2148 30668 2204
rect 30668 2148 30724 2204
rect 30724 2148 30728 2204
rect 30664 2144 30728 2148
rect 30744 2204 30808 2208
rect 30744 2148 30748 2204
rect 30748 2148 30804 2204
rect 30804 2148 30808 2204
rect 30744 2144 30808 2148
rect 30824 2204 30888 2208
rect 30824 2148 30828 2204
rect 30828 2148 30884 2204
rect 30884 2148 30888 2204
rect 30824 2144 30888 2148
rect 30904 2204 30968 2208
rect 30904 2148 30908 2204
rect 30908 2148 30964 2204
rect 30964 2148 30968 2204
rect 30904 2144 30968 2148
<< metal4 >>
rect 4658 28864 4978 29424
rect 4658 28800 4666 28864
rect 4730 28800 4746 28864
rect 4810 28800 4826 28864
rect 4890 28800 4906 28864
rect 4970 28800 4978 28864
rect 4658 27776 4978 28800
rect 4658 27712 4666 27776
rect 4730 27712 4746 27776
rect 4810 27712 4826 27776
rect 4890 27712 4906 27776
rect 4970 27712 4978 27776
rect 4658 26688 4978 27712
rect 4658 26624 4666 26688
rect 4730 26624 4746 26688
rect 4810 26624 4826 26688
rect 4890 26624 4906 26688
rect 4970 26624 4978 26688
rect 4658 25600 4978 26624
rect 4658 25536 4666 25600
rect 4730 25536 4746 25600
rect 4810 25536 4826 25600
rect 4890 25536 4906 25600
rect 4970 25536 4978 25600
rect 4658 24512 4978 25536
rect 4658 24448 4666 24512
rect 4730 24448 4746 24512
rect 4810 24448 4826 24512
rect 4890 24448 4906 24512
rect 4970 24448 4978 24512
rect 4658 23424 4978 24448
rect 4658 23360 4666 23424
rect 4730 23360 4746 23424
rect 4810 23360 4826 23424
rect 4890 23360 4906 23424
rect 4970 23360 4978 23424
rect 4658 22336 4978 23360
rect 4658 22272 4666 22336
rect 4730 22272 4746 22336
rect 4810 22272 4826 22336
rect 4890 22272 4906 22336
rect 4970 22272 4978 22336
rect 4658 21248 4978 22272
rect 4658 21184 4666 21248
rect 4730 21184 4746 21248
rect 4810 21184 4826 21248
rect 4890 21184 4906 21248
rect 4970 21184 4978 21248
rect 4658 20160 4978 21184
rect 4658 20096 4666 20160
rect 4730 20096 4746 20160
rect 4810 20096 4826 20160
rect 4890 20096 4906 20160
rect 4970 20096 4978 20160
rect 4658 19072 4978 20096
rect 4658 19008 4666 19072
rect 4730 19008 4746 19072
rect 4810 19008 4826 19072
rect 4890 19008 4906 19072
rect 4970 19008 4978 19072
rect 4658 17984 4978 19008
rect 4658 17920 4666 17984
rect 4730 17920 4746 17984
rect 4810 17920 4826 17984
rect 4890 17920 4906 17984
rect 4970 17920 4978 17984
rect 4658 16896 4978 17920
rect 4658 16832 4666 16896
rect 4730 16832 4746 16896
rect 4810 16832 4826 16896
rect 4890 16832 4906 16896
rect 4970 16832 4978 16896
rect 4658 15808 4978 16832
rect 4658 15744 4666 15808
rect 4730 15744 4746 15808
rect 4810 15744 4826 15808
rect 4890 15744 4906 15808
rect 4970 15744 4978 15808
rect 4658 14720 4978 15744
rect 4658 14656 4666 14720
rect 4730 14656 4746 14720
rect 4810 14656 4826 14720
rect 4890 14656 4906 14720
rect 4970 14656 4978 14720
rect 4658 13632 4978 14656
rect 4658 13568 4666 13632
rect 4730 13568 4746 13632
rect 4810 13568 4826 13632
rect 4890 13568 4906 13632
rect 4970 13568 4978 13632
rect 4658 12544 4978 13568
rect 4658 12480 4666 12544
rect 4730 12480 4746 12544
rect 4810 12480 4826 12544
rect 4890 12480 4906 12544
rect 4970 12480 4978 12544
rect 4658 11456 4978 12480
rect 4658 11392 4666 11456
rect 4730 11392 4746 11456
rect 4810 11392 4826 11456
rect 4890 11392 4906 11456
rect 4970 11392 4978 11456
rect 4658 10368 4978 11392
rect 4658 10304 4666 10368
rect 4730 10304 4746 10368
rect 4810 10304 4826 10368
rect 4890 10304 4906 10368
rect 4970 10304 4978 10368
rect 4658 9280 4978 10304
rect 4658 9216 4666 9280
rect 4730 9216 4746 9280
rect 4810 9216 4826 9280
rect 4890 9216 4906 9280
rect 4970 9216 4978 9280
rect 4658 8192 4978 9216
rect 4658 8128 4666 8192
rect 4730 8128 4746 8192
rect 4810 8128 4826 8192
rect 4890 8128 4906 8192
rect 4970 8128 4978 8192
rect 4658 7104 4978 8128
rect 4658 7040 4666 7104
rect 4730 7040 4746 7104
rect 4810 7040 4826 7104
rect 4890 7040 4906 7104
rect 4970 7040 4978 7104
rect 4658 6016 4978 7040
rect 4658 5952 4666 6016
rect 4730 5952 4746 6016
rect 4810 5952 4826 6016
rect 4890 5952 4906 6016
rect 4970 5952 4978 6016
rect 4658 4928 4978 5952
rect 4658 4864 4666 4928
rect 4730 4864 4746 4928
rect 4810 4864 4826 4928
rect 4890 4864 4906 4928
rect 4970 4864 4978 4928
rect 4658 3840 4978 4864
rect 4658 3776 4666 3840
rect 4730 3776 4746 3840
rect 4810 3776 4826 3840
rect 4890 3776 4906 3840
rect 4970 3776 4978 3840
rect 4658 2752 4978 3776
rect 4658 2688 4666 2752
rect 4730 2688 4746 2752
rect 4810 2688 4826 2752
rect 4890 2688 4906 2752
rect 4970 2688 4978 2752
rect 4658 2128 4978 2688
rect 8372 29408 8692 29424
rect 8372 29344 8380 29408
rect 8444 29344 8460 29408
rect 8524 29344 8540 29408
rect 8604 29344 8620 29408
rect 8684 29344 8692 29408
rect 8372 28320 8692 29344
rect 8372 28256 8380 28320
rect 8444 28256 8460 28320
rect 8524 28256 8540 28320
rect 8604 28256 8620 28320
rect 8684 28256 8692 28320
rect 8372 27232 8692 28256
rect 8372 27168 8380 27232
rect 8444 27168 8460 27232
rect 8524 27168 8540 27232
rect 8604 27168 8620 27232
rect 8684 27168 8692 27232
rect 8372 26144 8692 27168
rect 8372 26080 8380 26144
rect 8444 26080 8460 26144
rect 8524 26080 8540 26144
rect 8604 26080 8620 26144
rect 8684 26080 8692 26144
rect 8372 25056 8692 26080
rect 8372 24992 8380 25056
rect 8444 24992 8460 25056
rect 8524 24992 8540 25056
rect 8604 24992 8620 25056
rect 8684 24992 8692 25056
rect 8372 23968 8692 24992
rect 8372 23904 8380 23968
rect 8444 23904 8460 23968
rect 8524 23904 8540 23968
rect 8604 23904 8620 23968
rect 8684 23904 8692 23968
rect 8372 22880 8692 23904
rect 8372 22816 8380 22880
rect 8444 22816 8460 22880
rect 8524 22816 8540 22880
rect 8604 22816 8620 22880
rect 8684 22816 8692 22880
rect 8372 21792 8692 22816
rect 8372 21728 8380 21792
rect 8444 21728 8460 21792
rect 8524 21728 8540 21792
rect 8604 21728 8620 21792
rect 8684 21728 8692 21792
rect 8372 20704 8692 21728
rect 8372 20640 8380 20704
rect 8444 20640 8460 20704
rect 8524 20640 8540 20704
rect 8604 20640 8620 20704
rect 8684 20640 8692 20704
rect 8372 19616 8692 20640
rect 8372 19552 8380 19616
rect 8444 19552 8460 19616
rect 8524 19552 8540 19616
rect 8604 19552 8620 19616
rect 8684 19552 8692 19616
rect 8372 18528 8692 19552
rect 8372 18464 8380 18528
rect 8444 18464 8460 18528
rect 8524 18464 8540 18528
rect 8604 18464 8620 18528
rect 8684 18464 8692 18528
rect 8372 17440 8692 18464
rect 8372 17376 8380 17440
rect 8444 17376 8460 17440
rect 8524 17376 8540 17440
rect 8604 17376 8620 17440
rect 8684 17376 8692 17440
rect 8372 16352 8692 17376
rect 8372 16288 8380 16352
rect 8444 16288 8460 16352
rect 8524 16288 8540 16352
rect 8604 16288 8620 16352
rect 8684 16288 8692 16352
rect 8372 15264 8692 16288
rect 8372 15200 8380 15264
rect 8444 15200 8460 15264
rect 8524 15200 8540 15264
rect 8604 15200 8620 15264
rect 8684 15200 8692 15264
rect 8372 14176 8692 15200
rect 8372 14112 8380 14176
rect 8444 14112 8460 14176
rect 8524 14112 8540 14176
rect 8604 14112 8620 14176
rect 8684 14112 8692 14176
rect 8372 13088 8692 14112
rect 8372 13024 8380 13088
rect 8444 13024 8460 13088
rect 8524 13024 8540 13088
rect 8604 13024 8620 13088
rect 8684 13024 8692 13088
rect 8372 12000 8692 13024
rect 8372 11936 8380 12000
rect 8444 11936 8460 12000
rect 8524 11936 8540 12000
rect 8604 11936 8620 12000
rect 8684 11936 8692 12000
rect 8372 10912 8692 11936
rect 8372 10848 8380 10912
rect 8444 10848 8460 10912
rect 8524 10848 8540 10912
rect 8604 10848 8620 10912
rect 8684 10848 8692 10912
rect 8372 9824 8692 10848
rect 8372 9760 8380 9824
rect 8444 9760 8460 9824
rect 8524 9760 8540 9824
rect 8604 9760 8620 9824
rect 8684 9760 8692 9824
rect 8372 8736 8692 9760
rect 8372 8672 8380 8736
rect 8444 8672 8460 8736
rect 8524 8672 8540 8736
rect 8604 8672 8620 8736
rect 8684 8672 8692 8736
rect 8372 7648 8692 8672
rect 8372 7584 8380 7648
rect 8444 7584 8460 7648
rect 8524 7584 8540 7648
rect 8604 7584 8620 7648
rect 8684 7584 8692 7648
rect 8372 6560 8692 7584
rect 8372 6496 8380 6560
rect 8444 6496 8460 6560
rect 8524 6496 8540 6560
rect 8604 6496 8620 6560
rect 8684 6496 8692 6560
rect 8372 5472 8692 6496
rect 8372 5408 8380 5472
rect 8444 5408 8460 5472
rect 8524 5408 8540 5472
rect 8604 5408 8620 5472
rect 8684 5408 8692 5472
rect 8372 4384 8692 5408
rect 8372 4320 8380 4384
rect 8444 4320 8460 4384
rect 8524 4320 8540 4384
rect 8604 4320 8620 4384
rect 8684 4320 8692 4384
rect 8372 3296 8692 4320
rect 8372 3232 8380 3296
rect 8444 3232 8460 3296
rect 8524 3232 8540 3296
rect 8604 3232 8620 3296
rect 8684 3232 8692 3296
rect 8372 2208 8692 3232
rect 8372 2144 8380 2208
rect 8444 2144 8460 2208
rect 8524 2144 8540 2208
rect 8604 2144 8620 2208
rect 8684 2144 8692 2208
rect 8372 2128 8692 2144
rect 12086 28864 12406 29424
rect 12086 28800 12094 28864
rect 12158 28800 12174 28864
rect 12238 28800 12254 28864
rect 12318 28800 12334 28864
rect 12398 28800 12406 28864
rect 12086 27776 12406 28800
rect 12086 27712 12094 27776
rect 12158 27712 12174 27776
rect 12238 27712 12254 27776
rect 12318 27712 12334 27776
rect 12398 27712 12406 27776
rect 12086 26688 12406 27712
rect 12086 26624 12094 26688
rect 12158 26624 12174 26688
rect 12238 26624 12254 26688
rect 12318 26624 12334 26688
rect 12398 26624 12406 26688
rect 12086 25600 12406 26624
rect 12086 25536 12094 25600
rect 12158 25536 12174 25600
rect 12238 25536 12254 25600
rect 12318 25536 12334 25600
rect 12398 25536 12406 25600
rect 12086 24512 12406 25536
rect 12086 24448 12094 24512
rect 12158 24448 12174 24512
rect 12238 24448 12254 24512
rect 12318 24448 12334 24512
rect 12398 24448 12406 24512
rect 12086 23424 12406 24448
rect 12086 23360 12094 23424
rect 12158 23360 12174 23424
rect 12238 23360 12254 23424
rect 12318 23360 12334 23424
rect 12398 23360 12406 23424
rect 12086 22336 12406 23360
rect 12086 22272 12094 22336
rect 12158 22272 12174 22336
rect 12238 22272 12254 22336
rect 12318 22272 12334 22336
rect 12398 22272 12406 22336
rect 12086 21248 12406 22272
rect 12086 21184 12094 21248
rect 12158 21184 12174 21248
rect 12238 21184 12254 21248
rect 12318 21184 12334 21248
rect 12398 21184 12406 21248
rect 12086 20160 12406 21184
rect 12086 20096 12094 20160
rect 12158 20096 12174 20160
rect 12238 20096 12254 20160
rect 12318 20096 12334 20160
rect 12398 20096 12406 20160
rect 12086 19072 12406 20096
rect 12086 19008 12094 19072
rect 12158 19008 12174 19072
rect 12238 19008 12254 19072
rect 12318 19008 12334 19072
rect 12398 19008 12406 19072
rect 12086 17984 12406 19008
rect 12086 17920 12094 17984
rect 12158 17920 12174 17984
rect 12238 17920 12254 17984
rect 12318 17920 12334 17984
rect 12398 17920 12406 17984
rect 12086 16896 12406 17920
rect 12086 16832 12094 16896
rect 12158 16832 12174 16896
rect 12238 16832 12254 16896
rect 12318 16832 12334 16896
rect 12398 16832 12406 16896
rect 12086 15808 12406 16832
rect 12086 15744 12094 15808
rect 12158 15744 12174 15808
rect 12238 15744 12254 15808
rect 12318 15744 12334 15808
rect 12398 15744 12406 15808
rect 12086 14720 12406 15744
rect 12086 14656 12094 14720
rect 12158 14656 12174 14720
rect 12238 14656 12254 14720
rect 12318 14656 12334 14720
rect 12398 14656 12406 14720
rect 12086 13632 12406 14656
rect 12086 13568 12094 13632
rect 12158 13568 12174 13632
rect 12238 13568 12254 13632
rect 12318 13568 12334 13632
rect 12398 13568 12406 13632
rect 12086 12544 12406 13568
rect 12086 12480 12094 12544
rect 12158 12480 12174 12544
rect 12238 12480 12254 12544
rect 12318 12480 12334 12544
rect 12398 12480 12406 12544
rect 12086 11456 12406 12480
rect 12086 11392 12094 11456
rect 12158 11392 12174 11456
rect 12238 11392 12254 11456
rect 12318 11392 12334 11456
rect 12398 11392 12406 11456
rect 12086 10368 12406 11392
rect 12086 10304 12094 10368
rect 12158 10304 12174 10368
rect 12238 10304 12254 10368
rect 12318 10304 12334 10368
rect 12398 10304 12406 10368
rect 12086 9280 12406 10304
rect 12086 9216 12094 9280
rect 12158 9216 12174 9280
rect 12238 9216 12254 9280
rect 12318 9216 12334 9280
rect 12398 9216 12406 9280
rect 12086 8192 12406 9216
rect 12086 8128 12094 8192
rect 12158 8128 12174 8192
rect 12238 8128 12254 8192
rect 12318 8128 12334 8192
rect 12398 8128 12406 8192
rect 12086 7104 12406 8128
rect 12086 7040 12094 7104
rect 12158 7040 12174 7104
rect 12238 7040 12254 7104
rect 12318 7040 12334 7104
rect 12398 7040 12406 7104
rect 12086 6016 12406 7040
rect 12086 5952 12094 6016
rect 12158 5952 12174 6016
rect 12238 5952 12254 6016
rect 12318 5952 12334 6016
rect 12398 5952 12406 6016
rect 12086 4928 12406 5952
rect 12086 4864 12094 4928
rect 12158 4864 12174 4928
rect 12238 4864 12254 4928
rect 12318 4864 12334 4928
rect 12398 4864 12406 4928
rect 12086 3840 12406 4864
rect 12086 3776 12094 3840
rect 12158 3776 12174 3840
rect 12238 3776 12254 3840
rect 12318 3776 12334 3840
rect 12398 3776 12406 3840
rect 12086 2752 12406 3776
rect 12086 2688 12094 2752
rect 12158 2688 12174 2752
rect 12238 2688 12254 2752
rect 12318 2688 12334 2752
rect 12398 2688 12406 2752
rect 12086 2128 12406 2688
rect 15800 29408 16120 29424
rect 15800 29344 15808 29408
rect 15872 29344 15888 29408
rect 15952 29344 15968 29408
rect 16032 29344 16048 29408
rect 16112 29344 16120 29408
rect 15800 28320 16120 29344
rect 15800 28256 15808 28320
rect 15872 28256 15888 28320
rect 15952 28256 15968 28320
rect 16032 28256 16048 28320
rect 16112 28256 16120 28320
rect 15800 27232 16120 28256
rect 15800 27168 15808 27232
rect 15872 27168 15888 27232
rect 15952 27168 15968 27232
rect 16032 27168 16048 27232
rect 16112 27168 16120 27232
rect 15800 26144 16120 27168
rect 15800 26080 15808 26144
rect 15872 26080 15888 26144
rect 15952 26080 15968 26144
rect 16032 26080 16048 26144
rect 16112 26080 16120 26144
rect 15800 25056 16120 26080
rect 15800 24992 15808 25056
rect 15872 24992 15888 25056
rect 15952 24992 15968 25056
rect 16032 24992 16048 25056
rect 16112 24992 16120 25056
rect 15800 23968 16120 24992
rect 15800 23904 15808 23968
rect 15872 23904 15888 23968
rect 15952 23904 15968 23968
rect 16032 23904 16048 23968
rect 16112 23904 16120 23968
rect 15800 22880 16120 23904
rect 15800 22816 15808 22880
rect 15872 22816 15888 22880
rect 15952 22816 15968 22880
rect 16032 22816 16048 22880
rect 16112 22816 16120 22880
rect 15800 21792 16120 22816
rect 15800 21728 15808 21792
rect 15872 21728 15888 21792
rect 15952 21728 15968 21792
rect 16032 21728 16048 21792
rect 16112 21728 16120 21792
rect 15800 20704 16120 21728
rect 15800 20640 15808 20704
rect 15872 20640 15888 20704
rect 15952 20640 15968 20704
rect 16032 20640 16048 20704
rect 16112 20640 16120 20704
rect 15800 19616 16120 20640
rect 15800 19552 15808 19616
rect 15872 19552 15888 19616
rect 15952 19552 15968 19616
rect 16032 19552 16048 19616
rect 16112 19552 16120 19616
rect 15800 18528 16120 19552
rect 15800 18464 15808 18528
rect 15872 18464 15888 18528
rect 15952 18464 15968 18528
rect 16032 18464 16048 18528
rect 16112 18464 16120 18528
rect 15800 17440 16120 18464
rect 15800 17376 15808 17440
rect 15872 17376 15888 17440
rect 15952 17376 15968 17440
rect 16032 17376 16048 17440
rect 16112 17376 16120 17440
rect 15800 16352 16120 17376
rect 15800 16288 15808 16352
rect 15872 16288 15888 16352
rect 15952 16288 15968 16352
rect 16032 16288 16048 16352
rect 16112 16288 16120 16352
rect 15800 15264 16120 16288
rect 15800 15200 15808 15264
rect 15872 15200 15888 15264
rect 15952 15200 15968 15264
rect 16032 15200 16048 15264
rect 16112 15200 16120 15264
rect 15800 14176 16120 15200
rect 15800 14112 15808 14176
rect 15872 14112 15888 14176
rect 15952 14112 15968 14176
rect 16032 14112 16048 14176
rect 16112 14112 16120 14176
rect 15800 13088 16120 14112
rect 15800 13024 15808 13088
rect 15872 13024 15888 13088
rect 15952 13024 15968 13088
rect 16032 13024 16048 13088
rect 16112 13024 16120 13088
rect 15800 12000 16120 13024
rect 15800 11936 15808 12000
rect 15872 11936 15888 12000
rect 15952 11936 15968 12000
rect 16032 11936 16048 12000
rect 16112 11936 16120 12000
rect 15800 10912 16120 11936
rect 15800 10848 15808 10912
rect 15872 10848 15888 10912
rect 15952 10848 15968 10912
rect 16032 10848 16048 10912
rect 16112 10848 16120 10912
rect 15800 9824 16120 10848
rect 15800 9760 15808 9824
rect 15872 9760 15888 9824
rect 15952 9760 15968 9824
rect 16032 9760 16048 9824
rect 16112 9760 16120 9824
rect 15800 8736 16120 9760
rect 15800 8672 15808 8736
rect 15872 8672 15888 8736
rect 15952 8672 15968 8736
rect 16032 8672 16048 8736
rect 16112 8672 16120 8736
rect 15800 7648 16120 8672
rect 15800 7584 15808 7648
rect 15872 7584 15888 7648
rect 15952 7584 15968 7648
rect 16032 7584 16048 7648
rect 16112 7584 16120 7648
rect 15800 6560 16120 7584
rect 15800 6496 15808 6560
rect 15872 6496 15888 6560
rect 15952 6496 15968 6560
rect 16032 6496 16048 6560
rect 16112 6496 16120 6560
rect 15800 5472 16120 6496
rect 15800 5408 15808 5472
rect 15872 5408 15888 5472
rect 15952 5408 15968 5472
rect 16032 5408 16048 5472
rect 16112 5408 16120 5472
rect 15800 4384 16120 5408
rect 15800 4320 15808 4384
rect 15872 4320 15888 4384
rect 15952 4320 15968 4384
rect 16032 4320 16048 4384
rect 16112 4320 16120 4384
rect 15800 3296 16120 4320
rect 15800 3232 15808 3296
rect 15872 3232 15888 3296
rect 15952 3232 15968 3296
rect 16032 3232 16048 3296
rect 16112 3232 16120 3296
rect 15800 2208 16120 3232
rect 15800 2144 15808 2208
rect 15872 2144 15888 2208
rect 15952 2144 15968 2208
rect 16032 2144 16048 2208
rect 16112 2144 16120 2208
rect 15800 2128 16120 2144
rect 19514 28864 19834 29424
rect 19514 28800 19522 28864
rect 19586 28800 19602 28864
rect 19666 28800 19682 28864
rect 19746 28800 19762 28864
rect 19826 28800 19834 28864
rect 19514 27776 19834 28800
rect 19514 27712 19522 27776
rect 19586 27712 19602 27776
rect 19666 27712 19682 27776
rect 19746 27712 19762 27776
rect 19826 27712 19834 27776
rect 19514 26688 19834 27712
rect 19514 26624 19522 26688
rect 19586 26624 19602 26688
rect 19666 26624 19682 26688
rect 19746 26624 19762 26688
rect 19826 26624 19834 26688
rect 19514 25600 19834 26624
rect 19514 25536 19522 25600
rect 19586 25536 19602 25600
rect 19666 25536 19682 25600
rect 19746 25536 19762 25600
rect 19826 25536 19834 25600
rect 19514 24512 19834 25536
rect 19514 24448 19522 24512
rect 19586 24448 19602 24512
rect 19666 24448 19682 24512
rect 19746 24448 19762 24512
rect 19826 24448 19834 24512
rect 19514 23424 19834 24448
rect 19514 23360 19522 23424
rect 19586 23360 19602 23424
rect 19666 23360 19682 23424
rect 19746 23360 19762 23424
rect 19826 23360 19834 23424
rect 19514 22336 19834 23360
rect 19514 22272 19522 22336
rect 19586 22272 19602 22336
rect 19666 22272 19682 22336
rect 19746 22272 19762 22336
rect 19826 22272 19834 22336
rect 19514 21248 19834 22272
rect 19514 21184 19522 21248
rect 19586 21184 19602 21248
rect 19666 21184 19682 21248
rect 19746 21184 19762 21248
rect 19826 21184 19834 21248
rect 19514 20160 19834 21184
rect 19514 20096 19522 20160
rect 19586 20096 19602 20160
rect 19666 20096 19682 20160
rect 19746 20096 19762 20160
rect 19826 20096 19834 20160
rect 19514 19072 19834 20096
rect 19514 19008 19522 19072
rect 19586 19008 19602 19072
rect 19666 19008 19682 19072
rect 19746 19008 19762 19072
rect 19826 19008 19834 19072
rect 19514 17984 19834 19008
rect 19514 17920 19522 17984
rect 19586 17920 19602 17984
rect 19666 17920 19682 17984
rect 19746 17920 19762 17984
rect 19826 17920 19834 17984
rect 19514 16896 19834 17920
rect 19514 16832 19522 16896
rect 19586 16832 19602 16896
rect 19666 16832 19682 16896
rect 19746 16832 19762 16896
rect 19826 16832 19834 16896
rect 19514 15808 19834 16832
rect 19514 15744 19522 15808
rect 19586 15744 19602 15808
rect 19666 15744 19682 15808
rect 19746 15744 19762 15808
rect 19826 15744 19834 15808
rect 19514 14720 19834 15744
rect 19514 14656 19522 14720
rect 19586 14656 19602 14720
rect 19666 14656 19682 14720
rect 19746 14656 19762 14720
rect 19826 14656 19834 14720
rect 19514 13632 19834 14656
rect 19514 13568 19522 13632
rect 19586 13568 19602 13632
rect 19666 13568 19682 13632
rect 19746 13568 19762 13632
rect 19826 13568 19834 13632
rect 19514 12544 19834 13568
rect 19514 12480 19522 12544
rect 19586 12480 19602 12544
rect 19666 12480 19682 12544
rect 19746 12480 19762 12544
rect 19826 12480 19834 12544
rect 19514 11456 19834 12480
rect 19514 11392 19522 11456
rect 19586 11392 19602 11456
rect 19666 11392 19682 11456
rect 19746 11392 19762 11456
rect 19826 11392 19834 11456
rect 19514 10368 19834 11392
rect 19514 10304 19522 10368
rect 19586 10304 19602 10368
rect 19666 10304 19682 10368
rect 19746 10304 19762 10368
rect 19826 10304 19834 10368
rect 19514 9280 19834 10304
rect 19514 9216 19522 9280
rect 19586 9216 19602 9280
rect 19666 9216 19682 9280
rect 19746 9216 19762 9280
rect 19826 9216 19834 9280
rect 19514 8192 19834 9216
rect 19514 8128 19522 8192
rect 19586 8128 19602 8192
rect 19666 8128 19682 8192
rect 19746 8128 19762 8192
rect 19826 8128 19834 8192
rect 19514 7104 19834 8128
rect 19514 7040 19522 7104
rect 19586 7040 19602 7104
rect 19666 7040 19682 7104
rect 19746 7040 19762 7104
rect 19826 7040 19834 7104
rect 19514 6016 19834 7040
rect 19514 5952 19522 6016
rect 19586 5952 19602 6016
rect 19666 5952 19682 6016
rect 19746 5952 19762 6016
rect 19826 5952 19834 6016
rect 19514 4928 19834 5952
rect 19514 4864 19522 4928
rect 19586 4864 19602 4928
rect 19666 4864 19682 4928
rect 19746 4864 19762 4928
rect 19826 4864 19834 4928
rect 19514 3840 19834 4864
rect 19514 3776 19522 3840
rect 19586 3776 19602 3840
rect 19666 3776 19682 3840
rect 19746 3776 19762 3840
rect 19826 3776 19834 3840
rect 19514 2752 19834 3776
rect 19514 2688 19522 2752
rect 19586 2688 19602 2752
rect 19666 2688 19682 2752
rect 19746 2688 19762 2752
rect 19826 2688 19834 2752
rect 19514 2128 19834 2688
rect 23228 29408 23548 29424
rect 23228 29344 23236 29408
rect 23300 29344 23316 29408
rect 23380 29344 23396 29408
rect 23460 29344 23476 29408
rect 23540 29344 23548 29408
rect 23228 28320 23548 29344
rect 23228 28256 23236 28320
rect 23300 28256 23316 28320
rect 23380 28256 23396 28320
rect 23460 28256 23476 28320
rect 23540 28256 23548 28320
rect 23228 27232 23548 28256
rect 23228 27168 23236 27232
rect 23300 27168 23316 27232
rect 23380 27168 23396 27232
rect 23460 27168 23476 27232
rect 23540 27168 23548 27232
rect 23228 26144 23548 27168
rect 23228 26080 23236 26144
rect 23300 26080 23316 26144
rect 23380 26080 23396 26144
rect 23460 26080 23476 26144
rect 23540 26080 23548 26144
rect 23228 25056 23548 26080
rect 23228 24992 23236 25056
rect 23300 24992 23316 25056
rect 23380 24992 23396 25056
rect 23460 24992 23476 25056
rect 23540 24992 23548 25056
rect 23228 23968 23548 24992
rect 23228 23904 23236 23968
rect 23300 23904 23316 23968
rect 23380 23904 23396 23968
rect 23460 23904 23476 23968
rect 23540 23904 23548 23968
rect 23228 22880 23548 23904
rect 23228 22816 23236 22880
rect 23300 22816 23316 22880
rect 23380 22816 23396 22880
rect 23460 22816 23476 22880
rect 23540 22816 23548 22880
rect 23228 21792 23548 22816
rect 23228 21728 23236 21792
rect 23300 21728 23316 21792
rect 23380 21728 23396 21792
rect 23460 21728 23476 21792
rect 23540 21728 23548 21792
rect 23228 20704 23548 21728
rect 23228 20640 23236 20704
rect 23300 20640 23316 20704
rect 23380 20640 23396 20704
rect 23460 20640 23476 20704
rect 23540 20640 23548 20704
rect 23228 19616 23548 20640
rect 23228 19552 23236 19616
rect 23300 19552 23316 19616
rect 23380 19552 23396 19616
rect 23460 19552 23476 19616
rect 23540 19552 23548 19616
rect 23228 18528 23548 19552
rect 23228 18464 23236 18528
rect 23300 18464 23316 18528
rect 23380 18464 23396 18528
rect 23460 18464 23476 18528
rect 23540 18464 23548 18528
rect 23228 17440 23548 18464
rect 23228 17376 23236 17440
rect 23300 17376 23316 17440
rect 23380 17376 23396 17440
rect 23460 17376 23476 17440
rect 23540 17376 23548 17440
rect 23228 16352 23548 17376
rect 23228 16288 23236 16352
rect 23300 16288 23316 16352
rect 23380 16288 23396 16352
rect 23460 16288 23476 16352
rect 23540 16288 23548 16352
rect 23228 15264 23548 16288
rect 23228 15200 23236 15264
rect 23300 15200 23316 15264
rect 23380 15200 23396 15264
rect 23460 15200 23476 15264
rect 23540 15200 23548 15264
rect 23228 14176 23548 15200
rect 23228 14112 23236 14176
rect 23300 14112 23316 14176
rect 23380 14112 23396 14176
rect 23460 14112 23476 14176
rect 23540 14112 23548 14176
rect 23228 13088 23548 14112
rect 23228 13024 23236 13088
rect 23300 13024 23316 13088
rect 23380 13024 23396 13088
rect 23460 13024 23476 13088
rect 23540 13024 23548 13088
rect 23228 12000 23548 13024
rect 23228 11936 23236 12000
rect 23300 11936 23316 12000
rect 23380 11936 23396 12000
rect 23460 11936 23476 12000
rect 23540 11936 23548 12000
rect 23228 10912 23548 11936
rect 23228 10848 23236 10912
rect 23300 10848 23316 10912
rect 23380 10848 23396 10912
rect 23460 10848 23476 10912
rect 23540 10848 23548 10912
rect 23228 9824 23548 10848
rect 23228 9760 23236 9824
rect 23300 9760 23316 9824
rect 23380 9760 23396 9824
rect 23460 9760 23476 9824
rect 23540 9760 23548 9824
rect 23228 8736 23548 9760
rect 23228 8672 23236 8736
rect 23300 8672 23316 8736
rect 23380 8672 23396 8736
rect 23460 8672 23476 8736
rect 23540 8672 23548 8736
rect 23228 7648 23548 8672
rect 23228 7584 23236 7648
rect 23300 7584 23316 7648
rect 23380 7584 23396 7648
rect 23460 7584 23476 7648
rect 23540 7584 23548 7648
rect 23228 6560 23548 7584
rect 23228 6496 23236 6560
rect 23300 6496 23316 6560
rect 23380 6496 23396 6560
rect 23460 6496 23476 6560
rect 23540 6496 23548 6560
rect 23228 5472 23548 6496
rect 23228 5408 23236 5472
rect 23300 5408 23316 5472
rect 23380 5408 23396 5472
rect 23460 5408 23476 5472
rect 23540 5408 23548 5472
rect 23228 4384 23548 5408
rect 23228 4320 23236 4384
rect 23300 4320 23316 4384
rect 23380 4320 23396 4384
rect 23460 4320 23476 4384
rect 23540 4320 23548 4384
rect 23228 3296 23548 4320
rect 23228 3232 23236 3296
rect 23300 3232 23316 3296
rect 23380 3232 23396 3296
rect 23460 3232 23476 3296
rect 23540 3232 23548 3296
rect 23228 2208 23548 3232
rect 23228 2144 23236 2208
rect 23300 2144 23316 2208
rect 23380 2144 23396 2208
rect 23460 2144 23476 2208
rect 23540 2144 23548 2208
rect 23228 2128 23548 2144
rect 26942 28864 27262 29424
rect 26942 28800 26950 28864
rect 27014 28800 27030 28864
rect 27094 28800 27110 28864
rect 27174 28800 27190 28864
rect 27254 28800 27262 28864
rect 26942 27776 27262 28800
rect 26942 27712 26950 27776
rect 27014 27712 27030 27776
rect 27094 27712 27110 27776
rect 27174 27712 27190 27776
rect 27254 27712 27262 27776
rect 26942 26688 27262 27712
rect 26942 26624 26950 26688
rect 27014 26624 27030 26688
rect 27094 26624 27110 26688
rect 27174 26624 27190 26688
rect 27254 26624 27262 26688
rect 26942 25600 27262 26624
rect 26942 25536 26950 25600
rect 27014 25536 27030 25600
rect 27094 25536 27110 25600
rect 27174 25536 27190 25600
rect 27254 25536 27262 25600
rect 26942 24512 27262 25536
rect 26942 24448 26950 24512
rect 27014 24448 27030 24512
rect 27094 24448 27110 24512
rect 27174 24448 27190 24512
rect 27254 24448 27262 24512
rect 26942 23424 27262 24448
rect 26942 23360 26950 23424
rect 27014 23360 27030 23424
rect 27094 23360 27110 23424
rect 27174 23360 27190 23424
rect 27254 23360 27262 23424
rect 26942 22336 27262 23360
rect 26942 22272 26950 22336
rect 27014 22272 27030 22336
rect 27094 22272 27110 22336
rect 27174 22272 27190 22336
rect 27254 22272 27262 22336
rect 26942 21248 27262 22272
rect 26942 21184 26950 21248
rect 27014 21184 27030 21248
rect 27094 21184 27110 21248
rect 27174 21184 27190 21248
rect 27254 21184 27262 21248
rect 26942 20160 27262 21184
rect 26942 20096 26950 20160
rect 27014 20096 27030 20160
rect 27094 20096 27110 20160
rect 27174 20096 27190 20160
rect 27254 20096 27262 20160
rect 26942 19072 27262 20096
rect 26942 19008 26950 19072
rect 27014 19008 27030 19072
rect 27094 19008 27110 19072
rect 27174 19008 27190 19072
rect 27254 19008 27262 19072
rect 26942 17984 27262 19008
rect 26942 17920 26950 17984
rect 27014 17920 27030 17984
rect 27094 17920 27110 17984
rect 27174 17920 27190 17984
rect 27254 17920 27262 17984
rect 26942 16896 27262 17920
rect 26942 16832 26950 16896
rect 27014 16832 27030 16896
rect 27094 16832 27110 16896
rect 27174 16832 27190 16896
rect 27254 16832 27262 16896
rect 26942 15808 27262 16832
rect 26942 15744 26950 15808
rect 27014 15744 27030 15808
rect 27094 15744 27110 15808
rect 27174 15744 27190 15808
rect 27254 15744 27262 15808
rect 26942 14720 27262 15744
rect 26942 14656 26950 14720
rect 27014 14656 27030 14720
rect 27094 14656 27110 14720
rect 27174 14656 27190 14720
rect 27254 14656 27262 14720
rect 26942 13632 27262 14656
rect 26942 13568 26950 13632
rect 27014 13568 27030 13632
rect 27094 13568 27110 13632
rect 27174 13568 27190 13632
rect 27254 13568 27262 13632
rect 26942 12544 27262 13568
rect 26942 12480 26950 12544
rect 27014 12480 27030 12544
rect 27094 12480 27110 12544
rect 27174 12480 27190 12544
rect 27254 12480 27262 12544
rect 26942 11456 27262 12480
rect 26942 11392 26950 11456
rect 27014 11392 27030 11456
rect 27094 11392 27110 11456
rect 27174 11392 27190 11456
rect 27254 11392 27262 11456
rect 26942 10368 27262 11392
rect 26942 10304 26950 10368
rect 27014 10304 27030 10368
rect 27094 10304 27110 10368
rect 27174 10304 27190 10368
rect 27254 10304 27262 10368
rect 26942 9280 27262 10304
rect 26942 9216 26950 9280
rect 27014 9216 27030 9280
rect 27094 9216 27110 9280
rect 27174 9216 27190 9280
rect 27254 9216 27262 9280
rect 26942 8192 27262 9216
rect 26942 8128 26950 8192
rect 27014 8128 27030 8192
rect 27094 8128 27110 8192
rect 27174 8128 27190 8192
rect 27254 8128 27262 8192
rect 26942 7104 27262 8128
rect 26942 7040 26950 7104
rect 27014 7040 27030 7104
rect 27094 7040 27110 7104
rect 27174 7040 27190 7104
rect 27254 7040 27262 7104
rect 26942 6016 27262 7040
rect 26942 5952 26950 6016
rect 27014 5952 27030 6016
rect 27094 5952 27110 6016
rect 27174 5952 27190 6016
rect 27254 5952 27262 6016
rect 26942 4928 27262 5952
rect 26942 4864 26950 4928
rect 27014 4864 27030 4928
rect 27094 4864 27110 4928
rect 27174 4864 27190 4928
rect 27254 4864 27262 4928
rect 26942 3840 27262 4864
rect 26942 3776 26950 3840
rect 27014 3776 27030 3840
rect 27094 3776 27110 3840
rect 27174 3776 27190 3840
rect 27254 3776 27262 3840
rect 26942 2752 27262 3776
rect 26942 2688 26950 2752
rect 27014 2688 27030 2752
rect 27094 2688 27110 2752
rect 27174 2688 27190 2752
rect 27254 2688 27262 2752
rect 26942 2128 27262 2688
rect 30656 29408 30976 29424
rect 30656 29344 30664 29408
rect 30728 29344 30744 29408
rect 30808 29344 30824 29408
rect 30888 29344 30904 29408
rect 30968 29344 30976 29408
rect 30656 28320 30976 29344
rect 30656 28256 30664 28320
rect 30728 28256 30744 28320
rect 30808 28256 30824 28320
rect 30888 28256 30904 28320
rect 30968 28256 30976 28320
rect 30656 27232 30976 28256
rect 30656 27168 30664 27232
rect 30728 27168 30744 27232
rect 30808 27168 30824 27232
rect 30888 27168 30904 27232
rect 30968 27168 30976 27232
rect 30656 26144 30976 27168
rect 30656 26080 30664 26144
rect 30728 26080 30744 26144
rect 30808 26080 30824 26144
rect 30888 26080 30904 26144
rect 30968 26080 30976 26144
rect 30656 25056 30976 26080
rect 30656 24992 30664 25056
rect 30728 24992 30744 25056
rect 30808 24992 30824 25056
rect 30888 24992 30904 25056
rect 30968 24992 30976 25056
rect 30656 23968 30976 24992
rect 30656 23904 30664 23968
rect 30728 23904 30744 23968
rect 30808 23904 30824 23968
rect 30888 23904 30904 23968
rect 30968 23904 30976 23968
rect 30656 22880 30976 23904
rect 30656 22816 30664 22880
rect 30728 22816 30744 22880
rect 30808 22816 30824 22880
rect 30888 22816 30904 22880
rect 30968 22816 30976 22880
rect 30656 21792 30976 22816
rect 30656 21728 30664 21792
rect 30728 21728 30744 21792
rect 30808 21728 30824 21792
rect 30888 21728 30904 21792
rect 30968 21728 30976 21792
rect 30656 20704 30976 21728
rect 30656 20640 30664 20704
rect 30728 20640 30744 20704
rect 30808 20640 30824 20704
rect 30888 20640 30904 20704
rect 30968 20640 30976 20704
rect 30656 19616 30976 20640
rect 30656 19552 30664 19616
rect 30728 19552 30744 19616
rect 30808 19552 30824 19616
rect 30888 19552 30904 19616
rect 30968 19552 30976 19616
rect 30656 18528 30976 19552
rect 30656 18464 30664 18528
rect 30728 18464 30744 18528
rect 30808 18464 30824 18528
rect 30888 18464 30904 18528
rect 30968 18464 30976 18528
rect 30656 17440 30976 18464
rect 30656 17376 30664 17440
rect 30728 17376 30744 17440
rect 30808 17376 30824 17440
rect 30888 17376 30904 17440
rect 30968 17376 30976 17440
rect 30656 16352 30976 17376
rect 30656 16288 30664 16352
rect 30728 16288 30744 16352
rect 30808 16288 30824 16352
rect 30888 16288 30904 16352
rect 30968 16288 30976 16352
rect 30656 15264 30976 16288
rect 30656 15200 30664 15264
rect 30728 15200 30744 15264
rect 30808 15200 30824 15264
rect 30888 15200 30904 15264
rect 30968 15200 30976 15264
rect 30656 14176 30976 15200
rect 30656 14112 30664 14176
rect 30728 14112 30744 14176
rect 30808 14112 30824 14176
rect 30888 14112 30904 14176
rect 30968 14112 30976 14176
rect 30656 13088 30976 14112
rect 30656 13024 30664 13088
rect 30728 13024 30744 13088
rect 30808 13024 30824 13088
rect 30888 13024 30904 13088
rect 30968 13024 30976 13088
rect 30656 12000 30976 13024
rect 30656 11936 30664 12000
rect 30728 11936 30744 12000
rect 30808 11936 30824 12000
rect 30888 11936 30904 12000
rect 30968 11936 30976 12000
rect 30656 10912 30976 11936
rect 30656 10848 30664 10912
rect 30728 10848 30744 10912
rect 30808 10848 30824 10912
rect 30888 10848 30904 10912
rect 30968 10848 30976 10912
rect 30656 9824 30976 10848
rect 30656 9760 30664 9824
rect 30728 9760 30744 9824
rect 30808 9760 30824 9824
rect 30888 9760 30904 9824
rect 30968 9760 30976 9824
rect 30656 8736 30976 9760
rect 30656 8672 30664 8736
rect 30728 8672 30744 8736
rect 30808 8672 30824 8736
rect 30888 8672 30904 8736
rect 30968 8672 30976 8736
rect 30656 7648 30976 8672
rect 30656 7584 30664 7648
rect 30728 7584 30744 7648
rect 30808 7584 30824 7648
rect 30888 7584 30904 7648
rect 30968 7584 30976 7648
rect 30656 6560 30976 7584
rect 30656 6496 30664 6560
rect 30728 6496 30744 6560
rect 30808 6496 30824 6560
rect 30888 6496 30904 6560
rect 30968 6496 30976 6560
rect 30656 5472 30976 6496
rect 30656 5408 30664 5472
rect 30728 5408 30744 5472
rect 30808 5408 30824 5472
rect 30888 5408 30904 5472
rect 30968 5408 30976 5472
rect 30656 4384 30976 5408
rect 30656 4320 30664 4384
rect 30728 4320 30744 4384
rect 30808 4320 30824 4384
rect 30888 4320 30904 4384
rect 30968 4320 30976 4384
rect 30656 3296 30976 4320
rect 30656 3232 30664 3296
rect 30728 3232 30744 3296
rect 30808 3232 30824 3296
rect 30888 3232 30904 3296
rect 30968 3232 30976 3296
rect 30656 2208 30976 3232
rect 30656 2144 30664 2208
rect 30728 2144 30744 2208
rect 30808 2144 30824 2208
rect 30888 2144 30904 2208
rect 30968 2144 30976 2208
rect 30656 2128 30976 2144
use sky130_ef_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1676037725
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1676037725
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1676037725
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1676037725
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1676037725
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1676037725
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1676037725
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1676037725
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1676037725
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1676037725
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1676037725
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1676037725
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1676037725
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1676037725
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1676037725
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1676037725
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1676037725
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1676037725
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1676037725
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1676037725
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_309
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_318 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 30360 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1676037725
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1676037725
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1676037725
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1676037725
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1676037725
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1676037725
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1676037725
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1676037725
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1676037725
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1676037725
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1676037725
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1676037725
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1676037725
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1676037725
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1676037725
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1676037725
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1676037725
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_317
timestamp 1676037725
transform 1 0 30268 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1676037725
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1676037725
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1676037725
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1676037725
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1676037725
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1676037725
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1676037725
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1676037725
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1676037725
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1676037725
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_309 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_317
timestamp 1676037725
transform 1 0 30268 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_153
timestamp 1676037725
transform 1 0 15180 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_165
timestamp 1676037725
transform 1 0 16284 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1676037725
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1676037725
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1676037725
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1676037725
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1676037725
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1676037725
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1676037725
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_317
timestamp 1676037725
transform 1 0 30268 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_151
timestamp 1676037725
transform 1 0 14996 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_171
timestamp 1676037725
transform 1 0 16836 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_182
timestamp 1676037725
transform 1 0 17848 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1676037725
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_215
timestamp 1676037725
transform 1 0 20884 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_227
timestamp 1676037725
transform 1 0 21988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_239
timestamp 1676037725
transform 1 0 23092 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1676037725
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1676037725
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1676037725
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1676037725
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1676037725
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_317
timestamp 1676037725
transform 1 0 30268 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_145
timestamp 1676037725
transform 1 0 14444 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_157
timestamp 1676037725
transform 1 0 15548 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_165
timestamp 1676037725
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_188
timestamp 1676037725
transform 1 0 18400 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_208
timestamp 1676037725
transform 1 0 20240 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_220
timestamp 1676037725
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1676037725
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1676037725
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1676037725
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1676037725
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1676037725
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_285
timestamp 1676037725
transform 1 0 27324 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_291
timestamp 1676037725
transform 1 0 27876 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_299
timestamp 1676037725
transform 1 0 28612 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_303
timestamp 1676037725
transform 1 0 28980 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_315
timestamp 1676037725
transform 1 0 30084 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_319
timestamp 1676037725
transform 1 0 30452 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_105
timestamp 1676037725
transform 1 0 10764 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_159
timestamp 1676037725
transform 1 0 15732 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_171
timestamp 1676037725
transform 1 0 16836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_183
timestamp 1676037725
transform 1 0 17940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_206
timestamp 1676037725
transform 1 0 20056 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_218
timestamp 1676037725
transform 1 0 21160 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_242
timestamp 1676037725
transform 1 0 23368 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1676037725
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_271
timestamp 1676037725
transform 1 0 26036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_277
timestamp 1676037725
transform 1 0 26588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_288
timestamp 1676037725
transform 1 0 27600 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_299
timestamp 1676037725
transform 1 0 28612 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp 1676037725
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_318
timestamp 1676037725
transform 1 0 30360 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1676037725
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_62
timestamp 1676037725
transform 1 0 6808 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_74
timestamp 1676037725
transform 1 0 7912 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_98
timestamp 1676037725
transform 1 0 10120 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_106
timestamp 1676037725
transform 1 0 10856 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1676037725
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_136
timestamp 1676037725
transform 1 0 13616 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_148
timestamp 1676037725
transform 1 0 14720 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_160
timestamp 1676037725
transform 1 0 15824 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1676037725
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1676037725
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1676037725
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_248
timestamp 1676037725
transform 1 0 23920 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_268
timestamp 1676037725
transform 1 0 25760 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_274
timestamp 1676037725
transform 1 0 26312 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp 1676037725
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_300
timestamp 1676037725
transform 1 0 28704 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_311
timestamp 1676037725
transform 1 0 29716 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_318
timestamp 1676037725
transform 1 0 30360 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_45
timestamp 1676037725
transform 1 0 5244 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_67
timestamp 1676037725
transform 1 0 7268 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1676037725
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_108
timestamp 1676037725
transform 1 0 11040 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_120
timestamp 1676037725
transform 1 0 12144 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_132
timestamp 1676037725
transform 1 0 13248 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_164
timestamp 1676037725
transform 1 0 16192 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_174
timestamp 1676037725
transform 1 0 17112 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_181
timestamp 1676037725
transform 1 0 17756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_193
timestamp 1676037725
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_209
timestamp 1676037725
transform 1 0 20332 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_231
timestamp 1676037725
transform 1 0 22356 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_243
timestamp 1676037725
transform 1 0 23460 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1676037725
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_272
timestamp 1676037725
transform 1 0 26128 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_288
timestamp 1676037725
transform 1 0 27600 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_296
timestamp 1676037725
transform 1 0 28336 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_305
timestamp 1676037725
transform 1 0 29164 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_317
timestamp 1676037725
transform 1 0 30268 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_39
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1676037725
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_62
timestamp 1676037725
transform 1 0 6808 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_70
timestamp 1676037725
transform 1 0 7544 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_101
timestamp 1676037725
transform 1 0 10396 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_107
timestamp 1676037725
transform 1 0 10948 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_128
timestamp 1676037725
transform 1 0 12880 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_140
timestamp 1676037725
transform 1 0 13984 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_152
timestamp 1676037725
transform 1 0 15088 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_160
timestamp 1676037725
transform 1 0 15824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1676037725
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_191
timestamp 1676037725
transform 1 0 18676 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_203
timestamp 1676037725
transform 1 0 19780 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_215
timestamp 1676037725
transform 1 0 20884 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1676037725
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_230
timestamp 1676037725
transform 1 0 22264 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1676037725
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1676037725
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_261
timestamp 1676037725
transform 1 0 25116 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_265
timestamp 1676037725
transform 1 0 25484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_277
timestamp 1676037725
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_285
timestamp 1676037725
transform 1 0 27324 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_289
timestamp 1676037725
transform 1 0 27692 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_310
timestamp 1676037725
transform 1 0 29624 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_318
timestamp 1676037725
transform 1 0 30360 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_45
timestamp 1676037725
transform 1 0 5244 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_67
timestamp 1676037725
transform 1 0 7268 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_74
timestamp 1676037725
transform 1 0 7912 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1676037725
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_90
timestamp 1676037725
transform 1 0 9384 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_102
timestamp 1676037725
transform 1 0 10488 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_126
timestamp 1676037725
transform 1 0 12696 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_135
timestamp 1676037725
transform 1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_153
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_159
timestamp 1676037725
transform 1 0 15732 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_166
timestamp 1676037725
transform 1 0 16376 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_191
timestamp 1676037725
transform 1 0 18676 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1676037725
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_202
timestamp 1676037725
transform 1 0 19688 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_210
timestamp 1676037725
transform 1 0 20424 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_231
timestamp 1676037725
transform 1 0 22356 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_243
timestamp 1676037725
transform 1 0 23460 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1676037725
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_271
timestamp 1676037725
transform 1 0 26036 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_283
timestamp 1676037725
transform 1 0 27140 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_295
timestamp 1676037725
transform 1 0 28244 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_299
timestamp 1676037725
transform 1 0 28612 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1676037725
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_317
timestamp 1676037725
transform 1 0 30268 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_47
timestamp 1676037725
transform 1 0 5428 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1676037725
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_62
timestamp 1676037725
transform 1 0 6808 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_70
timestamp 1676037725
transform 1 0 7544 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1676037725
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_124
timestamp 1676037725
transform 1 0 12512 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_135
timestamp 1676037725
transform 1 0 13524 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_142
timestamp 1676037725
transform 1 0 14168 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_154
timestamp 1676037725
transform 1 0 15272 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1676037725
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_191
timestamp 1676037725
transform 1 0 18676 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_216
timestamp 1676037725
transform 1 0 20976 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_230
timestamp 1676037725
transform 1 0 22264 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_242
timestamp 1676037725
transform 1 0 23368 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_246
timestamp 1676037725
transform 1 0 23736 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_263
timestamp 1676037725
transform 1 0 25300 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_275
timestamp 1676037725
transform 1 0 26404 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1676037725
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_287
timestamp 1676037725
transform 1 0 27508 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_294
timestamp 1676037725
transform 1 0 28152 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_301
timestamp 1676037725
transform 1 0 28796 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_313
timestamp 1676037725
transform 1 0 29900 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_319
timestamp 1676037725
transform 1 0 30452 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1676037725
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_94
timestamp 1676037725
transform 1 0 9752 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_106
timestamp 1676037725
transform 1 0 10856 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_118
timestamp 1676037725
transform 1 0 11960 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_126
timestamp 1676037725
transform 1 0 12696 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_134
timestamp 1676037725
transform 1 0 13432 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_161
timestamp 1676037725
transform 1 0 15916 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_173
timestamp 1676037725
transform 1 0 17020 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_185
timestamp 1676037725
transform 1 0 18124 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_193
timestamp 1676037725
transform 1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_203
timestamp 1676037725
transform 1 0 19780 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_207
timestamp 1676037725
transform 1 0 20148 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_219
timestamp 1676037725
transform 1 0 21252 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_231
timestamp 1676037725
transform 1 0 22356 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_238
timestamp 1676037725
transform 1 0 23000 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1676037725
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_258
timestamp 1676037725
transform 1 0 24840 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_270
timestamp 1676037725
transform 1 0 25944 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_282
timestamp 1676037725
transform 1 0 27048 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_288
timestamp 1676037725
transform 1 0 27600 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_296
timestamp 1676037725
transform 1 0 28336 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_305
timestamp 1676037725
transform 1 0 29164 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_318
timestamp 1676037725
transform 1 0 30360 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_53
timestamp 1676037725
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_63
timestamp 1676037725
transform 1 0 6900 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_80
timestamp 1676037725
transform 1 0 8464 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_92
timestamp 1676037725
transform 1 0 9568 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1676037725
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_124
timestamp 1676037725
transform 1 0 12512 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_136
timestamp 1676037725
transform 1 0 13616 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_148
timestamp 1676037725
transform 1 0 14720 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_158
timestamp 1676037725
transform 1 0 15640 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1676037725
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_184
timestamp 1676037725
transform 1 0 18032 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_196
timestamp 1676037725
transform 1 0 19136 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_208
timestamp 1676037725
transform 1 0 20240 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 1676037725
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_243
timestamp 1676037725
transform 1 0 23460 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_251
timestamp 1676037725
transform 1 0 24196 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1676037725
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1676037725
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_289
timestamp 1676037725
transform 1 0 27692 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_308
timestamp 1676037725
transform 1 0 29440 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_318
timestamp 1676037725
transform 1 0 30360 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 1676037725
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_93
timestamp 1676037725
transform 1 0 9660 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_115
timestamp 1676037725
transform 1 0 11684 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_123
timestamp 1676037725
transform 1 0 12420 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_131
timestamp 1676037725
transform 1 0 13156 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1676037725
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_152
timestamp 1676037725
transform 1 0 15088 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_164
timestamp 1676037725
transform 1 0 16192 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_170
timestamp 1676037725
transform 1 0 16744 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_184
timestamp 1676037725
transform 1 0 18032 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_209
timestamp 1676037725
transform 1 0 20332 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1676037725
transform 1 0 20700 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_234
timestamp 1676037725
transform 1 0 22632 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_246
timestamp 1676037725
transform 1 0 23736 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_268
timestamp 1676037725
transform 1 0 25760 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_280
timestamp 1676037725
transform 1 0 26864 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_288
timestamp 1676037725
transform 1 0 27600 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_298
timestamp 1676037725
transform 1 0 28520 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_305
timestamp 1676037725
transform 1 0 29164 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1676037725
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_317
timestamp 1676037725
transform 1 0 30268 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1676037725
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_27
timestamp 1676037725
transform 1 0 3588 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1676037725
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_62
timestamp 1676037725
transform 1 0 6808 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_75
timestamp 1676037725
transform 1 0 8004 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_103
timestamp 1676037725
transform 1 0 10580 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1676037725
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_119
timestamp 1676037725
transform 1 0 12052 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_127
timestamp 1676037725
transform 1 0 12788 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_147
timestamp 1676037725
transform 1 0 14628 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_159
timestamp 1676037725
transform 1 0 15732 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1676037725
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_192
timestamp 1676037725
transform 1 0 18768 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_196
timestamp 1676037725
transform 1 0 19136 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_210
timestamp 1676037725
transform 1 0 20424 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1676037725
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_240
timestamp 1676037725
transform 1 0 23184 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_252
timestamp 1676037725
transform 1 0 24288 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_256
timestamp 1676037725
transform 1 0 24656 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_278
timestamp 1676037725
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_294
timestamp 1676037725
transform 1 0 28152 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_306
timestamp 1676037725
transform 1 0 29256 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_313
timestamp 1676037725
transform 1 0 29900 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_319
timestamp 1676037725
transform 1 0 30452 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_35
timestamp 1676037725
transform 1 0 4324 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_52
timestamp 1676037725
transform 1 0 5888 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_64
timestamp 1676037725
transform 1 0 6992 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_79
timestamp 1676037725
transform 1 0 8372 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_93
timestamp 1676037725
transform 1 0 9660 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_98
timestamp 1676037725
transform 1 0 10120 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_110
timestamp 1676037725
transform 1 0 11224 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_118
timestamp 1676037725
transform 1 0 11960 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_135
timestamp 1676037725
transform 1 0 13524 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1676037725
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_153
timestamp 1676037725
transform 1 0 15180 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_161
timestamp 1676037725
transform 1 0 15916 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_165
timestamp 1676037725
transform 1 0 16284 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_190
timestamp 1676037725
transform 1 0 18584 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_220
timestamp 1676037725
transform 1 0 21344 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1676037725
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1676037725
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_259
timestamp 1676037725
transform 1 0 24932 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_272
timestamp 1676037725
transform 1 0 26128 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_284
timestamp 1676037725
transform 1 0 27232 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_296
timestamp 1676037725
transform 1 0 28336 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_306
timestamp 1676037725
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1676037725
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_318
timestamp 1676037725
transform 1 0 30360 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_27
timestamp 1676037725
transform 1 0 3588 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1676037725
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_61
timestamp 1676037725
transform 1 0 6716 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_78
timestamp 1676037725
transform 1 0 8280 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_85
timestamp 1676037725
transform 1 0 8924 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_89
timestamp 1676037725
transform 1 0 9292 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_97
timestamp 1676037725
transform 1 0 10028 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_107
timestamp 1676037725
transform 1 0 10948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_134
timestamp 1676037725
transform 1 0 13432 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_146
timestamp 1676037725
transform 1 0 14536 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_158
timestamp 1676037725
transform 1 0 15640 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1676037725
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_173
timestamp 1676037725
transform 1 0 17020 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_190
timestamp 1676037725
transform 1 0 18584 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_197
timestamp 1676037725
transform 1 0 19228 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_201
timestamp 1676037725
transform 1 0 19596 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_205
timestamp 1676037725
transform 1 0 19964 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_216
timestamp 1676037725
transform 1 0 20976 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_230
timestamp 1676037725
transform 1 0 22264 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1676037725
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1676037725
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1676037725
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1676037725
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1676037725
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1676037725
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_317
timestamp 1676037725
transform 1 0 30268 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_37
timestamp 1676037725
transform 1 0 4508 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_43
timestamp 1676037725
transform 1 0 5060 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_50
timestamp 1676037725
transform 1 0 5704 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_62
timestamp 1676037725
transform 1 0 6808 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_66
timestamp 1676037725
transform 1 0 7176 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_78
timestamp 1676037725
transform 1 0 8280 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1676037725
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_121
timestamp 1676037725
transform 1 0 12236 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_125
timestamp 1676037725
transform 1 0 12604 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_137
timestamp 1676037725
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_153
timestamp 1676037725
transform 1 0 15180 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_159
timestamp 1676037725
transform 1 0 15732 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_176
timestamp 1676037725
transform 1 0 17296 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_183
timestamp 1676037725
transform 1 0 17940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1676037725
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1676037725
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_221
timestamp 1676037725
transform 1 0 21436 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1676037725
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_259
timestamp 1676037725
transform 1 0 24932 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_273
timestamp 1676037725
transform 1 0 26220 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_285
timestamp 1676037725
transform 1 0 27324 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_297
timestamp 1676037725
transform 1 0 28428 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_305
timestamp 1676037725
transform 1 0 29164 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_309
timestamp 1676037725
transform 1 0 29532 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_317
timestamp 1676037725
transform 1 0 30268 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_52
timestamp 1676037725
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_65
timestamp 1676037725
transform 1 0 7084 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_72
timestamp 1676037725
transform 1 0 7728 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_76
timestamp 1676037725
transform 1 0 8096 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_84
timestamp 1676037725
transform 1 0 8832 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_97
timestamp 1676037725
transform 1 0 10028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_109
timestamp 1676037725
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_125
timestamp 1676037725
transform 1 0 12604 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_144
timestamp 1676037725
transform 1 0 14352 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_157
timestamp 1676037725
transform 1 0 15548 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_165
timestamp 1676037725
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_180
timestamp 1676037725
transform 1 0 17664 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_192
timestamp 1676037725
transform 1 0 18768 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_198
timestamp 1676037725
transform 1 0 19320 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_206
timestamp 1676037725
transform 1 0 20056 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_218
timestamp 1676037725
transform 1 0 21160 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_233
timestamp 1676037725
transform 1 0 22540 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_238
timestamp 1676037725
transform 1 0 23000 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_245
timestamp 1676037725
transform 1 0 23644 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_249
timestamp 1676037725
transform 1 0 24012 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_253
timestamp 1676037725
transform 1 0 24380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1676037725
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_298
timestamp 1676037725
transform 1 0 28520 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_315
timestamp 1676037725
transform 1 0 30084 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_319
timestamp 1676037725
transform 1 0 30452 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_37
timestamp 1676037725
transform 1 0 4508 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_42
timestamp 1676037725
transform 1 0 4968 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_64
timestamp 1676037725
transform 1 0 6992 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_76
timestamp 1676037725
transform 1 0 8096 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_103
timestamp 1676037725
transform 1 0 10580 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_115
timestamp 1676037725
transform 1 0 11684 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_123
timestamp 1676037725
transform 1 0 12420 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_135
timestamp 1676037725
transform 1 0 13524 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1676037725
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_153
timestamp 1676037725
transform 1 0 15180 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_161
timestamp 1676037725
transform 1 0 15916 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_180
timestamp 1676037725
transform 1 0 17664 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_191
timestamp 1676037725
transform 1 0 18676 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1676037725
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_209
timestamp 1676037725
transform 1 0 20332 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_218
timestamp 1676037725
transform 1 0 21160 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_230
timestamp 1676037725
transform 1 0 22264 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_242
timestamp 1676037725
transform 1 0 23368 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_246
timestamp 1676037725
transform 1 0 23736 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1676037725
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_275
timestamp 1676037725
transform 1 0 26404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_302
timestamp 1676037725
transform 1 0 28888 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_309
timestamp 1676037725
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_314
timestamp 1676037725
transform 1 0 29992 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1676037725
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_27
timestamp 1676037725
transform 1 0 3588 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1676037725
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_66
timestamp 1676037725
transform 1 0 7176 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_78
timestamp 1676037725
transform 1 0 8280 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_90
timestamp 1676037725
transform 1 0 9384 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_102
timestamp 1676037725
transform 1 0 10488 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1676037725
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_137
timestamp 1676037725
transform 1 0 13708 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_144
timestamp 1676037725
transform 1 0 14352 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_156
timestamp 1676037725
transform 1 0 15456 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1676037725
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_180
timestamp 1676037725
transform 1 0 17664 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_192
timestamp 1676037725
transform 1 0 18768 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_204
timestamp 1676037725
transform 1 0 19872 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_214
timestamp 1676037725
transform 1 0 20792 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1676037725
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_238
timestamp 1676037725
transform 1 0 23000 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_262
timestamp 1676037725
transform 1 0 25208 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_272
timestamp 1676037725
transform 1 0 26128 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_286
timestamp 1676037725
transform 1 0 27416 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_294
timestamp 1676037725
transform 1 0 28152 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_317
timestamp 1676037725
transform 1 0 30268 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_35
timestamp 1676037725
transform 1 0 4324 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_39
timestamp 1676037725
transform 1 0 4692 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_66
timestamp 1676037725
transform 1 0 7176 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_73
timestamp 1676037725
transform 1 0 7820 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_81
timestamp 1676037725
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_95
timestamp 1676037725
transform 1 0 9844 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_103
timestamp 1676037725
transform 1 0 10580 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_108
timestamp 1676037725
transform 1 0 11040 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_121
timestamp 1676037725
transform 1 0 12236 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1676037725
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1676037725
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_146
timestamp 1676037725
transform 1 0 14536 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_166
timestamp 1676037725
transform 1 0 16376 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_178
timestamp 1676037725
transform 1 0 17480 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_190
timestamp 1676037725
transform 1 0 18584 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_217
timestamp 1676037725
transform 1 0 21068 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_227
timestamp 1676037725
transform 1 0 21988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_239
timestamp 1676037725
transform 1 0 23092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1676037725
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_262
timestamp 1676037725
transform 1 0 25208 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_274
timestamp 1676037725
transform 1 0 26312 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_282
timestamp 1676037725
transform 1 0 27048 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_287
timestamp 1676037725
transform 1 0 27508 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_294
timestamp 1676037725
transform 1 0 28152 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1676037725
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1676037725
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_309
timestamp 1676037725
transform 1 0 29532 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_318
timestamp 1676037725
transform 1 0 30360 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_39
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1676037725
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_79
timestamp 1676037725
transform 1 0 8372 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_91
timestamp 1676037725
transform 1 0 9476 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_103
timestamp 1676037725
transform 1 0 10580 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1676037725
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_140
timestamp 1676037725
transform 1 0 13984 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_148
timestamp 1676037725
transform 1 0 14720 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_156
timestamp 1676037725
transform 1 0 15456 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_180
timestamp 1676037725
transform 1 0 17664 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_188
timestamp 1676037725
transform 1 0 18400 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_195
timestamp 1676037725
transform 1 0 19044 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_206
timestamp 1676037725
transform 1 0 20056 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_218
timestamp 1676037725
transform 1 0 21160 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_235
timestamp 1676037725
transform 1 0 22724 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_239
timestamp 1676037725
transform 1 0 23092 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_256
timestamp 1676037725
transform 1 0 24656 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_260
timestamp 1676037725
transform 1 0 25024 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_268
timestamp 1676037725
transform 1 0 25760 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_281
timestamp 1676037725
transform 1 0 26956 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_289
timestamp 1676037725
transform 1 0 27692 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_312
timestamp 1676037725
transform 1 0 29808 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_46
timestamp 1676037725
transform 1 0 5336 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_54
timestamp 1676037725
transform 1 0 6072 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_71
timestamp 1676037725
transform 1 0 7636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_105
timestamp 1676037725
transform 1 0 10764 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_117
timestamp 1676037725
transform 1 0 11868 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_125
timestamp 1676037725
transform 1 0 12604 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_131
timestamp 1676037725
transform 1 0 13156 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1676037725
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1676037725
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_165
timestamp 1676037725
transform 1 0 16284 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_184
timestamp 1676037725
transform 1 0 18032 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_202
timestamp 1676037725
transform 1 0 19688 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_214
timestamp 1676037725
transform 1 0 20792 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_222
timestamp 1676037725
transform 1 0 21528 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_229
timestamp 1676037725
transform 1 0 22172 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1676037725
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_271
timestamp 1676037725
transform 1 0 26036 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_283
timestamp 1676037725
transform 1 0 27140 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_289
timestamp 1676037725
transform 1 0 27692 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_306
timestamp 1676037725
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_309
timestamp 1676037725
transform 1 0 29532 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_317
timestamp 1676037725
transform 1 0 30268 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_15
timestamp 1676037725
transform 1 0 2484 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_40
timestamp 1676037725
transform 1 0 4784 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1676037725
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_74
timestamp 1676037725
transform 1 0 7912 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_94
timestamp 1676037725
transform 1 0 9752 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_102
timestamp 1676037725
transform 1 0 10488 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_109
timestamp 1676037725
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_117
timestamp 1676037725
transform 1 0 11868 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_121
timestamp 1676037725
transform 1 0 12236 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_149
timestamp 1676037725
transform 1 0 14812 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_158
timestamp 1676037725
transform 1 0 15640 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_165
timestamp 1676037725
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_181
timestamp 1676037725
transform 1 0 17756 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_187
timestamp 1676037725
transform 1 0 18308 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_204
timestamp 1676037725
transform 1 0 19872 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_216
timestamp 1676037725
transform 1 0 20976 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_237
timestamp 1676037725
transform 1 0 22908 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_247
timestamp 1676037725
transform 1 0 23828 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_260
timestamp 1676037725
transform 1 0 25024 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_272
timestamp 1676037725
transform 1 0 26128 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_293
timestamp 1676037725
transform 1 0 28060 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_315
timestamp 1676037725
transform 1 0 30084 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_319
timestamp 1676037725
transform 1 0 30452 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_15
timestamp 1676037725
transform 1 0 2484 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_19
timestamp 1676037725
transform 1 0 2852 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_40
timestamp 1676037725
transform 1 0 4784 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_52
timestamp 1676037725
transform 1 0 5888 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_61
timestamp 1676037725
transform 1 0 6716 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_73
timestamp 1676037725
transform 1 0 7820 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_81
timestamp 1676037725
transform 1 0 8556 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_96
timestamp 1676037725
transform 1 0 9936 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_108
timestamp 1676037725
transform 1 0 11040 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_125
timestamp 1676037725
transform 1 0 12604 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1676037725
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_150
timestamp 1676037725
transform 1 0 14904 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_156
timestamp 1676037725
transform 1 0 15456 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_166
timestamp 1676037725
transform 1 0 16376 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_175
timestamp 1676037725
transform 1 0 17204 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_187
timestamp 1676037725
transform 1 0 18308 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1676037725
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_208
timestamp 1676037725
transform 1 0 20240 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_220
timestamp 1676037725
transform 1 0 21344 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_232
timestamp 1676037725
transform 1 0 22448 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_244
timestamp 1676037725
transform 1 0 23552 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_265
timestamp 1676037725
transform 1 0 25484 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_271
timestamp 1676037725
transform 1 0 26036 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_293
timestamp 1676037725
transform 1 0 28060 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_297
timestamp 1676037725
transform 1 0 28428 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1676037725
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1676037725
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1676037725
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_314
timestamp 1676037725
transform 1 0 29992 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_20
timestamp 1676037725
transform 1 0 2944 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_27
timestamp 1676037725
transform 1 0 3588 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1676037725
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_64
timestamp 1676037725
transform 1 0 6992 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_71
timestamp 1676037725
transform 1 0 7636 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_83
timestamp 1676037725
transform 1 0 8740 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_95
timestamp 1676037725
transform 1 0 9844 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_107
timestamp 1676037725
transform 1 0 10948 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1676037725
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_132
timestamp 1676037725
transform 1 0 13248 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_145
timestamp 1676037725
transform 1 0 14444 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1676037725
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_180
timestamp 1676037725
transform 1 0 17664 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_191
timestamp 1676037725
transform 1 0 18676 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_200
timestamp 1676037725
transform 1 0 19504 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_212
timestamp 1676037725
transform 1 0 20608 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_220
timestamp 1676037725
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_240
timestamp 1676037725
transform 1 0 23184 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_244
timestamp 1676037725
transform 1 0 23552 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_252
timestamp 1676037725
transform 1 0 24288 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_264
timestamp 1676037725
transform 1 0 25392 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_270
timestamp 1676037725
transform 1 0 25944 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_274
timestamp 1676037725
transform 1 0 26312 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_296
timestamp 1676037725
transform 1 0 28336 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_313
timestamp 1676037725
transform 1 0 29900 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_319
timestamp 1676037725
transform 1 0 30452 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_12
timestamp 1676037725
transform 1 0 2208 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_19
timestamp 1676037725
transform 1 0 2852 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1676037725
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_53
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_80
timestamp 1676037725
transform 1 0 8464 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_108
timestamp 1676037725
transform 1 0 11040 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_135
timestamp 1676037725
transform 1 0 13524 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1676037725
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_152
timestamp 1676037725
transform 1 0 15088 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_178
timestamp 1676037725
transform 1 0 17480 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_193
timestamp 1676037725
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_205
timestamp 1676037725
transform 1 0 19964 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_222
timestamp 1676037725
transform 1 0 21528 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_228
timestamp 1676037725
transform 1 0 22080 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1676037725
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1676037725
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_265
timestamp 1676037725
transform 1 0 25484 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_273
timestamp 1676037725
transform 1 0 26220 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_278
timestamp 1676037725
transform 1 0 26680 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_290
timestamp 1676037725
transform 1 0 27784 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_302
timestamp 1676037725
transform 1 0 28888 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_309
timestamp 1676037725
transform 1 0 29532 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_317
timestamp 1676037725
transform 1 0 30268 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_9
timestamp 1676037725
transform 1 0 1932 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_33
timestamp 1676037725
transform 1 0 4140 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_41
timestamp 1676037725
transform 1 0 4876 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_46
timestamp 1676037725
transform 1 0 5336 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_53
timestamp 1676037725
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_62
timestamp 1676037725
transform 1 0 6808 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_89
timestamp 1676037725
transform 1 0 9292 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_96
timestamp 1676037725
transform 1 0 9936 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_108
timestamp 1676037725
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_117
timestamp 1676037725
transform 1 0 11868 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_127
timestamp 1676037725
transform 1 0 12788 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_148
timestamp 1676037725
transform 1 0 14720 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_152
timestamp 1676037725
transform 1 0 15088 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1676037725
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1676037725
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_198
timestamp 1676037725
transform 1 0 19320 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_218
timestamp 1676037725
transform 1 0 21160 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_236
timestamp 1676037725
transform 1 0 22816 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_248
timestamp 1676037725
transform 1 0 23920 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_256
timestamp 1676037725
transform 1 0 24656 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_267
timestamp 1676037725
transform 1 0 25668 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1676037725
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1676037725
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1676037725
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_305
timestamp 1676037725
transform 1 0 29164 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_311
timestamp 1676037725
transform 1 0 29716 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_318
timestamp 1676037725
transform 1 0 30360 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_11
timestamp 1676037725
transform 1 0 2116 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_16
timestamp 1676037725
transform 1 0 2576 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_22
timestamp 1676037725
transform 1 0 3128 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1676037725
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1676037725
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1676037725
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_65
timestamp 1676037725
transform 1 0 7084 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_69
timestamp 1676037725
transform 1 0 7452 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_73
timestamp 1676037725
transform 1 0 7820 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1676037725
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_90
timestamp 1676037725
transform 1 0 9384 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_102
timestamp 1676037725
transform 1 0 10488 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_114
timestamp 1676037725
transform 1 0 11592 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_126
timestamp 1676037725
transform 1 0 12696 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1676037725
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_149
timestamp 1676037725
transform 1 0 14812 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_172
timestamp 1676037725
transform 1 0 16928 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_187
timestamp 1676037725
transform 1 0 18308 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1676037725
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_208
timestamp 1676037725
transform 1 0 20240 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1676037725
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1676037725
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1676037725
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1676037725
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_275
timestamp 1676037725
transform 1 0 26404 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_283
timestamp 1676037725
transform 1 0 27140 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_292
timestamp 1676037725
transform 1 0 27968 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_299
timestamp 1676037725
transform 1 0 28612 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1676037725
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1676037725
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_318
timestamp 1676037725
transform 1 0 30360 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_7
timestamp 1676037725
transform 1 0 1748 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_31
timestamp 1676037725
transform 1 0 3956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_43
timestamp 1676037725
transform 1 0 5060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1676037725
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1676037725
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1676037725
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1676037725
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1676037725
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1676037725
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_125
timestamp 1676037725
transform 1 0 12604 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_145
timestamp 1676037725
transform 1 0 14444 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1676037725
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_181
timestamp 1676037725
transform 1 0 17756 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_190
timestamp 1676037725
transform 1 0 18584 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_202
timestamp 1676037725
transform 1 0 19688 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_214
timestamp 1676037725
transform 1 0 20792 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1676037725
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_237
timestamp 1676037725
transform 1 0 22908 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_246
timestamp 1676037725
transform 1 0 23736 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_270
timestamp 1676037725
transform 1 0 25944 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1676037725
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_281
timestamp 1676037725
transform 1 0 26956 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_287
timestamp 1676037725
transform 1 0 27508 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_295
timestamp 1676037725
transform 1 0 28244 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_301
timestamp 1676037725
transform 1 0 28796 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_308
timestamp 1676037725
transform 1 0 29440 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_11
timestamp 1676037725
transform 1 0 2116 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_17
timestamp 1676037725
transform 1 0 2668 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_24
timestamp 1676037725
transform 1 0 3312 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_34
timestamp 1676037725
transform 1 0 4232 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_42
timestamp 1676037725
transform 1 0 4968 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_49
timestamp 1676037725
transform 1 0 5612 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_66
timestamp 1676037725
transform 1 0 7176 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_78
timestamp 1676037725
transform 1 0 8280 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_100
timestamp 1676037725
transform 1 0 10304 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_112
timestamp 1676037725
transform 1 0 11408 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_124
timestamp 1676037725
transform 1 0 12512 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1676037725
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1676037725
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1676037725
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_177
timestamp 1676037725
transform 1 0 17388 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1676037725
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_205
timestamp 1676037725
transform 1 0 19964 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_209
timestamp 1676037725
transform 1 0 20332 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_231
timestamp 1676037725
transform 1 0 22356 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_243
timestamp 1676037725
transform 1 0 23460 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1676037725
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1676037725
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_277
timestamp 1676037725
transform 1 0 26588 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_283
timestamp 1676037725
transform 1 0 27140 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_300
timestamp 1676037725
transform 1 0 28704 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_309
timestamp 1676037725
transform 1 0 29532 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_317
timestamp 1676037725
transform 1 0 30268 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_35
timestamp 1676037725
transform 1 0 4324 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_42
timestamp 1676037725
transform 1 0 4968 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_50
timestamp 1676037725
transform 1 0 5704 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1676037725
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_80
timestamp 1676037725
transform 1 0 8464 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_102
timestamp 1676037725
transform 1 0 10488 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1676037725
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1676037725
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_137
timestamp 1676037725
transform 1 0 13708 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_33_148
timestamp 1676037725
transform 1 0 14720 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_154
timestamp 1676037725
transform 1 0 15272 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_158
timestamp 1676037725
transform 1 0 15640 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1676037725
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_176
timestamp 1676037725
transform 1 0 17296 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_191
timestamp 1676037725
transform 1 0 18676 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_199
timestamp 1676037725
transform 1 0 19412 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_205
timestamp 1676037725
transform 1 0 19964 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1676037725
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_230
timestamp 1676037725
transform 1 0 22264 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_242
timestamp 1676037725
transform 1 0 23368 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_257
timestamp 1676037725
transform 1 0 24748 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_269
timestamp 1676037725
transform 1 0 25852 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_277
timestamp 1676037725
transform 1 0 26588 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1676037725
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1676037725
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1676037725
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_317
timestamp 1676037725
transform 1 0 30268 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_15
timestamp 1676037725
transform 1 0 2484 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_19
timestamp 1676037725
transform 1 0 2852 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1676037725
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_36
timestamp 1676037725
transform 1 0 4416 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_44
timestamp 1676037725
transform 1 0 5152 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_49
timestamp 1676037725
transform 1 0 5612 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_74
timestamp 1676037725
transform 1 0 7912 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1676037725
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_89
timestamp 1676037725
transform 1 0 9292 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_99
timestamp 1676037725
transform 1 0 10212 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_119
timestamp 1676037725
transform 1 0 12052 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_126
timestamp 1676037725
transform 1 0 12696 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1676037725
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_145
timestamp 1676037725
transform 1 0 14444 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_155
timestamp 1676037725
transform 1 0 15364 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_159
timestamp 1676037725
transform 1 0 15732 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_169
timestamp 1676037725
transform 1 0 16652 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_182
timestamp 1676037725
transform 1 0 17848 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_193
timestamp 1676037725
transform 1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_209
timestamp 1676037725
transform 1 0 20332 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_231
timestamp 1676037725
transform 1 0 22356 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_243
timestamp 1676037725
transform 1 0 23460 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1676037725
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_271
timestamp 1676037725
transform 1 0 26036 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_282
timestamp 1676037725
transform 1 0 27048 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_290
timestamp 1676037725
transform 1 0 27784 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_305
timestamp 1676037725
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_309
timestamp 1676037725
transform 1 0 29532 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_317
timestamp 1676037725
transform 1 0 30268 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_15
timestamp 1676037725
transform 1 0 2484 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_36
timestamp 1676037725
transform 1 0 4416 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_48
timestamp 1676037725
transform 1 0 5520 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1676037725
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_75
timestamp 1676037725
transform 1 0 8004 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_83
timestamp 1676037725
transform 1 0 8740 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_102
timestamp 1676037725
transform 1 0 10488 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1676037725
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_119
timestamp 1676037725
transform 1 0 12052 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_128
timestamp 1676037725
transform 1 0 12880 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_140
timestamp 1676037725
transform 1 0 13984 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_148
timestamp 1676037725
transform 1 0 14720 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1676037725
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_180
timestamp 1676037725
transform 1 0 17664 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_189
timestamp 1676037725
transform 1 0 18492 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_201
timestamp 1676037725
transform 1 0 19596 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_213
timestamp 1676037725
transform 1 0 20700 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_221
timestamp 1676037725
transform 1 0 21436 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_243
timestamp 1676037725
transform 1 0 23460 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_255
timestamp 1676037725
transform 1 0 24564 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_265
timestamp 1676037725
transform 1 0 25484 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_275
timestamp 1676037725
transform 1 0 26404 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1676037725
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_281
timestamp 1676037725
transform 1 0 26956 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_287
timestamp 1676037725
transform 1 0 27508 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_309
timestamp 1676037725
transform 1 0 29532 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_317
timestamp 1676037725
transform 1 0 30268 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_9
timestamp 1676037725
transform 1 0 1932 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1676037725
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_43
timestamp 1676037725
transform 1 0 5060 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_47
timestamp 1676037725
transform 1 0 5428 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_51
timestamp 1676037725
transform 1 0 5796 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_68
timestamp 1676037725
transform 1 0 7360 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_80
timestamp 1676037725
transform 1 0 8464 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_93
timestamp 1676037725
transform 1 0 9660 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_102
timestamp 1676037725
transform 1 0 10488 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_106
timestamp 1676037725
transform 1 0 10856 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_116
timestamp 1676037725
transform 1 0 11776 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_123
timestamp 1676037725
transform 1 0 12420 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_132
timestamp 1676037725
transform 1 0 13248 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_153
timestamp 1676037725
transform 1 0 15180 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_173
timestamp 1676037725
transform 1 0 17020 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_183
timestamp 1676037725
transform 1 0 17940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1676037725
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_209
timestamp 1676037725
transform 1 0 20332 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_215
timestamp 1676037725
transform 1 0 20884 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_232
timestamp 1676037725
transform 1 0 22448 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_242
timestamp 1676037725
transform 1 0 23368 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1676037725
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_266
timestamp 1676037725
transform 1 0 25576 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_277
timestamp 1676037725
transform 1 0 26588 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_285
timestamp 1676037725
transform 1 0 27324 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_289
timestamp 1676037725
transform 1 0 27692 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_306
timestamp 1676037725
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_309
timestamp 1676037725
transform 1 0 29532 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_318
timestamp 1676037725
transform 1 0 30360 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_13
timestamp 1676037725
transform 1 0 2300 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_33
timestamp 1676037725
transform 1 0 4140 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_43
timestamp 1676037725
transform 1 0 5060 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_52
timestamp 1676037725
transform 1 0 5888 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_62
timestamp 1676037725
transform 1 0 6808 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_84
timestamp 1676037725
transform 1 0 8832 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_95
timestamp 1676037725
transform 1 0 9844 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_107
timestamp 1676037725
transform 1 0 10948 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1676037725
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_124
timestamp 1676037725
transform 1 0 12512 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_132
timestamp 1676037725
transform 1 0 13248 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_144
timestamp 1676037725
transform 1 0 14352 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_153
timestamp 1676037725
transform 1 0 15180 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1676037725
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_182
timestamp 1676037725
transform 1 0 17848 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_190
timestamp 1676037725
transform 1 0 18584 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_209
timestamp 1676037725
transform 1 0 20332 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_217
timestamp 1676037725
transform 1 0 21068 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1676037725
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_236
timestamp 1676037725
transform 1 0 22816 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_245
timestamp 1676037725
transform 1 0 23644 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_253
timestamp 1676037725
transform 1 0 24380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_270
timestamp 1676037725
transform 1 0 25944 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1676037725
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1676037725
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_293
timestamp 1676037725
transform 1 0 28060 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_317
timestamp 1676037725
transform 1 0 30268 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_9
timestamp 1676037725
transform 1 0 1932 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_23
timestamp 1676037725
transform 1 0 3220 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1676037725
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_37
timestamp 1676037725
transform 1 0 4508 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_45
timestamp 1676037725
transform 1 0 5244 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_72
timestamp 1676037725
transform 1 0 7728 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_94
timestamp 1676037725
transform 1 0 9752 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_100
timestamp 1676037725
transform 1 0 10304 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_121
timestamp 1676037725
transform 1 0 12236 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_132
timestamp 1676037725
transform 1 0 13248 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_153
timestamp 1676037725
transform 1 0 15180 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1676037725
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1676037725
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1676037725
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1676037725
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_208
timestamp 1676037725
transform 1 0 20240 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_234
timestamp 1676037725
transform 1 0 22632 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_246
timestamp 1676037725
transform 1 0 23736 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_271
timestamp 1676037725
transform 1 0 26036 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_282
timestamp 1676037725
transform 1 0 27048 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_294
timestamp 1676037725
transform 1 0 28152 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_299
timestamp 1676037725
transform 1 0 28612 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_306
timestamp 1676037725
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_309
timestamp 1676037725
transform 1 0 29532 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_317
timestamp 1676037725
transform 1 0 30268 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_15
timestamp 1676037725
transform 1 0 2484 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_32
timestamp 1676037725
transform 1 0 4048 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_40
timestamp 1676037725
transform 1 0 4784 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_47
timestamp 1676037725
transform 1 0 5428 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1676037725
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_69
timestamp 1676037725
transform 1 0 7452 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_93
timestamp 1676037725
transform 1 0 9660 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_97
timestamp 1676037725
transform 1 0 10028 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_104
timestamp 1676037725
transform 1 0 10672 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_128
timestamp 1676037725
transform 1 0 12880 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_132
timestamp 1676037725
transform 1 0 13248 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_136
timestamp 1676037725
transform 1 0 13616 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_143
timestamp 1676037725
transform 1 0 14260 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_149
timestamp 1676037725
transform 1 0 14812 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1676037725
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_181
timestamp 1676037725
transform 1 0 17756 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_205
timestamp 1676037725
transform 1 0 19964 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_213
timestamp 1676037725
transform 1 0 20700 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_221
timestamp 1676037725
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_236
timestamp 1676037725
transform 1 0 22816 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_262
timestamp 1676037725
transform 1 0 25208 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_270
timestamp 1676037725
transform 1 0 25944 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_277
timestamp 1676037725
transform 1 0 26588 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1676037725
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_293
timestamp 1676037725
transform 1 0 28060 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_298
timestamp 1676037725
transform 1 0 28520 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_310
timestamp 1676037725
transform 1 0 29624 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_318
timestamp 1676037725
transform 1 0 30360 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_11
timestamp 1676037725
transform 1 0 2116 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_16
timestamp 1676037725
transform 1 0 2576 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1676037725
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_36
timestamp 1676037725
transform 1 0 4416 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_45
timestamp 1676037725
transform 1 0 5244 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_57
timestamp 1676037725
transform 1 0 6348 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_72
timestamp 1676037725
transform 1 0 7728 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1676037725
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_109
timestamp 1676037725
transform 1 0 11132 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_134
timestamp 1676037725
transform 1 0 13432 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_164
timestamp 1676037725
transform 1 0 16192 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_176
timestamp 1676037725
transform 1 0 17296 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_191
timestamp 1676037725
transform 1 0 18676 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1676037725
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_208
timestamp 1676037725
transform 1 0 20240 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_236
timestamp 1676037725
transform 1 0 22816 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1676037725
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1676037725
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_264
timestamp 1676037725
transform 1 0 25392 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_276
timestamp 1676037725
transform 1 0 26496 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_288
timestamp 1676037725
transform 1 0 27600 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_292
timestamp 1676037725
transform 1 0 27968 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_306
timestamp 1676037725
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_309
timestamp 1676037725
transform 1 0 29532 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_317
timestamp 1676037725
transform 1 0 30268 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_3
timestamp 1676037725
transform 1 0 1380 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_22
timestamp 1676037725
transform 1 0 3128 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_46
timestamp 1676037725
transform 1 0 5336 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_50
timestamp 1676037725
transform 1 0 5704 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_54
timestamp 1676037725
transform 1 0 6072 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_57
timestamp 1676037725
transform 1 0 6348 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_72
timestamp 1676037725
transform 1 0 7728 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_85
timestamp 1676037725
transform 1 0 8924 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_97
timestamp 1676037725
transform 1 0 10028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_109
timestamp 1676037725
transform 1 0 11132 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_113
timestamp 1676037725
transform 1 0 11500 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_119
timestamp 1676037725
transform 1 0 12052 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_126
timestamp 1676037725
transform 1 0 12696 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_138
timestamp 1676037725
transform 1 0 13800 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_153
timestamp 1676037725
transform 1 0 15180 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_164
timestamp 1676037725
transform 1 0 16192 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_169
timestamp 1676037725
transform 1 0 16652 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_175
timestamp 1676037725
transform 1 0 17204 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_192
timestamp 1676037725
transform 1 0 18768 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_200
timestamp 1676037725
transform 1 0 19504 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_210
timestamp 1676037725
transform 1 0 20424 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1676037725
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_225
timestamp 1676037725
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_231
timestamp 1676037725
transform 1 0 22356 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_239
timestamp 1676037725
transform 1 0 23092 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_261
timestamp 1676037725
transform 1 0 25116 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_272
timestamp 1676037725
transform 1 0 26128 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1676037725
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_293
timestamp 1676037725
transform 1 0 28060 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_315
timestamp 1676037725
transform 1 0 30084 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_319
timestamp 1676037725
transform 1 0 30452 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1676037725
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_15
timestamp 1676037725
transform 1 0 2484 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_24
timestamp 1676037725
transform 1 0 3312 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_29
timestamp 1676037725
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_34
timestamp 1676037725
transform 1 0 4232 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_46
timestamp 1676037725
transform 1 0 5336 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_58
timestamp 1676037725
transform 1 0 6440 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1676037725
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1676037725
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_85
timestamp 1676037725
transform 1 0 8924 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_100
timestamp 1676037725
transform 1 0 10304 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_104
timestamp 1676037725
transform 1 0 10672 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_125
timestamp 1676037725
transform 1 0 12604 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_137
timestamp 1676037725
transform 1 0 13708 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1676037725
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1676037725
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1676037725
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1676037725
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1676037725
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1676037725
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1676037725
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_206
timestamp 1676037725
transform 1 0 20056 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_218
timestamp 1676037725
transform 1 0 21160 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_230
timestamp 1676037725
transform 1 0 22264 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_234
timestamp 1676037725
transform 1 0 22632 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_238
timestamp 1676037725
transform 1 0 23000 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1676037725
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_253
timestamp 1676037725
transform 1 0 24380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_266
timestamp 1676037725
transform 1 0 25576 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1676037725
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_289
timestamp 1676037725
transform 1 0 27692 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_294
timestamp 1676037725
transform 1 0 28152 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1676037725
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1676037725
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_309
timestamp 1676037725
transform 1 0 29532 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_318
timestamp 1676037725
transform 1 0 30360 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1676037725
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_15
timestamp 1676037725
transform 1 0 2484 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_36
timestamp 1676037725
transform 1 0 4416 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_48
timestamp 1676037725
transform 1 0 5520 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_57
timestamp 1676037725
transform 1 0 6348 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_80
timestamp 1676037725
transform 1 0 8464 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_100
timestamp 1676037725
transform 1 0 10304 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_113
timestamp 1676037725
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_124
timestamp 1676037725
transform 1 0 12512 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_134
timestamp 1676037725
transform 1 0 13432 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_146
timestamp 1676037725
transform 1 0 14536 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_158
timestamp 1676037725
transform 1 0 15640 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_166
timestamp 1676037725
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1676037725
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_181
timestamp 1676037725
transform 1 0 17756 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_187
timestamp 1676037725
transform 1 0 18308 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_211
timestamp 1676037725
transform 1 0 20516 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_218
timestamp 1676037725
transform 1 0 21160 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_225
timestamp 1676037725
transform 1 0 21804 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_229
timestamp 1676037725
transform 1 0 22172 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_239
timestamp 1676037725
transform 1 0 23092 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_251
timestamp 1676037725
transform 1 0 24196 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_271
timestamp 1676037725
transform 1 0 26036 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1676037725
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1676037725
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_293
timestamp 1676037725
transform 1 0 28060 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_315
timestamp 1676037725
transform 1 0 30084 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_319
timestamp 1676037725
transform 1 0 30452 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1676037725
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_15
timestamp 1676037725
transform 1 0 2484 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_21
timestamp 1676037725
transform 1 0 3036 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_26
timestamp 1676037725
transform 1 0 3496 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_29
timestamp 1676037725
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_39
timestamp 1676037725
transform 1 0 4692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_51
timestamp 1676037725
transform 1 0 5796 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_68
timestamp 1676037725
transform 1 0 7360 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_79
timestamp 1676037725
transform 1 0 8372 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1676037725
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1676037725
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_94
timestamp 1676037725
transform 1 0 9752 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_106
timestamp 1676037725
transform 1 0 10856 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_125
timestamp 1676037725
transform 1 0 12604 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_137
timestamp 1676037725
transform 1 0 13708 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_141
timestamp 1676037725
transform 1 0 14076 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_145
timestamp 1676037725
transform 1 0 14444 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_153
timestamp 1676037725
transform 1 0 15180 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_166
timestamp 1676037725
transform 1 0 16376 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_178
timestamp 1676037725
transform 1 0 17480 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_193
timestamp 1676037725
transform 1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1676037725
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_212
timestamp 1676037725
transform 1 0 20608 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_224
timestamp 1676037725
transform 1 0 21712 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_241
timestamp 1676037725
transform 1 0 23276 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_249
timestamp 1676037725
transform 1 0 24012 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_253
timestamp 1676037725
transform 1 0 24380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_257
timestamp 1676037725
transform 1 0 24748 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_267
timestamp 1676037725
transform 1 0 25668 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1676037725
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_289
timestamp 1676037725
transform 1 0 27692 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_306
timestamp 1676037725
transform 1 0 29256 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_309
timestamp 1676037725
transform 1 0 29532 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_314
timestamp 1676037725
transform 1 0 29992 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1676037725
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_15
timestamp 1676037725
transform 1 0 2484 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_35
timestamp 1676037725
transform 1 0 4324 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_45
timestamp 1676037725
transform 1 0 5244 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_53
timestamp 1676037725
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_57
timestamp 1676037725
transform 1 0 6348 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_63
timestamp 1676037725
transform 1 0 6900 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_70
timestamp 1676037725
transform 1 0 7544 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_82
timestamp 1676037725
transform 1 0 8648 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_94
timestamp 1676037725
transform 1 0 9752 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_106
timestamp 1676037725
transform 1 0 10856 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_113
timestamp 1676037725
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_122
timestamp 1676037725
transform 1 0 12328 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_45_143
timestamp 1676037725
transform 1 0 14260 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_149
timestamp 1676037725
transform 1 0 14812 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1676037725
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1676037725
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_181
timestamp 1676037725
transform 1 0 17756 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_200
timestamp 1676037725
transform 1 0 19504 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_212
timestamp 1676037725
transform 1 0 20608 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1676037725
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_237
timestamp 1676037725
transform 1 0 22908 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_45_250
timestamp 1676037725
transform 1 0 24104 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_45_272
timestamp 1676037725
transform 1 0 26128 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1676037725
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_293
timestamp 1676037725
transform 1 0 28060 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_317
timestamp 1676037725
transform 1 0 30268 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_3
timestamp 1676037725
transform 1 0 1380 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_16
timestamp 1676037725
transform 1 0 2576 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_26
timestamp 1676037725
transform 1 0 3496 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1676037725
transform 1 0 3772 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_47
timestamp 1676037725
transform 1 0 5428 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_55
timestamp 1676037725
transform 1 0 6164 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_59
timestamp 1676037725
transform 1 0 6532 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_81
timestamp 1676037725
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_85
timestamp 1676037725
transform 1 0 8924 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_100
timestamp 1676037725
transform 1 0 10304 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_127
timestamp 1676037725
transform 1 0 12788 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1676037725
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_141
timestamp 1676037725
transform 1 0 14076 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_158
timestamp 1676037725
transform 1 0 15640 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_170
timestamp 1676037725
transform 1 0 16744 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_178
timestamp 1676037725
transform 1 0 17480 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1676037725
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1676037725
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_202
timestamp 1676037725
transform 1 0 19688 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_210
timestamp 1676037725
transform 1 0 20424 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_232
timestamp 1676037725
transform 1 0 22448 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_239
timestamp 1676037725
transform 1 0 23092 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_246
timestamp 1676037725
transform 1 0 23736 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1676037725
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_272
timestamp 1676037725
transform 1 0 26128 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_279
timestamp 1676037725
transform 1 0 26772 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_296
timestamp 1676037725
transform 1 0 28336 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_303
timestamp 1676037725
transform 1 0 28980 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1676037725
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_309
timestamp 1676037725
transform 1 0 29532 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_317
timestamp 1676037725
transform 1 0 30268 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1676037725
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_15
timestamp 1676037725
transform 1 0 2484 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_33
timestamp 1676037725
transform 1 0 4140 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_47_53
timestamp 1676037725
transform 1 0 5980 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_57
timestamp 1676037725
transform 1 0 6348 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_74
timestamp 1676037725
transform 1 0 7912 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_99
timestamp 1676037725
transform 1 0 10212 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_110
timestamp 1676037725
transform 1 0 11224 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_113
timestamp 1676037725
transform 1 0 11500 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_140
timestamp 1676037725
transform 1 0 13984 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_47_165
timestamp 1676037725
transform 1 0 16284 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_169
timestamp 1676037725
transform 1 0 16652 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_180
timestamp 1676037725
transform 1 0 17664 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_205
timestamp 1676037725
transform 1 0 19964 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_222
timestamp 1676037725
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_225
timestamp 1676037725
transform 1 0 21804 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_231
timestamp 1676037725
transform 1 0 22356 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_253
timestamp 1676037725
transform 1 0 24380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_265
timestamp 1676037725
transform 1 0 25484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_277
timestamp 1676037725
transform 1 0 26588 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_281
timestamp 1676037725
transform 1 0 26956 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_304
timestamp 1676037725
transform 1 0 29072 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_311
timestamp 1676037725
transform 1 0 29716 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_319
timestamp 1676037725
transform 1 0 30452 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1676037725
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_15
timestamp 1676037725
transform 1 0 2484 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_21
timestamp 1676037725
transform 1 0 3036 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_26
timestamp 1676037725
transform 1 0 3496 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_29
timestamp 1676037725
transform 1 0 3772 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_43
timestamp 1676037725
transform 1 0 5060 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_55
timestamp 1676037725
transform 1 0 6164 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_67
timestamp 1676037725
transform 1 0 7268 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_73
timestamp 1676037725
transform 1 0 7820 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_80
timestamp 1676037725
transform 1 0 8464 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_85
timestamp 1676037725
transform 1 0 8924 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_89
timestamp 1676037725
transform 1 0 9292 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_93
timestamp 1676037725
transform 1 0 9660 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_99
timestamp 1676037725
transform 1 0 10212 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_103
timestamp 1676037725
transform 1 0 10580 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_120
timestamp 1676037725
transform 1 0 12144 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_127
timestamp 1676037725
transform 1 0 12788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1676037725
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_141
timestamp 1676037725
transform 1 0 14076 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_150
timestamp 1676037725
transform 1 0 14904 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_157
timestamp 1676037725
transform 1 0 15548 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_169
timestamp 1676037725
transform 1 0 16652 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_181
timestamp 1676037725
transform 1 0 17756 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_191
timestamp 1676037725
transform 1 0 18676 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1676037725
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1676037725
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_209
timestamp 1676037725
transform 1 0 20332 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_213
timestamp 1676037725
transform 1 0 20700 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_217
timestamp 1676037725
transform 1 0 21068 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_221
timestamp 1676037725
transform 1 0 21436 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_225
timestamp 1676037725
transform 1 0 21804 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_233
timestamp 1676037725
transform 1 0 22540 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_247
timestamp 1676037725
transform 1 0 23828 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1676037725
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1676037725
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1676037725
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_277
timestamp 1676037725
transform 1 0 26588 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_281
timestamp 1676037725
transform 1 0 26956 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_285
timestamp 1676037725
transform 1 0 27324 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_306
timestamp 1676037725
transform 1 0 29256 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_309
timestamp 1676037725
transform 1 0 29532 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_317
timestamp 1676037725
transform 1 0 30268 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1676037725
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_15
timestamp 1676037725
transform 1 0 2484 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_21
timestamp 1676037725
transform 1 0 3036 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_25
timestamp 1676037725
transform 1 0 3404 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_29
timestamp 1676037725
transform 1 0 3772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_41
timestamp 1676037725
transform 1 0 4876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_53
timestamp 1676037725
transform 1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_57
timestamp 1676037725
transform 1 0 6348 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_65
timestamp 1676037725
transform 1 0 7084 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_77
timestamp 1676037725
transform 1 0 8188 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_83
timestamp 1676037725
transform 1 0 8740 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_85
timestamp 1676037725
transform 1 0 8924 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_97
timestamp 1676037725
transform 1 0 10028 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_107
timestamp 1676037725
transform 1 0 10948 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1676037725
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1676037725
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1676037725
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_137
timestamp 1676037725
transform 1 0 13708 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_141
timestamp 1676037725
transform 1 0 14076 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_152
timestamp 1676037725
transform 1 0 15088 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_164
timestamp 1676037725
transform 1 0 16192 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1676037725
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_181
timestamp 1676037725
transform 1 0 17756 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_188
timestamp 1676037725
transform 1 0 18400 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_197
timestamp 1676037725
transform 1 0 19228 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_209
timestamp 1676037725
transform 1 0 20332 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_221
timestamp 1676037725
transform 1 0 21436 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1676037725
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_231
timestamp 1676037725
transform 1 0 22356 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_243
timestamp 1676037725
transform 1 0 23460 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_251
timestamp 1676037725
transform 1 0 24196 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_253
timestamp 1676037725
transform 1 0 24380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_265
timestamp 1676037725
transform 1 0 25484 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_269
timestamp 1676037725
transform 1 0 25852 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_274
timestamp 1676037725
transform 1 0 26312 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1676037725
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_293
timestamp 1676037725
transform 1 0 28060 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_306
timestamp 1676037725
transform 1 0 29256 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_309
timestamp 1676037725
transform 1 0 29532 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_318
timestamp 1676037725
transform 1 0 30360 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 30820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 30820 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 30820 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 30820 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 30820 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 30820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 30820 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 30820 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 30820 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 30820 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 30820 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 30820 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 30820 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 30820 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 30820 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 30820 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 30820 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 30820 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 30820 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 30820 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 30820 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 30820 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 30820 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 30820 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 30820 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 30820 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 30820 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 30820 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 30820 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 30820 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 30820 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 30820 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 30820 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 30820 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 30820 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 30820 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 30820 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 30820 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 30820 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 30820 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 30820 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1676037725
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1676037725
transform -1 0 30820 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1676037725
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1676037725
transform -1 0 30820 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1676037725
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1676037725
transform -1 0 30820 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1676037725
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1676037725
transform -1 0 30820 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1676037725
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1676037725
transform -1 0 30820 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1676037725
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1676037725
transform -1 0 30820 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1676037725
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1676037725
transform -1 0 30820 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1676037725
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1676037725
transform -1 0 30820 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1676037725
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1676037725
transform -1 0 30820 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 3680 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 8832 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 13984 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 19136 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 24288 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 29440 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _308_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10856 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _309_
timestamp 1676037725
transform -1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 1676037725
transform 1 0 4692 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _311_
timestamp 1676037725
transform -1 0 27508 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _312_
timestamp 1676037725
transform -1 0 24104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _313_
timestamp 1676037725
transform -1 0 23000 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _314_
timestamp 1676037725
transform -1 0 22264 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _315_
timestamp 1676037725
transform -1 0 19964 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _316_
timestamp 1676037725
transform -1 0 17940 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _317_
timestamp 1676037725
transform -1 0 16376 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _318_
timestamp 1676037725
transform -1 0 26680 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _319_
timestamp 1676037725
transform 1 0 28520 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _320_
timestamp 1676037725
transform 1 0 27416 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _321_
timestamp 1676037725
transform -1 0 29992 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _322_
timestamp 1676037725
transform -1 0 23000 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _323_
timestamp 1676037725
transform -1 0 25484 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _324_
timestamp 1676037725
transform 1 0 28888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _325_
timestamp 1676037725
transform -1 0 28612 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _326_
timestamp 1676037725
transform 1 0 28980 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _327_
timestamp 1676037725
transform -1 0 4324 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _328_
timestamp 1676037725
transform -1 0 5060 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _329_
timestamp 1676037725
transform -1 0 5336 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _330_
timestamp 1676037725
transform 1 0 7544 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _331_
timestamp 1676037725
transform 1 0 10948 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _332_
timestamp 1676037725
transform 1 0 8280 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _333_
timestamp 1676037725
transform 1 0 6532 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _334_
timestamp 1676037725
transform -1 0 6808 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _335_
timestamp 1676037725
transform -1 0 9384 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _336_
timestamp 1676037725
transform -1 0 11224 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _337_
timestamp 1676037725
transform 1 0 9844 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _338_
timestamp 1676037725
transform -1 0 28612 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _339_
timestamp 1676037725
transform -1 0 23092 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _340_
timestamp 1676037725
transform 1 0 20792 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _341_
timestamp 1676037725
transform -1 0 17664 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _342_
timestamp 1676037725
transform 1 0 20884 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _343_
timestamp 1676037725
transform -1 0 22264 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _344_
timestamp 1676037725
transform 1 0 27416 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 1676037725
transform -1 0 29256 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp 1676037725
transform -1 0 28796 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 1676037725
transform -1 0 29992 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _348_
timestamp 1676037725
transform 1 0 27048 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _349_
timestamp 1676037725
transform 1 0 29440 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _350_
timestamp 1676037725
transform -1 0 18584 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _351_
timestamp 1676037725
transform -1 0 13800 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _352_
timestamp 1676037725
transform 1 0 14628 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _353_
timestamp 1676037725
transform 1 0 13984 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _354_
timestamp 1676037725
transform -1 0 12052 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _355_
timestamp 1676037725
transform 1 0 5796 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _356_
timestamp 1676037725
transform 1 0 5796 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _357_
timestamp 1676037725
transform -1 0 6808 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _358_
timestamp 1676037725
transform -1 0 6900 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _359_
timestamp 1676037725
transform -1 0 7820 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _360_
timestamp 1676037725
transform -1 0 9660 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _361_
timestamp 1676037725
transform -1 0 11224 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _362_
timestamp 1676037725
transform -1 0 7820 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _363_
timestamp 1676037725
transform 1 0 6716 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _364_
timestamp 1676037725
transform -1 0 14536 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _365_
timestamp 1676037725
transform -1 0 2668 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _366_
timestamp 1676037725
transform -1 0 2208 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _367_
timestamp 1676037725
transform -1 0 2944 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _368_
timestamp 1676037725
transform 1 0 4508 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _369_
timestamp 1676037725
transform -1 0 9936 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _370_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15548 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _371_
timestamp 1676037725
transform 1 0 16928 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _372_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 20240 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _373_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25300 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _374_
timestamp 1676037725
transform 1 0 24932 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _375_
timestamp 1676037725
transform 1 0 24840 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _376_
timestamp 1676037725
transform 1 0 24656 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_8  _377_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4508 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_2  _378_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _379__1
timestamp 1676037725
transform -1 0 12236 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _379__2
timestamp 1676037725
transform -1 0 11040 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _380_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15180 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _381_
timestamp 1676037725
transform -1 0 16192 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _382_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12052 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _383_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12420 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _384_
timestamp 1676037725
transform 1 0 9200 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _385_
timestamp 1676037725
transform 1 0 9108 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _386_
timestamp 1676037725
transform 1 0 9108 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _387_
timestamp 1676037725
transform -1 0 13248 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _388_
timestamp 1676037725
transform 1 0 12144 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _389_
timestamp 1676037725
transform 1 0 9844 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _390_
timestamp 1676037725
transform -1 0 13248 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _391_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10120 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _392_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12144 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _393_
timestamp 1676037725
transform 1 0 7728 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _394_
timestamp 1676037725
transform 1 0 11684 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _395_
timestamp 1676037725
transform 1 0 12880 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _396_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 13248 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_4  _397_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16376 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__o211ai_4  _398_
timestamp 1676037725
transform 1 0 14812 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _399_
timestamp 1676037725
transform -1 0 15640 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_2  _400_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14536 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_2  _401_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10948 0 1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _402_
timestamp 1676037725
transform 1 0 20792 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _403_
timestamp 1676037725
transform -1 0 26588 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _404_
timestamp 1676037725
transform 1 0 19412 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _405_
timestamp 1676037725
transform 1 0 23184 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _406_
timestamp 1676037725
transform 1 0 22724 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _407_
timestamp 1676037725
transform 1 0 25484 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _408_
timestamp 1676037725
transform 1 0 23460 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _409_
timestamp 1676037725
transform 1 0 19780 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _410_
timestamp 1676037725
transform 1 0 25944 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _411_
timestamp 1676037725
transform -1 0 27048 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _412_
timestamp 1676037725
transform -1 0 26588 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _413_
timestamp 1676037725
transform 1 0 21252 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _414_
timestamp 1676037725
transform -1 0 23644 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _415_
timestamp 1676037725
transform 1 0 23000 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _416_
timestamp 1676037725
transform 1 0 25484 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _417_
timestamp 1676037725
transform 1 0 26036 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_2  _418_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 26496 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_4  _419_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17296 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__and3b_1  _420_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18032 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _421_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18216 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _422_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28060 0 1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _423_
timestamp 1676037725
transform -1 0 12512 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _424_
timestamp 1676037725
transform 1 0 12972 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _425_
timestamp 1676037725
transform -1 0 14168 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _426_
timestamp 1676037725
transform -1 0 13524 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _427_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 13524 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _428_
timestamp 1676037725
transform 1 0 9200 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _429_
timestamp 1676037725
transform 1 0 11868 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _430_
timestamp 1676037725
transform -1 0 13156 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _431_
timestamp 1676037725
transform -1 0 8924 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _432_
timestamp 1676037725
transform -1 0 8004 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _433_
timestamp 1676037725
transform 1 0 8188 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _434_
timestamp 1676037725
transform 1 0 9384 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _435_
timestamp 1676037725
transform 1 0 7268 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _436_
timestamp 1676037725
transform -1 0 7176 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _437_
timestamp 1676037725
transform 1 0 6532 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _438_
timestamp 1676037725
transform 1 0 9108 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _439_
timestamp 1676037725
transform 1 0 7544 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _440_
timestamp 1676037725
transform 1 0 10396 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _441_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12144 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _442_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 12604 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _443_
timestamp 1676037725
transform -1 0 17664 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_4  _444_
timestamp 1676037725
transform -1 0 16192 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__a21boi_1  _445_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13248 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_2  _446_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11408 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _447_
timestamp 1676037725
transform 1 0 9844 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _448_
timestamp 1676037725
transform -1 0 21528 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _449_
timestamp 1676037725
transform -1 0 22172 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _450_
timestamp 1676037725
transform 1 0 25116 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _451_
timestamp 1676037725
transform 1 0 18032 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _452_
timestamp 1676037725
transform 1 0 23644 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _453_
timestamp 1676037725
transform 1 0 19412 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _454_
timestamp 1676037725
transform 1 0 22356 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _455_
timestamp 1676037725
transform 1 0 20700 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _456_
timestamp 1676037725
transform 1 0 20516 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _457_
timestamp 1676037725
transform 1 0 19412 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _458_
timestamp 1676037725
transform 1 0 21436 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _459_
timestamp 1676037725
transform 1 0 19412 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _460_
timestamp 1676037725
transform 1 0 18584 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _461_
timestamp 1676037725
transform 1 0 20424 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _462_
timestamp 1676037725
transform 1 0 24564 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _463_
timestamp 1676037725
transform 1 0 25576 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_2  _464_
timestamp 1676037725
transform 1 0 21988 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _465_
timestamp 1676037725
transform 1 0 18860 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _466_
timestamp 1676037725
transform -1 0 18676 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _467_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17572 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_2  _468_
timestamp 1676037725
transform 1 0 28888 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__and4_2  _469_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26864 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _470_
timestamp 1676037725
transform 1 0 27968 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _471_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27416 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _472_
timestamp 1676037725
transform -1 0 30360 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _473_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29072 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _474_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27692 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _475_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27600 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _476_
timestamp 1676037725
transform 1 0 28704 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _477_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28428 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _478_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 30268 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _479_
timestamp 1676037725
transform -1 0 30360 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _480_
timestamp 1676037725
transform 1 0 27876 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _481_
timestamp 1676037725
transform 1 0 27508 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _482_
timestamp 1676037725
transform 1 0 28704 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _483_
timestamp 1676037725
transform -1 0 29900 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _484_
timestamp 1676037725
transform 1 0 29716 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _485_
timestamp 1676037725
transform 1 0 27416 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _486_
timestamp 1676037725
transform 1 0 27600 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _487_
timestamp 1676037725
transform -1 0 29256 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _488_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 29256 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _489_
timestamp 1676037725
transform -1 0 30360 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _490_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 29440 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_2  _491_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 27600 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _492_
timestamp 1676037725
transform 1 0 28704 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _493_
timestamp 1676037725
transform 1 0 14352 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _494_
timestamp 1676037725
transform -1 0 17848 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _495_
timestamp 1676037725
transform 1 0 19412 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and4_4  _496_
timestamp 1676037725
transform -1 0 14444 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _497_
timestamp 1676037725
transform -1 0 13800 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _498_
timestamp 1676037725
transform 1 0 9108 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _499_
timestamp 1676037725
transform 1 0 9752 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _500_
timestamp 1676037725
transform 1 0 7084 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _501_
timestamp 1676037725
transform -1 0 3404 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _502_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3128 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _503_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2944 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _504_
timestamp 1676037725
transform 1 0 5796 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _505_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2116 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _506_
timestamp 1676037725
transform -1 0 3496 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and4_2  _507_
timestamp 1676037725
transform -1 0 4692 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _508_
timestamp 1676037725
transform -1 0 4232 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _509_
timestamp 1676037725
transform -1 0 5244 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _510_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 5244 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _511_
timestamp 1676037725
transform -1 0 2576 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _512_
timestamp 1676037725
transform 1 0 2944 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _513_
timestamp 1676037725
transform 1 0 3956 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _514_
timestamp 1676037725
transform 1 0 5152 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _515_
timestamp 1676037725
transform 1 0 2760 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _516_
timestamp 1676037725
transform -1 0 5888 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _517_
timestamp 1676037725
transform -1 0 1932 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _518_
timestamp 1676037725
transform 1 0 2668 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _519_
timestamp 1676037725
transform -1 0 2300 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _520_
timestamp 1676037725
transform 1 0 2944 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _521_
timestamp 1676037725
transform 1 0 19044 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _522_
timestamp 1676037725
transform 1 0 19964 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _523_
timestamp 1676037725
transform 1 0 23276 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _524_
timestamp 1676037725
transform 1 0 19412 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _525_
timestamp 1676037725
transform -1 0 25024 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_4  _526_
timestamp 1676037725
transform 1 0 17848 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__nand2_2  _527_
timestamp 1676037725
transform -1 0 17204 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _528_
timestamp 1676037725
transform 1 0 16836 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _529_
timestamp 1676037725
transform 1 0 16836 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _530_
timestamp 1676037725
transform 1 0 16836 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _531_
timestamp 1676037725
transform 1 0 15548 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_2  _532_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 14904 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _533_
timestamp 1676037725
transform 1 0 11776 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _534_
timestamp 1676037725
transform 1 0 11960 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _535_
timestamp 1676037725
transform 1 0 12972 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _536_
timestamp 1676037725
transform 1 0 14260 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _537_
timestamp 1676037725
transform 1 0 16836 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _538_
timestamp 1676037725
transform 1 0 16836 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _539_
timestamp 1676037725
transform 1 0 15456 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _540_
timestamp 1676037725
transform -1 0 16376 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _541_
timestamp 1676037725
transform 1 0 9200 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _542_
timestamp 1676037725
transform 1 0 14812 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _543_
timestamp 1676037725
transform 1 0 7636 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _544_
timestamp 1676037725
transform 1 0 7544 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _545_
timestamp 1676037725
transform -1 0 15640 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _546_
timestamp 1676037725
transform 1 0 12696 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _547_
timestamp 1676037725
transform 1 0 14260 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _548_
timestamp 1676037725
transform 1 0 12604 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _549_
timestamp 1676037725
transform 1 0 14720 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _550_
timestamp 1676037725
transform 1 0 21988 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _551_
timestamp 1676037725
transform 1 0 22356 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _552_
timestamp 1676037725
transform 1 0 20608 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _553_
timestamp 1676037725
transform 1 0 19504 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _554_
timestamp 1676037725
transform 1 0 21988 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _555_
timestamp 1676037725
transform 1 0 24656 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _556_
timestamp 1676037725
transform 1 0 24748 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _557_
timestamp 1676037725
transform 1 0 24564 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _558_
timestamp 1676037725
transform -1 0 20332 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _559_
timestamp 1676037725
transform 1 0 24748 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _560_
timestamp 1676037725
transform 1 0 24840 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _561_
timestamp 1676037725
transform 1 0 21988 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _562_
timestamp 1676037725
transform 1 0 22264 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _563_
timestamp 1676037725
transform 1 0 18032 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _564_
timestamp 1676037725
transform 1 0 19412 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _565_
timestamp 1676037725
transform 1 0 17848 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _566_
timestamp 1676037725
transform 1 0 19412 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _567_
timestamp 1676037725
transform -1 0 14720 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _568_
timestamp 1676037725
transform 1 0 9476 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _569_
timestamp 1676037725
transform 1 0 9384 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _570_
timestamp 1676037725
transform 1 0 8096 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _571_
timestamp 1676037725
transform 1 0 6900 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _572_
timestamp 1676037725
transform -1 0 16652 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _573_
timestamp 1676037725
transform 1 0 9476 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _574_
timestamp 1676037725
transform 1 0 11684 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _575_
timestamp 1676037725
transform 1 0 10948 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _576_
timestamp 1676037725
transform -1 0 16376 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _577_
timestamp 1676037725
transform 1 0 17388 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _578_
timestamp 1676037725
transform 1 0 19504 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _579_
timestamp 1676037725
transform -1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _580_
timestamp 1676037725
transform 1 0 3312 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _581_
timestamp 1676037725
transform 1 0 2576 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _582_
timestamp 1676037725
transform -1 0 3496 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _583_
timestamp 1676037725
transform -1 0 4232 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _584_
timestamp 1676037725
transform 1 0 7360 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _585_
timestamp 1676037725
transform 1 0 8188 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _586_
timestamp 1676037725
transform -1 0 10304 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _587_
timestamp 1676037725
transform 1 0 6716 0 -1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _588_
timestamp 1676037725
transform 1 0 6164 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _589_
timestamp 1676037725
transform -1 0 7728 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _590_
timestamp 1676037725
transform 1 0 6164 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _591_
timestamp 1676037725
transform 1 0 11684 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _592_
timestamp 1676037725
transform 1 0 13984 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _593_
timestamp 1676037725
transform 1 0 14444 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _594_
timestamp 1676037725
transform -1 0 14260 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _595_
timestamp 1676037725
transform 1 0 27140 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _596_
timestamp 1676037725
transform 1 0 28060 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _597_
timestamp 1676037725
transform 1 0 28060 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _598_
timestamp 1676037725
transform 1 0 28060 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _599_
timestamp 1676037725
transform 1 0 27968 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _600_
timestamp 1676037725
transform -1 0 20608 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _601_
timestamp 1676037725
transform 1 0 17756 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _602_
timestamp 1676037725
transform 1 0 20332 0 -1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _603_
timestamp 1676037725
transform 1 0 22632 0 1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _604_
timestamp 1676037725
transform -1 0 12880 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _605_
timestamp 1676037725
transform 1 0 7452 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _606_
timestamp 1676037725
transform 1 0 4876 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _607_
timestamp 1676037725
transform 1 0 4876 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _608_
timestamp 1676037725
transform 1 0 8924 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _609_
timestamp 1676037725
transform 1 0 4876 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _610_
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _611_
timestamp 1676037725
transform 1 0 4692 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _612_
timestamp 1676037725
transform -1 0 5980 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _613_
timestamp 1676037725
transform 1 0 28060 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _614_
timestamp 1676037725
transform 1 0 28704 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _615_
timestamp 1676037725
transform -1 0 28336 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _616_
timestamp 1676037725
transform 1 0 16836 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _617_
timestamp 1676037725
transform 1 0 19228 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _618_
timestamp 1676037725
transform 1 0 21988 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _619_
timestamp 1676037725
transform 1 0 22816 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _620_
timestamp 1676037725
transform 1 0 25024 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _621_
timestamp 1676037725
transform 1 0 27324 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _622_
timestamp 1676037725
transform -1 0 16376 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _623_
timestamp 1676037725
transform 1 0 17480 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _624_
timestamp 1676037725
transform -1 0 19688 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _625_
timestamp 1676037725
transform 1 0 19872 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _626_
timestamp 1676037725
transform -1 0 22264 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _627_
timestamp 1676037725
transform 1 0 21252 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _628_
timestamp 1676037725
transform 1 0 21988 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _629_
timestamp 1676037725
transform -1 0 22908 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _630_
timestamp 1676037725
transform 1 0 27140 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _631_
timestamp 1676037725
transform 1 0 24104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _632_
timestamp 1676037725
transform 1 0 23368 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _633_
timestamp 1676037725
transform 1 0 20700 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _634_
timestamp 1676037725
transform 1 0 18952 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _635_
timestamp 1676037725
transform -1 0 16284 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _636_
timestamp 1676037725
transform 1 0 16836 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _637_
timestamp 1676037725
transform 1 0 26036 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _638_
timestamp 1676037725
transform 1 0 29716 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _639_
timestamp 1676037725
transform -1 0 28152 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _640_
timestamp 1676037725
transform -1 0 28796 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _641_
timestamp 1676037725
transform -1 0 6808 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _642_
timestamp 1676037725
transform -1 0 5704 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _643_
timestamp 1676037725
transform -1 0 4968 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _644_
timestamp 1676037725
transform -1 0 4692 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _645_
timestamp 1676037725
transform 1 0 11040 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _646_
timestamp 1676037725
transform -1 0 8648 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _647_
timestamp 1676037725
transform -1 0 6808 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _648_
timestamp 1676037725
transform -1 0 5888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _649_
timestamp 1676037725
transform 1 0 7636 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _650_
timestamp 1676037725
transform 1 0 10672 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _651_
timestamp 1676037725
transform -1 0 11224 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _652_
timestamp 1676037725
transform 1 0 28520 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _653_
timestamp 1676037725
transform -1 0 27692 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _654_
timestamp 1676037725
transform 1 0 26404 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _655_
timestamp 1676037725
transform -1 0 23736 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _656_
timestamp 1676037725
transform -1 0 21804 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _657_
timestamp 1676037725
transform -1 0 19688 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _658_
timestamp 1676037725
transform -1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _659_
timestamp 1676037725
transform 1 0 20332 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _660_
timestamp 1676037725
transform 1 0 26772 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _661_
timestamp 1676037725
transform -1 0 28612 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _662_
timestamp 1676037725
transform -1 0 28520 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _663_
timestamp 1676037725
transform 1 0 27876 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _664_
timestamp 1676037725
transform 1 0 26496 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _665_
timestamp 1676037725
transform 1 0 28704 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _666_
timestamp 1676037725
transform 1 0 12512 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _667_
timestamp 1676037725
transform 1 0 15272 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _668_
timestamp 1676037725
transform 1 0 13340 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _669_
timestamp 1676037725
transform -1 0 12696 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _670_
timestamp 1676037725
transform 1 0 5980 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _671_
timestamp 1676037725
transform -1 0 5612 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _672_
timestamp 1676037725
transform -1 0 5796 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _673_
timestamp 1676037725
transform -1 0 6072 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _674_
timestamp 1676037725
transform -1 0 7544 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _675_
timestamp 1676037725
transform 1 0 8188 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _676_
timestamp 1676037725
transform 1 0 10304 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _677_
timestamp 1676037725
transform 1 0 23460 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _678_
timestamp 1676037725
transform 1 0 24472 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _679_
timestamp 1676037725
transform 1 0 24564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _680_
timestamp 1676037725
transform 1 0 24656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _681_
timestamp 1676037725
transform 1 0 6532 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _682_
timestamp 1676037725
transform -1 0 11224 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _683_
timestamp 1676037725
transform 1 0 14076 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _684_
timestamp 1676037725
transform -1 0 3312 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _685_
timestamp 1676037725
transform -1 0 2576 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _686_
timestamp 1676037725
transform -1 0 2852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _687_
timestamp 1676037725
transform -1 0 3496 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _688_
timestamp 1676037725
transform -1 0 5336 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _689_
timestamp 1676037725
transform 1 0 9108 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _690_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 9752 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _691_
timestamp 1676037725
transform 1 0 9292 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _692_
timestamp 1676037725
transform -1 0 7636 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _693_
timestamp 1676037725
transform 1 0 4508 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _694_
timestamp 1676037725
transform 1 0 2668 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _695_
timestamp 1676037725
transform 1 0 3956 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _696_
timestamp 1676037725
transform 1 0 2852 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _697_
timestamp 1676037725
transform -1 0 3128 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _698_
timestamp 1676037725
transform 1 0 2576 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _699_
timestamp 1676037725
transform 1 0 2024 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _700_
timestamp 1676037725
transform 1 0 2668 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _701_
timestamp 1676037725
transform -1 0 14444 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _702_
timestamp 1676037725
transform 1 0 24564 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _703_
timestamp 1676037725
transform 1 0 24288 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _704_
timestamp 1676037725
transform 1 0 24564 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _705_
timestamp 1676037725
transform 1 0 23828 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _706_
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _707_
timestamp 1676037725
transform 1 0 15364 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _708_
timestamp 1676037725
transform 1 0 16928 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _709_
timestamp 1676037725
transform 1 0 18768 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _710_
timestamp 1676037725
transform -1 0 20884 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _711_
timestamp 1676037725
transform -1 0 15732 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_1  _712_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _713_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _714_
timestamp 1676037725
transform -1 0 18676 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _715_
timestamp 1676037725
transform 1 0 16836 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _716_
timestamp 1676037725
transform 1 0 19044 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _717_
timestamp 1676037725
transform 1 0 20516 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _718_
timestamp 1676037725
transform 1 0 20424 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _719_
timestamp 1676037725
transform 1 0 21988 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _720_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21436 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _721_
timestamp 1676037725
transform 1 0 19596 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _722_
timestamp 1676037725
transform 1 0 23184 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _723_
timestamp 1676037725
transform 1 0 18400 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _724_
timestamp 1676037725
transform 1 0 24564 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _725_
timestamp 1676037725
transform 1 0 16560 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _726_
timestamp 1676037725
transform 1 0 15824 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _727_
timestamp 1676037725
transform 1 0 16192 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _728_
timestamp 1676037725
transform 1 0 14904 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _729_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11684 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _730_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11776 0 1 17408
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _731_
timestamp 1676037725
transform 1 0 12880 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _732_
timestamp 1676037725
transform 1 0 13156 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _733_
timestamp 1676037725
transform 1 0 21988 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_2  _734_
timestamp 1676037725
transform 1 0 26956 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _735_
timestamp 1676037725
transform 1 0 24748 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _736_
timestamp 1676037725
transform 1 0 22172 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _737_
timestamp 1676037725
transform 1 0 21712 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _738_
timestamp 1676037725
transform 1 0 19412 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _739_
timestamp 1676037725
transform 1 0 16652 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _740_
timestamp 1676037725
transform 1 0 16836 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _741_
timestamp 1676037725
transform 1 0 26128 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _742_
timestamp 1676037725
transform -1 0 30084 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _743_
timestamp 1676037725
transform 1 0 27876 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _744_
timestamp 1676037725
transform 1 0 28336 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _745_
timestamp 1676037725
transform -1 0 6072 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _746_
timestamp 1676037725
transform 1 0 4140 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _747_
timestamp 1676037725
transform 1 0 4140 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _748_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5060 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _749_
timestamp 1676037725
transform -1 0 13616 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _750_
timestamp 1676037725
transform 1 0 9108 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _751_
timestamp 1676037725
transform -1 0 7268 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _752_
timestamp 1676037725
transform 1 0 5336 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _753_
timestamp 1676037725
transform 1 0 7728 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _754_
timestamp 1676037725
transform 1 0 10764 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _755_
timestamp 1676037725
transform 1 0 9752 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_2  _756_
timestamp 1676037725
transform 1 0 24564 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _757_
timestamp 1676037725
transform -1 0 29440 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _758_
timestamp 1676037725
transform 1 0 28060 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _759_
timestamp 1676037725
transform 1 0 27140 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _760_
timestamp 1676037725
transform -1 0 16376 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _761_
timestamp 1676037725
transform 1 0 14904 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _762_
timestamp 1676037725
transform -1 0 17020 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _763_
timestamp 1676037725
transform 1 0 9108 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _764_
timestamp 1676037725
transform -1 0 15916 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _765_
timestamp 1676037725
transform 1 0 6992 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _766_
timestamp 1676037725
transform 1 0 6808 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _767_
timestamp 1676037725
transform 1 0 12236 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _768_
timestamp 1676037725
transform 1 0 13156 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _769_
timestamp 1676037725
transform 1 0 12052 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _770_
timestamp 1676037725
transform 1 0 12880 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_2  _771_
timestamp 1676037725
transform 1 0 22448 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _772_
timestamp 1676037725
transform -1 0 22448 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _773_
timestamp 1676037725
transform -1 0 19964 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _774_
timestamp 1676037725
transform 1 0 18400 0 -1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _775_
timestamp 1676037725
transform 1 0 20424 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _776_
timestamp 1676037725
transform 1 0 27600 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _777_
timestamp 1676037725
transform 1 0 28336 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _778_
timestamp 1676037725
transform 1 0 28152 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _779_
timestamp 1676037725
transform 1 0 28152 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _780_
timestamp 1676037725
transform 1 0 27140 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _781_
timestamp 1676037725
transform -1 0 30268 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _782_
timestamp 1676037725
transform 1 0 27232 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _783_
timestamp 1676037725
transform 1 0 20056 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _784_
timestamp 1676037725
transform 1 0 22172 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _785_
timestamp 1676037725
transform 1 0 19688 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _786_
timestamp 1676037725
transform 1 0 21988 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _787_
timestamp 1676037725
transform 1 0 24564 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _788_
timestamp 1676037725
transform 1 0 24472 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _789_
timestamp 1676037725
transform 1 0 24564 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _790_
timestamp 1676037725
transform 1 0 24564 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _791_
timestamp 1676037725
transform 1 0 24656 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _792_
timestamp 1676037725
transform 1 0 21344 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _793_
timestamp 1676037725
transform 1 0 21804 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_2  _794_
timestamp 1676037725
transform 1 0 12052 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _795_
timestamp 1676037725
transform -1 0 16284 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _796_
timestamp 1676037725
transform 1 0 14260 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _797_
timestamp 1676037725
transform 1 0 11316 0 1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _798_
timestamp 1676037725
transform 1 0 6532 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _799_
timestamp 1676037725
transform 1 0 5980 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _800_
timestamp 1676037725
transform 1 0 5796 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _801_
timestamp 1676037725
transform 1 0 6532 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _802_
timestamp 1676037725
transform 1 0 6624 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _803_
timestamp 1676037725
transform 1 0 8280 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _804_
timestamp 1676037725
transform 1 0 10856 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _805_
timestamp 1676037725
transform 1 0 17480 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _806_
timestamp 1676037725
transform 1 0 18860 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _807_
timestamp 1676037725
transform 1 0 17296 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _808_
timestamp 1676037725
transform 1 0 18492 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _809_
timestamp 1676037725
transform 1 0 9016 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _810_
timestamp 1676037725
transform 1 0 9016 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _811_
timestamp 1676037725
transform 1 0 7360 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _812_
timestamp 1676037725
transform 1 0 6716 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _813_
timestamp 1676037725
transform 1 0 8832 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _814_
timestamp 1676037725
transform 1 0 11132 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _815_
timestamp 1676037725
transform 1 0 10580 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _816_
timestamp 1676037725
transform -1 0 16376 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _817_
timestamp 1676037725
transform 1 0 18032 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _818_
timestamp 1676037725
transform 1 0 20884 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _819_
timestamp 1676037725
transform 1 0 24104 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _820_
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _821_
timestamp 1676037725
transform 1 0 24288 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _822_
timestamp 1676037725
transform 1 0 24748 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _823_
timestamp 1676037725
transform 1 0 7176 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _824_
timestamp 1676037725
transform -1 0 8464 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _825_
timestamp 1676037725
transform 1 0 11868 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _826_
timestamp 1676037725
transform 1 0 2484 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _827_
timestamp 1676037725
transform 1 0 1840 0 -1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _828_
timestamp 1676037725
transform 1 0 2024 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _829_
timestamp 1676037725
transform 1 0 2668 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _830_
timestamp 1676037725
transform -1 0 6072 0 -1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _831_
timestamp 1676037725
transform 1 0 9108 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__183_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15088 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__203_
timestamp 1676037725
transform -1 0 12604 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__222_
timestamp 1676037725
transform 1 0 23276 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__245_
timestamp 1676037725
transform -1 0 10580 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__264_
timestamp 1676037725
transform 1 0 23368 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1676037725
transform 1 0 3496 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__183_
timestamp 1676037725
transform -1 0 14812 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__203_
timestamp 1676037725
transform -1 0 9660 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__222_
timestamp 1676037725
transform -1 0 22632 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__245_
timestamp 1676037725
transform -1 0 9660 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__264_
timestamp 1676037725
transform -1 0 22632 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1676037725
transform -1 0 4416 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__183_
timestamp 1676037725
transform 1 0 15640 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__203_
timestamp 1676037725
transform 1 0 10396 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__222_
timestamp 1676037725
transform 1 0 23368 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__245_
timestamp 1676037725
transform -1 0 7084 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__264_
timestamp 1676037725
transform 1 0 24564 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1676037725
transform -1 0 4416 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_4  fanout16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 12604 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15824 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  fanout18 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 6992 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  fanout19
timestamp 1676037725
transform 1 0 6532 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  fanout20
timestamp 1676037725
transform 1 0 6532 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_12  fanout21
timestamp 1676037725
transform 1 0 20976 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  fanout22
timestamp 1676037725
transform -1 0 18584 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  fanout23
timestamp 1676037725
transform 1 0 6164 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 5060 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  fanout25
timestamp 1676037725
transform 1 0 4508 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout26
timestamp 1676037725
transform -1 0 4508 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout27
timestamp 1676037725
transform -1 0 23828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout28
timestamp 1676037725
transform 1 0 14904 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout29
timestamp 1676037725
transform 1 0 22816 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout30 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21988 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout31
timestamp 1676037725
transform -1 0 15180 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout32
timestamp 1676037725
transform 1 0 14628 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout33
timestamp 1676037725
transform 1 0 16560 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout34
timestamp 1676037725
transform -1 0 5060 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_8  fanout35 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 17848 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout36
timestamp 1676037725
transform 1 0 25852 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout37
timestamp 1676037725
transform -1 0 17940 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout38 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18308 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold1
timestamp 1676037725
transform -1 0 4784 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold2
timestamp 1676037725
transform 1 0 5244 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold3
timestamp 1676037725
transform 1 0 10120 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold4
timestamp 1676037725
transform -1 0 13340 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold5
timestamp 1676037725
transform -1 0 5244 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10120 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  input2
timestamp 1676037725
transform 1 0 14260 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1676037725
transform 1 0 18032 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 1676037725
transform 1 0 21988 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1676037725
transform 1 0 25944 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  input6
timestamp 1676037725
transform -1 0 29256 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  input7
timestamp 1676037725
transform 1 0 6532 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output8
timestamp 1676037725
transform 1 0 29808 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output9
timestamp 1676037725
transform 1 0 29808 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output10
timestamp 1676037725
transform 1 0 29808 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output11
timestamp 1676037725
transform -1 0 30360 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output12
timestamp 1676037725
transform 1 0 29808 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output13
timestamp 1676037725
transform 1 0 29808 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output14
timestamp 1676037725
transform 1 0 29808 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output15
timestamp 1676037725
transform 1 0 29808 0 -1 29376
box -38 -48 590 592
<< labels >>
flabel metal2 s 2134 31200 2190 32000 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 10046 31200 10102 32000 0 FreeSans 224 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 14002 31200 14058 32000 0 FreeSans 224 90 0 0 io_in[1]
port 2 nsew signal input
flabel metal2 s 17958 31200 18014 32000 0 FreeSans 224 90 0 0 io_in[2]
port 3 nsew signal input
flabel metal2 s 21914 31200 21970 32000 0 FreeSans 224 90 0 0 io_in[3]
port 4 nsew signal input
flabel metal2 s 25870 31200 25926 32000 0 FreeSans 224 90 0 0 io_in[4]
port 5 nsew signal input
flabel metal2 s 29826 31200 29882 32000 0 FreeSans 224 90 0 0 io_in[5]
port 6 nsew signal input
flabel metal3 s 31200 2048 32000 2168 0 FreeSans 480 0 0 0 io_out[0]
port 7 nsew signal tristate
flabel metal3 s 31200 5992 32000 6112 0 FreeSans 480 0 0 0 io_out[1]
port 8 nsew signal tristate
flabel metal3 s 31200 9936 32000 10056 0 FreeSans 480 0 0 0 io_out[2]
port 9 nsew signal tristate
flabel metal3 s 31200 13880 32000 14000 0 FreeSans 480 0 0 0 io_out[3]
port 10 nsew signal tristate
flabel metal3 s 31200 17824 32000 17944 0 FreeSans 480 0 0 0 io_out[4]
port 11 nsew signal tristate
flabel metal3 s 31200 21768 32000 21888 0 FreeSans 480 0 0 0 io_out[5]
port 12 nsew signal tristate
flabel metal3 s 31200 25712 32000 25832 0 FreeSans 480 0 0 0 io_out[6]
port 13 nsew signal tristate
flabel metal3 s 31200 29656 32000 29776 0 FreeSans 480 0 0 0 io_out[7]
port 14 nsew signal tristate
flabel metal2 s 6090 31200 6146 32000 0 FreeSans 224 90 0 0 rst
port 15 nsew signal input
flabel metal4 s 4658 2128 4978 29424 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 12086 2128 12406 29424 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 19514 2128 19834 29424 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 26942 2128 27262 29424 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 8372 2128 8692 29424 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 15800 2128 16120 29424 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 23228 2128 23548 29424 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 30656 2128 30976 29424 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32000 32000
<< end >>
