magic
tech sky130B
magscale 1 2
timestamp 1680173957
<< nwell >>
rect 1066 32901 34906 33467
rect 1066 31813 34906 32379
rect 1066 30725 34906 31291
rect 1066 29637 34906 30203
rect 1066 28549 34906 29115
rect 1066 27461 34906 28027
rect 1066 26373 34906 26939
rect 1066 25285 34906 25851
rect 1066 24197 34906 24763
rect 1066 23109 34906 23675
rect 1066 22021 34906 22587
rect 1066 20933 34906 21499
rect 1066 19845 34906 20411
rect 1066 18757 34906 19323
rect 1066 17669 34906 18235
rect 1066 16581 34906 17147
rect 1066 15493 34906 16059
rect 1066 14405 34906 14971
rect 1066 13317 34906 13883
rect 1066 12229 34906 12795
rect 1066 11141 34906 11707
rect 1066 10053 34906 10619
rect 1066 8965 34906 9531
rect 1066 7877 34906 8443
rect 1066 6789 34906 7355
rect 1066 5701 34906 6267
rect 1066 4613 34906 5179
rect 1066 3525 34906 4091
rect 1066 2437 34906 3003
<< obsli1 >>
rect 1104 2159 34868 33745
<< obsm1 >>
rect 1104 2128 35027 33776
<< metal2 >>
rect 1766 35200 1822 36000
rect 4710 35200 4766 36000
rect 7654 35200 7710 36000
rect 10598 35200 10654 36000
rect 13542 35200 13598 36000
rect 16486 35200 16542 36000
rect 19430 35200 19486 36000
rect 22374 35200 22430 36000
rect 25318 35200 25374 36000
rect 28262 35200 28318 36000
rect 31206 35200 31262 36000
rect 34150 35200 34206 36000
rect 1214 0 1270 800
rect 2502 0 2558 800
rect 3790 0 3846 800
rect 5078 0 5134 800
rect 6366 0 6422 800
rect 7654 0 7710 800
rect 8942 0 8998 800
rect 10230 0 10286 800
rect 11518 0 11574 800
rect 12806 0 12862 800
rect 14094 0 14150 800
rect 15382 0 15438 800
rect 16670 0 16726 800
rect 17958 0 18014 800
rect 19246 0 19302 800
rect 20534 0 20590 800
rect 21822 0 21878 800
rect 23110 0 23166 800
rect 24398 0 24454 800
rect 25686 0 25742 800
rect 26974 0 27030 800
rect 28262 0 28318 800
rect 29550 0 29606 800
rect 30838 0 30894 800
rect 32126 0 32182 800
rect 33414 0 33470 800
rect 34702 0 34758 800
<< obsm2 >>
rect 1216 35144 1710 35306
rect 1878 35144 4654 35306
rect 4822 35144 7598 35306
rect 7766 35144 10542 35306
rect 10710 35144 13486 35306
rect 13654 35144 16430 35306
rect 16598 35144 19374 35306
rect 19542 35144 22318 35306
rect 22486 35144 25262 35306
rect 25430 35144 28206 35306
rect 28374 35144 31150 35306
rect 31318 35144 34094 35306
rect 34262 35144 35021 35306
rect 1216 856 35021 35144
rect 1326 734 2446 856
rect 2614 734 3734 856
rect 3902 734 5022 856
rect 5190 734 6310 856
rect 6478 734 7598 856
rect 7766 734 8886 856
rect 9054 734 10174 856
rect 10342 734 11462 856
rect 11630 734 12750 856
rect 12918 734 14038 856
rect 14206 734 15326 856
rect 15494 734 16614 856
rect 16782 734 17902 856
rect 18070 734 19190 856
rect 19358 734 20478 856
rect 20646 734 21766 856
rect 21934 734 23054 856
rect 23222 734 24342 856
rect 24510 734 25630 856
rect 25798 734 26918 856
rect 27086 734 28206 856
rect 28374 734 29494 856
rect 29662 734 30782 856
rect 30950 734 32070 856
rect 32238 734 33358 856
rect 33526 734 34646 856
rect 34814 734 35021 856
<< metal3 >>
rect 35200 17824 36000 17944
<< obsm3 >>
rect 5166 18024 35200 33761
rect 5166 17744 35120 18024
rect 5166 2143 35200 17744
<< metal4 >>
rect 5164 2128 5484 33776
rect 9384 2128 9704 33776
rect 13605 2128 13925 33776
rect 17825 2128 18145 33776
rect 22046 2128 22366 33776
rect 26266 2128 26586 33776
rect 30487 2128 30807 33776
rect 34707 2128 35027 33776
<< obsm4 >>
rect 24899 23155 24965 30837
<< labels >>
rlabel metal2 s 1766 35200 1822 36000 6 clk
port 1 nsew signal input
rlabel metal2 s 7654 35200 7710 36000 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 10598 35200 10654 36000 6 io_in[1]
port 3 nsew signal input
rlabel metal2 s 13542 35200 13598 36000 6 io_in[2]
port 4 nsew signal input
rlabel metal2 s 16486 35200 16542 36000 6 io_in[3]
port 5 nsew signal input
rlabel metal2 s 19430 35200 19486 36000 6 io_in[4]
port 6 nsew signal input
rlabel metal2 s 22374 35200 22430 36000 6 io_in[5]
port 7 nsew signal input
rlabel metal2 s 25318 35200 25374 36000 6 io_in[6]
port 8 nsew signal input
rlabel metal2 s 28262 35200 28318 36000 6 io_in[7]
port 9 nsew signal input
rlabel metal2 s 31206 35200 31262 36000 6 io_in[8]
port 10 nsew signal input
rlabel metal2 s 34150 35200 34206 36000 6 io_in[9]
port 11 nsew signal input
rlabel metal3 s 35200 17824 36000 17944 6 io_oeb
port 12 nsew signal output
rlabel metal2 s 1214 0 1270 800 6 io_out[0]
port 13 nsew signal output
rlabel metal2 s 14094 0 14150 800 6 io_out[10]
port 14 nsew signal output
rlabel metal2 s 15382 0 15438 800 6 io_out[11]
port 15 nsew signal output
rlabel metal2 s 16670 0 16726 800 6 io_out[12]
port 16 nsew signal output
rlabel metal2 s 17958 0 18014 800 6 io_out[13]
port 17 nsew signal output
rlabel metal2 s 19246 0 19302 800 6 io_out[14]
port 18 nsew signal output
rlabel metal2 s 20534 0 20590 800 6 io_out[15]
port 19 nsew signal output
rlabel metal2 s 21822 0 21878 800 6 io_out[16]
port 20 nsew signal output
rlabel metal2 s 23110 0 23166 800 6 io_out[17]
port 21 nsew signal output
rlabel metal2 s 24398 0 24454 800 6 io_out[18]
port 22 nsew signal output
rlabel metal2 s 25686 0 25742 800 6 io_out[19]
port 23 nsew signal output
rlabel metal2 s 2502 0 2558 800 6 io_out[1]
port 24 nsew signal output
rlabel metal2 s 26974 0 27030 800 6 io_out[20]
port 25 nsew signal output
rlabel metal2 s 28262 0 28318 800 6 io_out[21]
port 26 nsew signal output
rlabel metal2 s 29550 0 29606 800 6 io_out[22]
port 27 nsew signal output
rlabel metal2 s 30838 0 30894 800 6 io_out[23]
port 28 nsew signal output
rlabel metal2 s 32126 0 32182 800 6 io_out[24]
port 29 nsew signal output
rlabel metal2 s 33414 0 33470 800 6 io_out[25]
port 30 nsew signal output
rlabel metal2 s 34702 0 34758 800 6 io_out[26]
port 31 nsew signal output
rlabel metal2 s 3790 0 3846 800 6 io_out[2]
port 32 nsew signal output
rlabel metal2 s 5078 0 5134 800 6 io_out[3]
port 33 nsew signal output
rlabel metal2 s 6366 0 6422 800 6 io_out[4]
port 34 nsew signal output
rlabel metal2 s 7654 0 7710 800 6 io_out[5]
port 35 nsew signal output
rlabel metal2 s 8942 0 8998 800 6 io_out[6]
port 36 nsew signal output
rlabel metal2 s 10230 0 10286 800 6 io_out[7]
port 37 nsew signal output
rlabel metal2 s 11518 0 11574 800 6 io_out[8]
port 38 nsew signal output
rlabel metal2 s 12806 0 12862 800 6 io_out[9]
port 39 nsew signal output
rlabel metal2 s 4710 35200 4766 36000 6 rst
port 40 nsew signal input
rlabel metal4 s 5164 2128 5484 33776 6 vccd1
port 41 nsew power bidirectional
rlabel metal4 s 13605 2128 13925 33776 6 vccd1
port 41 nsew power bidirectional
rlabel metal4 s 22046 2128 22366 33776 6 vccd1
port 41 nsew power bidirectional
rlabel metal4 s 30487 2128 30807 33776 6 vccd1
port 41 nsew power bidirectional
rlabel metal4 s 9384 2128 9704 33776 6 vssd1
port 42 nsew ground bidirectional
rlabel metal4 s 17825 2128 18145 33776 6 vssd1
port 42 nsew ground bidirectional
rlabel metal4 s 26266 2128 26586 33776 6 vssd1
port 42 nsew ground bidirectional
rlabel metal4 s 34707 2128 35027 33776 6 vssd1
port 42 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 36000 36000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2913376
string GDS_FILE /run/media/tholin/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/AS5401/runs/23_03_30_12_55/results/signoff/tholin_avalonsemi_5401.magic.gds
string GDS_START 884056
<< end >>

